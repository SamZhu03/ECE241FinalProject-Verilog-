module rom_w0(
input  clk,
input [16:0] addr,
output signed [15:0] dout);
(*rom_style = "block" *) reg signed [15:0] data;
always @(posedge clk) 
begin
    case(addr)
      0:data<=16'd80;
      1:data<=-16'd209;
      2:data<=-16'd1392;
      3:data<=-16'd2403;
      4:data<=-16'd2322;
      5:data<=-16'd3031;
      6:data<=-16'd5844;
      7:data<=-16'd9119;
      8:data<=-16'd9652;
      9:data<=-16'd8859;
      10:data<=-16'd10134;
      11:data<=-16'd11201;
      12:data<=-16'd10712;
      13:data<=-16'd10487;
      14:data<=-16'd10049;
      15:data<=-16'd10921;
      16:data<=-16'd13678;
      17:data<=-16'd14257;
      18:data<=-16'd13673;
      19:data<=-16'd14827;
      20:data<=-16'd15418;
      21:data<=-16'd15121;
      22:data<=-16'd14775;
      23:data<=-16'd13794;
      24:data<=-16'd13794;
      25:data<=-16'd13873;
      26:data<=-16'd12474;
      27:data<=-16'd12681;
      28:data<=-16'd14020;
      29:data<=-16'd13700;
      30:data<=-16'd13412;
      31:data<=-16'd13292;
      32:data<=-16'd12605;
      33:data<=-16'd12618;
      34:data<=-16'd12245;
      35:data<=-16'd11732;
      36:data<=-16'd12451;
      37:data<=-16'd12267;
      38:data<=-16'd11674;
      39:data<=-16'd12283;
      40:data<=-16'd11747;
      41:data<=-16'd10646;
      42:data<=-16'd10607;
      43:data<=-16'd8915;
      44:data<=-16'd5727;
      45:data<=-16'd4573;
      46:data<=-16'd5018;
      47:data<=-16'd4595;
      48:data<=-16'd4041;
      49:data<=-16'd4707;
      50:data<=-16'd4758;
      51:data<=-16'd3792;
      52:data<=-16'd4071;
      53:data<=-16'd3988;
      54:data<=-16'd1986;
      55:data<=-16'd1269;
      56:data<=-16'd1944;
      57:data<=-16'd1572;
      58:data<=-16'd1283;
      59:data<=-16'd1679;
      60:data<=-16'd2079;
      61:data<=-16'd3040;
      62:data<=-16'd3694;
      63:data<=-16'd3397;
      64:data<=-16'd3310;
      65:data<=-16'd3139;
      66:data<=-16'd2699;
      67:data<=-16'd2883;
      68:data<=-16'd3204;
      69:data<=-16'd3673;
      70:data<=-16'd4308;
      71:data<=-16'd3826;
      72:data<=-16'd3466;
      73:data<=-16'd4262;
      74:data<=-16'd4138;
      75:data<=-16'd3479;
      76:data<=-16'd3556;
      77:data<=-16'd3739;
      78:data<=-16'd4701;
      79:data<=-16'd5203;
      80:data<=-16'd4399;
      81:data<=-16'd6604;
      82:data<=-16'd10604;
      83:data<=-16'd10558;
      84:data<=-16'd9154;
      85:data<=-16'd9940;
      86:data<=-16'd10349;
      87:data<=-16'd10108;
      88:data<=-16'd9884;
      89:data<=-16'd8766;
      90:data<=-16'd9172;
      91:data<=-16'd11897;
      92:data<=-16'd12754;
      93:data<=-16'd11414;
      94:data<=-16'd11301;
      95:data<=-16'd11997;
      96:data<=-16'd11847;
      97:data<=-16'd11209;
      98:data<=-16'd10322;
      99:data<=-16'd9682;
      100:data<=-16'd9271;
      101:data<=-16'd8508;
      102:data<=-16'd8543;
      103:data<=-16'd9207;
      104:data<=-16'd9075;
      105:data<=-16'd8871;
      106:data<=-16'd8454;
      107:data<=-16'd7545;
      108:data<=-16'd7241;
      109:data<=-16'd6587;
      110:data<=-16'd6214;
      111:data<=-16'd7715;
      112:data<=-16'd8031;
      113:data<=-16'd6874;
      114:data<=-16'd7131;
      115:data<=-16'd6583;
      116:data<=-16'd5218;
      117:data<=-16'd5835;
      118:data<=-16'd4208;
      119:data<=16'd732;
      120:data<=16'd2182;
      121:data<=16'd1221;
      122:data<=16'd2660;
      123:data<=16'd3190;
      124:data<=16'd1868;
      125:data<=16'd1865;
      126:data<=16'd2074;
      127:data<=16'd3485;
      128:data<=16'd7391;
      129:data<=16'd9139;
      130:data<=16'd8346;
      131:data<=16'd8445;
      132:data<=16'd8484;
      133:data<=16'd8184;
      134:data<=16'd8059;
      135:data<=16'd7758;
      136:data<=16'd8715;
      137:data<=16'd9826;
      138:data<=16'd9401;
      139:data<=16'd8997;
      140:data<=16'd8622;
      141:data<=16'd8331;
      142:data<=16'd8593;
      143:data<=16'd8058;
      144:data<=16'd8310;
      145:data<=16'd10008;
      146:data<=16'd10202;
      147:data<=16'd9582;
      148:data<=16'd9374;
      149:data<=16'd8727;
      150:data<=16'd8422;
      151:data<=16'd8382;
      152:data<=16'd8633;
      153:data<=16'd9632;
      154:data<=16'd10032;
      155:data<=16'd9752;
      156:data<=16'd7503;
      157:data<=16'd3183;
      158:data<=16'd2138;
      159:data<=16'd3087;
      160:data<=16'd1968;
      161:data<=16'd3042;
      162:data<=16'd5398;
      163:data<=16'd5095;
      164:data<=16'd5068;
      165:data<=16'd3768;
      166:data<=16'd441;
      167:data<=16'd65;
      168:data<=16'd566;
      169:data<=16'd532;
      170:data<=16'd2446;
      171:data<=16'd3116;
      172:data<=16'd2350;
      173:data<=16'd2617;
      174:data<=16'd2472;
      175:data<=16'd2692;
      176:data<=16'd2980;
      177:data<=16'd2499;
      178:data<=16'd3812;
      179:data<=16'd4836;
      180:data<=16'd4284;
      181:data<=16'd5053;
      182:data<=16'd4784;
      183:data<=16'd3163;
      184:data<=16'd3412;
      185:data<=16'd3626;
      186:data<=16'd3897;
      187:data<=16'd5739;
      188:data<=16'd6055;
      189:data<=16'd4787;
      190:data<=16'd4748;
      191:data<=16'd4980;
      192:data<=16'd4167;
      193:data<=16'd5030;
      194:data<=16'd9277;
      195:data<=16'd12292;
      196:data<=16'd11822;
      197:data<=16'd11521;
      198:data<=16'd11306;
      199:data<=16'd10524;
      200:data<=16'd10463;
      201:data<=16'd9433;
      202:data<=16'd9814;
      203:data<=16'd13676;
      204:data<=16'd15211;
      205:data<=16'd14113;
      206:data<=16'd13900;
      207:data<=16'd12913;
      208:data<=16'd12310;
      209:data<=16'd12584;
      210:data<=16'd11242;
      211:data<=16'd10904;
      212:data<=16'd12005;
      213:data<=16'd11394;
      214:data<=16'd10457;
      215:data<=16'd10226;
      216:data<=16'd9868;
      217:data<=16'd9421;
      218:data<=16'd8699;
      219:data<=16'd8930;
      220:data<=16'd9871;
      221:data<=16'd9805;
      222:data<=16'd9849;
      223:data<=16'd9802;
      224:data<=16'd8877;
      225:data<=16'd8370;
      226:data<=16'd7726;
      227:data<=16'd7250;
      228:data<=16'd7970;
      229:data<=16'd8681;
      230:data<=16'd9047;
      231:data<=16'd6872;
      232:data<=16'd1924;
      233:data<=16'd291;
      234:data<=16'd1322;
      235:data<=16'd561;
      236:data<=16'd898;
      237:data<=16'd2507;
      238:data<=16'd2566;
      239:data<=16'd1777;
      240:data<=-16'd397;
      241:data<=-16'd2745;
      242:data<=-16'd2852;
      243:data<=-16'd2587;
      244:data<=-16'd2305;
      245:data<=-16'd1225;
      246:data<=-16'd699;
      247:data<=-16'd702;
      248:data<=-16'd1195;
      249:data<=-16'd1905;
      250:data<=-16'd1789;
      251:data<=-16'd1764;
      252:data<=-16'd1744;
      253:data<=-16'd1048;
      254:data<=-16'd870;
      255:data<=-16'd1242;
      256:data<=-16'd1635;
      257:data<=-16'd1935;
      258:data<=-16'd1909;
      259:data<=-16'd1977;
      260:data<=-16'd1974;
      261:data<=-16'd2388;
      262:data<=-16'd3469;
      263:data<=-16'd3732;
      264:data<=-16'd4029;
      265:data<=-16'd4287;
      266:data<=-16'd3519;
      267:data<=-16'd4182;
      268:data<=-16'd3533;
      269:data<=16'd466;
      270:data<=16'd1137;
      271:data<=-16'd187;
      272:data<=16'd722;
      273:data<=-16'd259;
      274:data<=-16'd1263;
      275:data<=-16'd499;
      276:data<=-16'd1283;
      277:data<=16'd287;
      278:data<=16'd2987;
      279:data<=16'd1359;
      280:data<=16'd522;
      281:data<=16'd1510;
      282:data<=16'd902;
      283:data<=16'd1154;
      284:data<=16'd1313;
      285:data<=16'd638;
      286:data<=16'd607;
      287:data<=-16'd1049;
      288:data<=-16'd2361;
      289:data<=-16'd1597;
      290:data<=-16'd1850;
      291:data<=-16'd1941;
      292:data<=-16'd1568;
      293:data<=-16'd2159;
      294:data<=-16'd2150;
      295:data<=-16'd2787;
      296:data<=-16'd4056;
      297:data<=-16'd4026;
      298:data<=-16'd4340;
      299:data<=-16'd4434;
      300:data<=-16'd3882;
      301:data<=-16'd3973;
      302:data<=-16'd3500;
      303:data<=-16'd4222;
      304:data<=-16'd5894;
      305:data<=-16'd5292;
      306:data<=-16'd6422;
      307:data<=-16'd9682;
      308:data<=-16'd10038;
      309:data<=-16'd9465;
      310:data<=-16'd9241;
      311:data<=-16'd8884;
      312:data<=-16'd9956;
      313:data<=-16'd10248;
      314:data<=-16'd10572;
      315:data<=-16'd13065;
      316:data<=-16'd13708;
      317:data<=-16'd12775;
      318:data<=-16'd12411;
      319:data<=-16'd11235;
      320:data<=-16'd11756;
      321:data<=-16'd13661;
      322:data<=-16'd13341;
      323:data<=-16'd12713;
      324:data<=-16'd12219;
      325:data<=-16'd11054;
      326:data<=-16'd10825;
      327:data<=-16'd10383;
      328:data<=-16'd10343;
      329:data<=-16'd11753;
      330:data<=-16'd11480;
      331:data<=-16'd10405;
      332:data<=-16'd10439;
      333:data<=-16'd10040;
      334:data<=-16'd9868;
      335:data<=-16'd9429;
      336:data<=-16'd8479;
      337:data<=-16'd9397;
      338:data<=-16'd10128;
      339:data<=-16'd9668;
      340:data<=-16'd9823;
      341:data<=-16'd9191;
      342:data<=-16'd8755;
      343:data<=-16'd7829;
      344:data<=-16'd3865;
      345:data<=-16'd2729;
      346:data<=-16'd5175;
      347:data<=-16'd4758;
      348:data<=-16'd3662;
      349:data<=-16'd3632;
      350:data<=-16'd3219;
      351:data<=-16'd3066;
      352:data<=-16'd378;
      353:data<=16'd1912;
      354:data<=-16'd520;
      355:data<=-16'd1339;
      356:data<=-16'd359;
      357:data<=-16'd1221;
      358:data<=-16'd381;
      359:data<=16'd285;
      360:data<=-16'd412;
      361:data<=16'd400;
      362:data<=-16'd511;
      363:data<=-16'd2224;
      364:data<=-16'd1780;
      365:data<=-16'd1818;
      366:data<=-16'd1360;
      367:data<=-16'd479;
      368:data<=-16'd999;
      369:data<=-16'd923;
      370:data<=-16'd1685;
      371:data<=-16'd3037;
      372:data<=-16'd2297;
      373:data<=-16'd2197;
      374:data<=-16'd2569;
      375:data<=-16'd1953;
      376:data<=-16'd1876;
      377:data<=-16'd1142;
      378:data<=-16'd1351;
      379:data<=-16'd3281;
      380:data<=-16'd3078;
      381:data<=-16'd3553;
      382:data<=-16'd6602;
      383:data<=-16'd7370;
      384:data<=-16'd6172;
      385:data<=-16'd6029;
      386:data<=-16'd6566;
      387:data<=-16'd5974;
      388:data<=-16'd4431;
      389:data<=-16'd5529;
      390:data<=-16'd8244;
      391:data<=-16'd8335;
      392:data<=-16'd7241;
      393:data<=-16'd6854;
      394:data<=-16'd6943;
      395:data<=-16'd6514;
      396:data<=-16'd4358;
      397:data<=-16'd3206;
      398:data<=-16'd3363;
      399:data<=-16'd2334;
      400:data<=-16'd2270;
      401:data<=-16'd2453;
      402:data<=-16'd1242;
      403:data<=-16'd1131;
      404:data<=-16'd320;
      405:data<=16'd1401;
      406:data<=16'd1055;
      407:data<=16'd857;
      408:data<=16'd940;
      409:data<=16'd547;
      410:data<=16'd1469;
      411:data<=16'd1648;
      412:data<=16'd1691;
      413:data<=16'd3262;
      414:data<=16'd3503;
      415:data<=16'd3850;
      416:data<=16'd4681;
      417:data<=16'd3239;
      418:data<=16'd3048;
      419:data<=16'd5419;
      420:data<=16'd7926;
      421:data<=16'd10287;
      422:data<=16'd10299;
      423:data<=16'd9025;
      424:data<=16'd9144;
      425:data<=16'd8812;
      426:data<=16'd9787;
      427:data<=16'd12322;
      428:data<=16'd12240;
      429:data<=16'd12141;
      430:data<=16'd13641;
      431:data<=16'd13429;
      432:data<=16'd12484;
      433:data<=16'd11946;
      434:data<=16'd11568;
      435:data<=16'd11549;
      436:data<=16'd10642;
      437:data<=16'd10316;
      438:data<=16'd11617;
      439:data<=16'd12231;
      440:data<=16'd12337;
      441:data<=16'd12029;
      442:data<=16'd10810;
      443:data<=16'd10214;
      444:data<=16'd9885;
      445:data<=16'd10009;
      446:data<=16'd11191;
      447:data<=16'd11003;
      448:data<=16'd9840;
      449:data<=16'd9559;
      450:data<=16'd9333;
      451:data<=16'd9424;
      452:data<=16'd9188;
      453:data<=16'd7949;
      454:data<=16'd8640;
      455:data<=16'd10411;
      456:data<=16'd8757;
      457:data<=16'd4993;
      458:data<=16'd3290;
      459:data<=16'd3541;
      460:data<=16'd3635;
      461:data<=16'd3469;
      462:data<=16'd3956;
      463:data<=16'd4229;
      464:data<=16'd2814;
      465:data<=16'd934;
      466:data<=16'd305;
      467:data<=16'd140;
      468:data<=16'd50;
      469:data<=16'd117;
      470:data<=-16'd76;
      471:data<=16'd826;
      472:data<=16'd2102;
      473:data<=16'd1577;
      474:data<=16'd1265;
      475:data<=16'd1562;
      476:data<=16'd1218;
      477:data<=16'd1618;
      478:data<=16'd1509;
      479:data<=16'd1048;
      480:data<=16'd2275;
      481:data<=16'd2594;
      482:data<=16'd2419;
      483:data<=16'd2886;
      484:data<=16'd1768;
      485:data<=16'd1293;
      486:data<=16'd1351;
      487:data<=16'd731;
      488:data<=16'd2528;
      489:data<=16'd3486;
      490:data<=16'd2491;
      491:data<=16'd2863;
      492:data<=16'd1677;
      493:data<=16'd1900;
      494:data<=16'd5682;
      495:data<=16'd6310;
      496:data<=16'd6128;
      497:data<=16'd7448;
      498:data<=16'd6946;
      499:data<=16'd6661;
      500:data<=16'd6065;
      501:data<=16'd6382;
      502:data<=16'd9238;
      503:data<=16'd8822;
      504:data<=16'd8235;
      505:data<=16'd10238;
      506:data<=16'd9118;
      507:data<=16'd8745;
      508:data<=16'd9796;
      509:data<=16'd7896;
      510:data<=16'd7238;
      511:data<=16'd6949;
      512:data<=16'd5959;
      513:data<=16'd7439;
      514:data<=16'd7497;
      515:data<=16'd6332;
      516:data<=16'd6300;
      517:data<=16'd5321;
      518:data<=16'd5612;
      519:data<=16'd6009;
      520:data<=16'd4341;
      521:data<=16'd3711;
      522:data<=16'd2939;
      523:data<=16'd2428;
      524:data<=16'd3439;
      525:data<=16'd2655;
      526:data<=16'd2359;
      527:data<=16'd3280;
      528:data<=16'd1413;
      529:data<=-16'd379;
      530:data<=-16'd176;
      531:data<=-16'd1409;
      532:data<=-16'd4455;
      533:data<=-16'd6194;
      534:data<=-16'd5651;
      535:data<=-16'd5794;
      536:data<=-16'd5659;
      537:data<=-16'd4205;
      538:data<=-16'd7051;
      539:data<=-16'd11900;
      540:data<=-16'd12263;
      541:data<=-16'd11395;
      542:data<=-16'd11250;
      543:data<=-16'd10705;
      544:data<=-16'd10662;
      545:data<=-16'd10348;
      546:data<=-16'd10857;
      547:data<=-16'd12243;
      548:data<=-16'd11994;
      549:data<=-16'd11411;
      550:data<=-16'd11130;
      551:data<=-16'd10868;
      552:data<=-16'd11048;
      553:data<=-16'd10028;
      554:data<=-16'd9774;
      555:data<=-16'd11768;
      556:data<=-16'd12249;
      557:data<=-16'd11676;
      558:data<=-16'd11784;
      559:data<=-16'd11057;
      560:data<=-16'd10014;
      561:data<=-16'd9266;
      562:data<=-16'd9291;
      563:data<=-16'd10674;
      564:data<=-16'd11177;
      565:data<=-16'd10534;
      566:data<=-16'd10525;
      567:data<=-16'd10513;
      568:data<=-16'd9791;
      569:data<=-16'd7574;
      570:data<=-16'd4532;
      571:data<=-16'd4866;
      572:data<=-16'd7527;
      573:data<=-16'd7186;
      574:data<=-16'd6179;
      575:data<=-16'd6940;
      576:data<=-16'd4921;
      577:data<=-16'd1459;
      578:data<=-16'd1371;
      579:data<=-16'd2499;
      580:data<=-16'd3644;
      581:data<=-16'd5160;
      582:data<=-16'd4896;
      583:data<=-16'd4176;
      584:data<=-16'd4032;
      585:data<=-16'd3418;
      586:data<=-16'd4018;
      587:data<=-16'd4746;
      588:data<=-16'd4003;
      589:data<=-16'd4278;
      590:data<=-16'd5174;
      591:data<=-16'd5272;
      592:data<=-16'd5404;
      593:data<=-16'd5133;
      594:data<=-16'd4525;
      595:data<=-16'd4290;
      596:data<=-16'd4869;
      597:data<=-16'd6282;
      598:data<=-16'd6557;
      599:data<=-16'd6003;
      600:data<=-16'd6341;
      601:data<=-16'd5803;
      602:data<=-16'd4520;
      603:data<=-16'd4690;
      604:data<=-16'd5190;
      605:data<=-16'd5359;
      606:data<=-16'd6933;
      607:data<=-16'd9371;
      608:data<=-16'd9735;
      609:data<=-16'd8637;
      610:data<=-16'd9028;
      611:data<=-16'd8473;
      612:data<=-16'd5733;
      613:data<=-16'd6858;
      614:data<=-16'd11740;
      615:data<=-16'd13297;
      616:data<=-16'd11828;
      617:data<=-16'd11496;
      618:data<=-16'd11741;
      619:data<=-16'd11354;
      620:data<=-16'd10871;
      621:data<=-16'd10414;
      622:data<=-16'd10140;
      623:data<=-16'd10279;
      624:data<=-16'd10299;
      625:data<=-16'd9867;
      626:data<=-16'd9125;
      627:data<=-16'd8193;
      628:data<=-16'd7650;
      629:data<=-16'd7803;
      630:data<=-16'd8109;
      631:data<=-16'd8252;
      632:data<=-16'd8084;
      633:data<=-16'd7400;
      634:data<=-16'd6590;
      635:data<=-16'd6399;
      636:data<=-16'd6269;
      637:data<=-16'd5169;
      638:data<=-16'd4990;
      639:data<=-16'd6610;
      640:data<=-16'd6628;
      641:data<=-16'd5520;
      642:data<=-16'd6263;
      643:data<=-16'd5580;
      644:data<=-16'd1697;
      645:data<=16'd644;
      646:data<=-16'd226;
      647:data<=-16'd1524;
      648:data<=-16'd1999;
      649:data<=-16'd1820;
      650:data<=-16'd112;
      651:data<=16'd2905;
      652:data<=16'd4285;
      653:data<=16'd3739;
      654:data<=16'd4034;
      655:data<=16'd4598;
      656:data<=16'd4356;
      657:data<=16'd4696;
      658:data<=16'd4821;
      659:data<=16'd4067;
      660:data<=16'd4326;
      661:data<=16'd4805;
      662:data<=16'd4269;
      663:data<=16'd4575;
      664:data<=16'd5513;
      665:data<=16'd6290;
      666:data<=16'd7686;
      667:data<=16'd7333;
      668:data<=16'd5738;
      669:data<=16'd6796;
      670:data<=16'd7514;
      671:data<=16'd6783;
      672:data<=16'd8251;
      673:data<=16'd9367;
      674:data<=16'd9348;
      675:data<=16'd9629;
      676:data<=16'd8034;
      677:data<=16'd7630;
      678:data<=16'd8887;
      679:data<=16'd8152;
      680:data<=16'd9172;
      681:data<=16'd9671;
      682:data<=16'd5667;
      683:data<=16'd4614;
      684:data<=16'd6038;
      685:data<=16'd5002;
      686:data<=16'd5121;
      687:data<=16'd5435;
      688:data<=16'd4449;
      689:data<=16'd4551;
      690:data<=16'd4106;
      691:data<=16'd3518;
      692:data<=16'd3776;
      693:data<=16'd3421;
      694:data<=16'd3407;
      695:data<=16'd3418;
      696:data<=16'd3958;
      697:data<=16'd6149;
      698:data<=16'd6684;
      699:data<=16'd5962;
      700:data<=16'd6205;
      701:data<=16'd5655;
      702:data<=16'd5400;
      703:data<=16'd5741;
      704:data<=16'd4716;
      705:data<=16'd5127;
      706:data<=16'd7450;
      707:data<=16'd7524;
      708:data<=16'd6213;
      709:data<=16'd6575;
      710:data<=16'd6816;
      711:data<=16'd5800;
      712:data<=16'd6266;
      713:data<=16'd7746;
      714:data<=16'd7787;
      715:data<=16'd7561;
      716:data<=16'd7401;
      717:data<=16'd6875;
      718:data<=16'd7997;
      719:data<=16'd10076;
      720:data<=16'd10332;
      721:data<=16'd10026;
      722:data<=16'd11590;
      723:data<=16'd12725;
      724:data<=16'd11461;
      725:data<=16'd11978;
      726:data<=16'd14850;
      727:data<=16'd15044;
      728:data<=16'd13532;
      729:data<=16'd12986;
      730:data<=16'd12792;
      731:data<=16'd13717;
      732:data<=16'd14607;
      733:data<=16'd14038;
      734:data<=16'd13282;
      735:data<=16'd12158;
      736:data<=16'd11335;
      737:data<=16'd11232;
      738:data<=16'd10780;
      739:data<=16'd11300;
      740:data<=16'd12058;
      741:data<=16'd11147;
      742:data<=16'd9915;
      743:data<=16'd9224;
      744:data<=16'd9142;
      745:data<=16'd8740;
      746:data<=16'd8015;
      747:data<=16'd9169;
      748:data<=16'd10056;
      749:data<=16'd9215;
      750:data<=16'd8857;
      751:data<=16'd8313;
      752:data<=16'd8213;
      753:data<=16'd7964;
      754:data<=16'd6097;
      755:data<=16'd6854;
      756:data<=16'd7468;
      757:data<=16'd3909;
      758:data<=16'd2682;
      759:data<=16'd3290;
      760:data<=16'd2541;
      761:data<=16'd3151;
      762:data<=16'd1723;
      763:data<=-16'd1259;
      764:data<=-16'd810;
      765:data<=-16'd224;
      766:data<=-16'd684;
      767:data<=-16'd825;
      768:data<=-16'd1466;
      769:data<=-16'd1055;
      770:data<=-16'd858;
      771:data<=-16'd1662;
      772:data<=-16'd1172;
      773:data<=-16'd904;
      774:data<=-16'd831;
      775:data<=-16'd277;
      776:data<=-16'd949;
      777:data<=-16'd899;
      778:data<=-16'd258;
      779:data<=-16'd948;
      780:data<=-16'd318;
      781:data<=16'd1057;
      782:data<=16'd719;
      783:data<=16'd305;
      784:data<=16'd12;
      785:data<=-16'd414;
      786:data<=16'd473;
      787:data<=16'd773;
      788:data<=-16'd1024;
      789:data<=-16'd1171;
      790:data<=16'd196;
      791:data<=-16'd2179;
      792:data<=-16'd5662;
      793:data<=-16'd5233;
      794:data<=-16'd4337;
      795:data<=-16'd4910;
      796:data<=-16'd4972;
      797:data<=-16'd5251;
      798:data<=-16'd6438;
      799:data<=-16'd7671;
      800:data<=-16'd6246;
      801:data<=-16'd3233;
      802:data<=-16'd3707;
      803:data<=-16'd2049;
      804:data<=16'd4981;
      805:data<=16'd6111;
      806:data<=16'd2510;
      807:data<=16'd2972;
      808:data<=16'd3015;
      809:data<=16'd1745;
      810:data<=16'd2094;
      811:data<=16'd1791;
      812:data<=16'd2206;
      813:data<=16'd2331;
      814:data<=16'd1642;
      815:data<=16'd4408;
      816:data<=16'd4598;
      817:data<=-16'd99;
      818:data<=-16'd378;
      819:data<=16'd1249;
      820:data<=16'd412;
      821:data<=16'd681;
      822:data<=-16'd188;
      823:data<=-16'd1360;
      824:data<=-16'd508;
      825:data<=-16'd1706;
      826:data<=-16'd2399;
      827:data<=-16'd1744;
      828:data<=-16'd2526;
      829:data<=-16'd628;
      830:data<=-16'd2826;
      831:data<=-16'd13776;
      832:data<=-16'd18372;
      833:data<=-16'd15899;
      834:data<=-16'd15705;
      835:data<=-16'd14173;
      836:data<=-16'd12809;
      837:data<=-16'd12695;
      838:data<=-16'd10618;
      839:data<=-16'd11230;
      840:data<=-16'd11917;
      841:data<=-16'd10466;
      842:data<=-16'd11402;
      843:data<=-16'd9655;
      844:data<=-16'd8305;
      845:data<=-16'd11118;
      846:data<=-16'd8718;
      847:data<=-16'd11047;
      848:data<=-16'd23643;
      849:data<=-16'd27155;
      850:data<=-16'd24809;
      851:data<=-16'd26554;
      852:data<=-16'd24178;
      853:data<=-16'd23003;
      854:data<=-16'd27671;
      855:data<=-16'd28650;
      856:data<=-16'd26852;
      857:data<=-16'd26090;
      858:data<=-16'd25023;
      859:data<=-16'd24069;
      860:data<=-16'd22530;
      861:data<=-16'd20883;
      862:data<=-16'd19946;
      863:data<=-16'd19162;
      864:data<=-16'd18677;
      865:data<=-16'd17528;
      866:data<=-16'd16909;
      867:data<=-16'd16970;
      868:data<=-16'd15673;
      869:data<=-16'd15879;
      870:data<=-16'd16433;
      871:data<=-16'd13991;
      872:data<=-16'd12863;
      873:data<=-16'd13241;
      874:data<=-16'd12539;
      875:data<=-16'd12216;
      876:data<=-16'd11280;
      877:data<=-16'd10229;
      878:data<=-16'd9923;
      879:data<=-16'd8916;
      880:data<=-16'd8671;
      881:data<=-16'd8287;
      882:data<=-16'd7230;
      883:data<=-16'd7909;
      884:data<=-16'd8686;
      885:data<=-16'd9094;
      886:data<=-16'd8358;
      887:data<=-16'd6742;
      888:data<=-16'd8222;
      889:data<=-16'd3850;
      890:data<=16'd8878;
      891:data<=16'd12336;
      892:data<=16'd9257;
      893:data<=16'd11283;
      894:data<=16'd10953;
      895:data<=16'd9248;
      896:data<=16'd10248;
      897:data<=16'd8886;
      898:data<=16'd8843;
      899:data<=16'd9803;
      900:data<=16'd7295;
      901:data<=16'd6390;
      902:data<=16'd6364;
      903:data<=16'd6529;
      904:data<=16'd11632;
      905:data<=16'd15582;
      906:data<=16'd14337;
      907:data<=16'd13496;
      908:data<=16'd13593;
      909:data<=16'd13118;
      910:data<=16'd12463;
      911:data<=16'd11427;
      912:data<=16'd11133;
      913:data<=16'd11662;
      914:data<=16'd11652;
      915:data<=16'd11129;
      916:data<=16'd10402;
      917:data<=16'd9063;
      918:data<=16'd7964;
      919:data<=16'd8457;
      920:data<=16'd8566;
      921:data<=16'd7579;
      922:data<=16'd8019;
      923:data<=16'd8643;
      924:data<=16'd8070;
      925:data<=16'd7307;
      926:data<=16'd6953;
      927:data<=16'd8102;
      928:data<=16'd7413;
      929:data<=16'd5579;
      930:data<=16'd7964;
      931:data<=16'd4187;
      932:data<=-16'd8264;
      933:data<=-16'd11966;
      934:data<=-16'd9784;
      935:data<=-16'd11370;
      936:data<=-16'd10531;
      937:data<=-16'd9461;
      938:data<=-16'd10111;
      939:data<=-16'd8320;
      940:data<=-16'd7920;
      941:data<=-16'd8075;
      942:data<=-16'd7330;
      943:data<=-16'd8103;
      944:data<=-16'd6766;
      945:data<=-16'd5291;
      946:data<=-16'd5598;
      947:data<=-16'd4002;
      948:data<=-16'd3999;
      949:data<=-16'd4673;
      950:data<=-16'd3755;
      951:data<=-16'd5465;
      952:data<=-16'd5206;
      953:data<=-16'd3380;
      954:data<=-16'd8240;
      955:data<=-16'd13564;
      956:data<=-16'd13345;
      957:data<=-16'd11947;
      958:data<=-16'd11032;
      959:data<=-16'd10358;
      960:data<=-16'd10032;
      961:data<=-16'd9884;
      962:data<=-16'd8950;
      963:data<=-16'd7197;
      964:data<=-16'd7010;
      965:data<=-16'd6951;
      966:data<=-16'd6331;
      967:data<=-16'd6825;
      968:data<=-16'd6752;
      969:data<=-16'd7624;
      970:data<=-16'd8076;
      971:data<=-16'd5789;
      972:data<=-16'd6222;
      973:data<=-16'd2282;
      974:data<=16'd10355;
      975:data<=16'd14945;
      976:data<=16'd11985;
      977:data<=16'd12528;
      978:data<=16'd12354;
      979:data<=16'd12099;
      980:data<=16'd12765;
      981:data<=16'd11241;
      982:data<=16'd11039;
      983:data<=16'd10237;
      984:data<=16'd7773;
      985:data<=16'd7603;
      986:data<=16'd7072;
      987:data<=16'd6523;
      988:data<=16'd7268;
      989:data<=16'd7013;
      990:data<=16'd7189;
      991:data<=16'd6764;
      992:data<=16'd6070;
      993:data<=16'd7283;
      994:data<=16'd6846;
      995:data<=16'd6226;
      996:data<=16'd7216;
      997:data<=16'd6382;
      998:data<=16'd6062;
      999:data<=16'd6605;
      1000:data<=16'd5603;
      1001:data<=16'd4883;
      1002:data<=16'd3714;
      1003:data<=16'd3369;
      1004:data<=16'd7192;
      1005:data<=16'd11844;
      1006:data<=16'd13027;
      1007:data<=16'd11662;
      1008:data<=16'd11708;
      1009:data<=16'd12176;
      1010:data<=16'd10554;
      1011:data<=16'd10571;
      1012:data<=16'd10502;
      1013:data<=16'd9030;
      1014:data<=16'd10530;
      1015:data<=16'd6087;
      1016:data<=-16'd6260;
      1017:data<=-16'd11388;
      1018:data<=-16'd10577;
      1019:data<=-16'd10398;
      1020:data<=-16'd8178;
      1021:data<=-16'd7602;
      1022:data<=-16'd8702;
      1023:data<=-16'd7811;
      1024:data<=-16'd7407;
      1025:data<=-16'd6837;
      1026:data<=-16'd5929;
      1027:data<=-16'd5736;
      1028:data<=-16'd4537;
      1029:data<=-16'd4417;
      1030:data<=-16'd5250;
      1031:data<=-16'd4608;
      1032:data<=-16'd4564;
      1033:data<=-16'd5198;
      1034:data<=-16'd5611;
      1035:data<=-16'd5949;
      1036:data<=-16'd5462;
      1037:data<=-16'd5103;
      1038:data<=-16'd4576;
      1039:data<=-16'd4087;
      1040:data<=-16'd4611;
      1041:data<=-16'd3582;
      1042:data<=-16'd2466;
      1043:data<=-16'd3306;
      1044:data<=-16'd3019;
      1045:data<=-16'd2760;
      1046:data<=-16'd3092;
      1047:data<=-16'd1730;
      1048:data<=-16'd698;
      1049:data<=-16'd393;
      1050:data<=-16'd1057;
      1051:data<=-16'd3224;
      1052:data<=-16'd2980;
      1053:data<=-16'd1877;
      1054:data<=-16'd3982;
      1055:data<=-16'd8156;
      1056:data<=-16'd11778;
      1057:data<=-16'd6862;
      1058:data<=16'd6034;
      1059:data<=16'd11403;
      1060:data<=16'd9121;
      1061:data<=16'd9357;
      1062:data<=16'd9617;
      1063:data<=16'd8931;
      1064:data<=16'd9279;
      1065:data<=16'd8426;
      1066:data<=16'd7956;
      1067:data<=16'd7715;
      1068:data<=16'd6115;
      1069:data<=16'd5477;
      1070:data<=16'd4287;
      1071:data<=16'd2690;
      1072:data<=16'd3856;
      1073:data<=16'd4868;
      1074:data<=16'd4831;
      1075:data<=16'd5313;
      1076:data<=16'd4831;
      1077:data<=16'd5422;
      1078:data<=16'd6915;
      1079:data<=16'd5703;
      1080:data<=16'd5015;
      1081:data<=16'd6454;
      1082:data<=16'd6492;
      1083:data<=16'd6067;
      1084:data<=16'd6243;
      1085:data<=16'd5638;
      1086:data<=16'd5492;
      1087:data<=16'd6044;
      1088:data<=16'd5664;
      1089:data<=16'd5316;
      1090:data<=16'd5468;
      1091:data<=16'd4911;
      1092:data<=16'd4804;
      1093:data<=16'd4989;
      1094:data<=16'd4313;
      1095:data<=16'd5121;
      1096:data<=16'd5523;
      1097:data<=16'd4147;
      1098:data<=16'd5755;
      1099:data<=16'd2830;
      1100:data<=-16'd9332;
      1101:data<=-16'd13911;
      1102:data<=-16'd10063;
      1103:data<=-16'd10772;
      1104:data<=-16'd8599;
      1105:data<=-16'd1322;
      1106:data<=16'd564;
      1107:data<=-16'd83;
      1108:data<=16'd644;
      1109:data<=16'd845;
      1110:data<=16'd1607;
      1111:data<=16'd2130;
      1112:data<=16'd1851;
      1113:data<=16'd1492;
      1114:data<=16'd1309;
      1115:data<=16'd2170;
      1116:data<=16'd2035;
      1117:data<=16'd1747;
      1118:data<=16'd3645;
      1119:data<=16'd4043;
      1120:data<=16'd3570;
      1121:data<=16'd4717;
      1122:data<=16'd4476;
      1123:data<=16'd3940;
      1124:data<=16'd4561;
      1125:data<=16'd4472;
      1126:data<=16'd4763;
      1127:data<=16'd5168;
      1128:data<=16'd4487;
      1129:data<=16'd3811;
      1130:data<=16'd3588;
      1131:data<=16'd4040;
      1132:data<=16'd4173;
      1133:data<=16'd3516;
      1134:data<=16'd4137;
      1135:data<=16'd6088;
      1136:data<=16'd6822;
      1137:data<=16'd5136;
      1138:data<=16'd4817;
      1139:data<=16'd6460;
      1140:data<=16'd4511;
      1141:data<=16'd6558;
      1142:data<=16'd18642;
      1143:data<=16'd24410;
      1144:data<=16'd21030;
      1145:data<=16'd21179;
      1146:data<=16'd21014;
      1147:data<=16'd18782;
      1148:data<=16'd19326;
      1149:data<=16'd18571;
      1150:data<=16'd17411;
      1151:data<=16'd18313;
      1152:data<=16'd18713;
      1153:data<=16'd18762;
      1154:data<=16'd15170;
      1155:data<=16'd8605;
      1156:data<=16'd6724;
      1157:data<=16'd7365;
      1158:data<=16'd6551;
      1159:data<=16'd6310;
      1160:data<=16'd6170;
      1161:data<=16'd6017;
      1162:data<=16'd6140;
      1163:data<=16'd5758;
      1164:data<=16'd5914;
      1165:data<=16'd5764;
      1166:data<=16'd4590;
      1167:data<=16'd4698;
      1168:data<=16'd6202;
      1169:data<=16'd6672;
      1170:data<=16'd5497;
      1171:data<=16'd4811;
      1172:data<=16'd5057;
      1173:data<=16'd4648;
      1174:data<=16'd4461;
      1175:data<=16'd4702;
      1176:data<=16'd4105;
      1177:data<=16'd3275;
      1178:data<=16'd2930;
      1179:data<=16'd3466;
      1180:data<=16'd3432;
      1181:data<=16'd2851;
      1182:data<=16'd4466;
      1183:data<=16'd1836;
      1184:data<=-16'd8243;
      1185:data<=-16'd13386;
      1186:data<=-16'd11815;
      1187:data<=-16'd11629;
      1188:data<=-16'd11089;
      1189:data<=-16'd10410;
      1190:data<=-16'd11279;
      1191:data<=-16'd10536;
      1192:data<=-16'd9470;
      1193:data<=-16'd8895;
      1194:data<=-16'd8022;
      1195:data<=-16'd8156;
      1196:data<=-16'd7706;
      1197:data<=-16'd7103;
      1198:data<=-16'd7595;
      1199:data<=-16'd7326;
      1200:data<=-16'd6940;
      1201:data<=-16'd5395;
      1202:data<=-16'd3090;
      1203:data<=-16'd4024;
      1204:data<=-16'd3231;
      1205:data<=16'd2181;
      1206:data<=16'd4654;
      1207:data<=16'd3792;
      1208:data<=16'd3923;
      1209:data<=16'd3997;
      1210:data<=16'd3519;
      1211:data<=16'd3820;
      1212:data<=16'd4607;
      1213:data<=16'd4124;
      1214:data<=16'd2799;
      1215:data<=16'd2720;
      1216:data<=16'd3193;
      1217:data<=16'd3738;
      1218:data<=16'd4607;
      1219:data<=16'd5356;
      1220:data<=16'd6209;
      1221:data<=16'd5174;
      1222:data<=16'd3519;
      1223:data<=16'd3955;
      1224:data<=16'd2205;
      1225:data<=16'd3210;
      1226:data<=16'd14131;
      1227:data<=16'd21652;
      1228:data<=16'd19347;
      1229:data<=16'd17882;
      1230:data<=16'd17741;
      1231:data<=16'd16311;
      1232:data<=16'd16004;
      1233:data<=16'd15054;
      1234:data<=16'd13920;
      1235:data<=16'd14832;
      1236:data<=16'd15547;
      1237:data<=16'd14173;
      1238:data<=16'd12005;
      1239:data<=16'd11200;
      1240:data<=16'd10968;
      1241:data<=16'd10571;
      1242:data<=16'd11097;
      1243:data<=16'd9765;
      1244:data<=16'd6940;
      1245:data<=16'd7512;
      1246:data<=16'd8698;
      1247:data<=16'd7453;
      1248:data<=16'd6821;
      1249:data<=16'd6657;
      1250:data<=16'd5882;
      1251:data<=16'd5767;
      1252:data<=16'd6270;
      1253:data<=16'd6578;
      1254:data<=16'd4989;
      1255:data<=16'd675;
      1256:data<=-16'd3306;
      1257:data<=-16'd4297;
      1258:data<=-16'd4006;
      1259:data<=-16'd4206;
      1260:data<=-16'd3724;
      1261:data<=-16'd3336;
      1262:data<=-16'd4461;
      1263:data<=-16'd4592;
      1264:data<=-16'd3792;
      1265:data<=-16'd3560;
      1266:data<=-16'd1955;
      1267:data<=-16'd2998;
      1268:data<=-16'd11291;
      1269:data<=-16'd18988;
      1270:data<=-16'd19707;
      1271:data<=-16'd18128;
      1272:data<=-16'd17650;
      1273:data<=-16'd17241;
      1274:data<=-16'd16772;
      1275:data<=-16'd15954;
      1276:data<=-16'd14822;
      1277:data<=-16'd15083;
      1278:data<=-16'd15693;
      1279:data<=-16'd14342;
      1280:data<=-16'd13117;
      1281:data<=-16'd13103;
      1282:data<=-16'd12352;
      1283:data<=-16'd11699;
      1284:data<=-16'd11012;
      1285:data<=-16'd9080;
      1286:data<=-16'd8399;
      1287:data<=-16'd9147;
      1288:data<=-16'd9094;
      1289:data<=-16'd8836;
      1290:data<=-16'd8355;
      1291:data<=-16'd7705;
      1292:data<=-16'd7867;
      1293:data<=-16'd7597;
      1294:data<=-16'd7089;
      1295:data<=-16'd7473;
      1296:data<=-16'd7389;
      1297:data<=-16'd7062;
      1298:data<=-16'd6984;
      1299:data<=-16'd6285;
      1300:data<=-16'd5962;
      1301:data<=-16'd5163;
      1302:data<=-16'd3262;
      1303:data<=-16'd3472;
      1304:data<=-16'd3312;
      1305:data<=16'd829;
      1306:data<=16'd4056;
      1307:data<=16'd3974;
      1308:data<=16'd2635;
      1309:data<=16'd3065;
      1310:data<=16'd10857;
      1311:data<=16'd20151;
      1312:data<=16'd20583;
      1313:data<=16'd18310;
      1314:data<=16'd18340;
      1315:data<=16'd16707;
      1316:data<=16'd15485;
      1317:data<=16'd15173;
      1318:data<=16'd14175;
      1319:data<=16'd14560;
      1320:data<=16'd14516;
      1321:data<=16'd13559;
      1322:data<=16'd13294;
      1323:data<=16'd11649;
      1324:data<=16'd9935;
      1325:data<=16'd9687;
      1326:data<=16'd9403;
      1327:data<=16'd9617;
      1328:data<=16'd9320;
      1329:data<=16'd8282;
      1330:data<=16'd8337;
      1331:data<=16'd7923;
      1332:data<=16'd6622;
      1333:data<=16'd5841;
      1334:data<=16'd5658;
      1335:data<=16'd6137;
      1336:data<=16'd6134;
      1337:data<=16'd5683;
      1338:data<=16'd5959;
      1339:data<=16'd6012;
      1340:data<=16'd5259;
      1341:data<=16'd4009;
      1342:data<=16'd3430;
      1343:data<=16'd3339;
      1344:data<=16'd2282;
      1345:data<=16'd2414;
      1346:data<=16'd2576;
      1347:data<=16'd1069;
      1348:data<=16'd1959;
      1349:data<=16'd2144;
      1350:data<=16'd746;
      1351:data<=16'd1316;
      1352:data<=-16'd6041;
      1353:data<=-16'd17532;
      1354:data<=-16'd17655;
      1355:data<=-16'd17699;
      1356:data<=-16'd24283;
      1357:data<=-16'd24914;
      1358:data<=-16'd22492;
      1359:data<=-16'd22221;
      1360:data<=-16'd21182;
      1361:data<=-16'd20615;
      1362:data<=-16'd20043;
      1363:data<=-16'd19811;
      1364:data<=-16'd19934;
      1365:data<=-16'd18055;
      1366:data<=-16'd17317;
      1367:data<=-16'd17373;
      1368:data<=-16'd16362;
      1369:data<=-16'd17356;
      1370:data<=-16'd17588;
      1371:data<=-16'd16134;
      1372:data<=-16'd16587;
      1373:data<=-16'd16616;
      1374:data<=-16'd15453;
      1375:data<=-16'd14352;
      1376:data<=-16'd13406;
      1377:data<=-16'd14029;
      1378:data<=-16'd14098;
      1379:data<=-16'd12834;
      1380:data<=-16'd12648;
      1381:data<=-16'd12801;
      1382:data<=-16'd12625;
      1383:data<=-16'd11392;
      1384:data<=-16'd10126;
      1385:data<=-16'd11194;
      1386:data<=-16'd12079;
      1387:data<=-16'd12222;
      1388:data<=-16'd11768;
      1389:data<=-16'd9931;
      1390:data<=-16'd10428;
      1391:data<=-16'd10543;
      1392:data<=-16'd9171;
      1393:data<=-16'd10226;
      1394:data<=-16'd3583;
      1395:data<=16'd8793;
      1396:data<=16'd9841;
      1397:data<=16'd6657;
      1398:data<=16'd7633;
      1399:data<=16'd6843;
      1400:data<=16'd6314;
      1401:data<=16'd5586;
      1402:data<=16'd3606;
      1403:data<=16'd3551;
      1404:data<=16'd2793;
      1405:data<=16'd5515;
      1406:data<=16'd12041;
      1407:data<=16'd12075;
      1408:data<=16'd9759;
      1409:data<=16'd10131;
      1410:data<=16'd9436;
      1411:data<=16'd9750;
      1412:data<=16'd9591;
      1413:data<=16'd8031;
      1414:data<=16'd8846;
      1415:data<=16'd8596;
      1416:data<=16'd7042;
      1417:data<=16'd6918;
      1418:data<=16'd5685;
      1419:data<=16'd4455;
      1420:data<=16'd4341;
      1421:data<=16'd3956;
      1422:data<=16'd3943;
      1423:data<=16'd3883;
      1424:data<=16'd3682;
      1425:data<=16'd2684;
      1426:data<=16'd1098;
      1427:data<=16'd1530;
      1428:data<=16'd2056;
      1429:data<=16'd1416;
      1430:data<=16'd1184;
      1431:data<=16'd1242;
      1432:data<=16'd2400;
      1433:data<=16'd1877;
      1434:data<=16'd411;
      1435:data<=16'd1688;
      1436:data<=-16'd4504;
      1437:data<=-16'd17161;
      1438:data<=-16'd19423;
      1439:data<=-16'd16246;
      1440:data<=-16'd16625;
      1441:data<=-16'd15576;
      1442:data<=-16'd14622;
      1443:data<=-16'd14783;
      1444:data<=-16'd13570;
      1445:data<=-16'd12663;
      1446:data<=-16'd11975;
      1447:data<=-16'd12236;
      1448:data<=-16'd12518;
      1449:data<=-16'd11106;
      1450:data<=-16'd10853;
      1451:data<=-16'd10722;
      1452:data<=-16'd11072;
      1453:data<=-16'd12743;
      1454:data<=-16'd11165;
      1455:data<=-16'd12185;
      1456:data<=-16'd18616;
      1457:data<=-16'd19667;
      1458:data<=-16'd16970;
      1459:data<=-16'd16681;
      1460:data<=-16'd16257;
      1461:data<=-16'd16005;
      1462:data<=-16'd15541;
      1463:data<=-16'd14349;
      1464:data<=-16'd13982;
      1465:data<=-16'd13251;
      1466:data<=-16'd12551;
      1467:data<=-16'd11797;
      1468:data<=-16'd11242;
      1469:data<=-16'd12167;
      1470:data<=-16'd11840;
      1471:data<=-16'd11324;
      1472:data<=-16'd11151;
      1473:data<=-16'd9544;
      1474:data<=-16'd10517;
      1475:data<=-16'd10392;
      1476:data<=-16'd8241;
      1477:data<=-16'd10607;
      1478:data<=-16'd5306;
      1479:data<=16'd8652;
      1480:data<=16'd11597;
      1481:data<=16'd8666;
      1482:data<=16'd9233;
      1483:data<=16'd7891;
      1484:data<=16'd7465;
      1485:data<=16'd7623;
      1486:data<=16'd5515;
      1487:data<=16'd5027;
      1488:data<=16'd5027;
      1489:data<=16'd5257;
      1490:data<=16'd5940;
      1491:data<=16'd5351;
      1492:data<=16'd5756;
      1493:data<=16'd5159;
      1494:data<=16'd3944;
      1495:data<=16'd5300;
      1496:data<=16'd4602;
      1497:data<=16'd3392;
      1498:data<=16'd4435;
      1499:data<=16'd4156;
      1500:data<=16'd4639;
      1501:data<=16'd4637;
      1502:data<=16'd2927;
      1503:data<=16'd3021;
      1504:data<=16'd1527;
      1505:data<=16'd2531;
      1506:data<=16'd9755;
      1507:data<=16'd12148;
      1508:data<=16'd10287;
      1509:data<=16'd10252;
      1510:data<=16'd9101;
      1511:data<=16'd8669;
      1512:data<=16'd8737;
      1513:data<=16'd7702;
      1514:data<=16'd7830;
      1515:data<=16'd7548;
      1516:data<=16'd7861;
      1517:data<=16'd7900;
      1518:data<=16'd6426;
      1519:data<=16'd7459;
      1520:data<=16'd2285;
      1521:data<=-16'd10584;
      1522:data<=-16'd14290;
      1523:data<=-16'd11580;
      1524:data<=-16'd11386;
      1525:data<=-16'd9718;
      1526:data<=-16'd9276;
      1527:data<=-16'd9812;
      1528:data<=-16'd7973;
      1529:data<=-16'd7935;
      1530:data<=-16'd8079;
      1531:data<=-16'd6913;
      1532:data<=-16'd7107;
      1533:data<=-16'd6569;
      1534:data<=-16'd5692;
      1535:data<=-16'd6426;
      1536:data<=-16'd7269;
      1537:data<=-16'd6824;
      1538:data<=-16'd5827;
      1539:data<=-16'd6431;
      1540:data<=-16'd6487;
      1541:data<=-16'd5263;
      1542:data<=-16'd5829;
      1543:data<=-16'd5389;
      1544:data<=-16'd4303;
      1545:data<=-16'd4757;
      1546:data<=-16'd3130;
      1547:data<=-16'd2209;
      1548:data<=-16'd3001;
      1549:data<=-16'd2196;
      1550:data<=-16'd2402;
      1551:data<=-16'd1682;
      1552:data<=-16'd1099;
      1553:data<=-16'd3453;
      1554:data<=-16'd2393;
      1555:data<=-16'd3542;
      1556:data<=-16'd9776;
      1557:data<=-16'd10331;
      1558:data<=-16'd9864;
      1559:data<=-16'd10196;
      1560:data<=-16'd7953;
      1561:data<=-16'd10047;
      1562:data<=-16'd5567;
      1563:data<=16'd8470;
      1564:data<=16'd11429;
      1565:data<=16'd8366;
      1566:data<=16'd10111;
      1567:data<=16'd9579;
      1568:data<=16'd8396;
      1569:data<=16'd7621;
      1570:data<=16'd6140;
      1571:data<=16'd7339;
      1572:data<=16'd7335;
      1573:data<=16'd6552;
      1574:data<=16'd7661;
      1575:data<=16'd6865;
      1576:data<=16'd6381;
      1577:data<=16'd7189;
      1578:data<=16'd6623;
      1579:data<=16'd6598;
      1580:data<=16'd6845;
      1581:data<=16'd7183;
      1582:data<=16'd7981;
      1583:data<=16'd7608;
      1584:data<=16'd7494;
      1585:data<=16'd7130;
      1586:data<=16'd5476;
      1587:data<=16'd4672;
      1588:data<=16'd4115;
      1589:data<=16'd3682;
      1590:data<=16'd4085;
      1591:data<=16'd4740;
      1592:data<=16'd5300;
      1593:data<=16'd4205;
      1594:data<=16'd3726;
      1595:data<=16'd4895;
      1596:data<=16'd4081;
      1597:data<=16'd4065;
      1598:data<=16'd4563;
      1599:data<=16'd3142;
      1600:data<=16'd4695;
      1601:data<=16'd5009;
      1602:data<=16'd3162;
      1603:data<=16'd5532;
      1604:data<=16'd276;
      1605:data<=-16'd11176;
      1606:data<=-16'd9300;
      1607:data<=-16'd3351;
      1608:data<=-16'd4570;
      1609:data<=-16'd3686;
      1610:data<=-16'd2047;
      1611:data<=-16'd2958;
      1612:data<=-16'd2736;
      1613:data<=-16'd2775;
      1614:data<=-16'd2544;
      1615:data<=-16'd1434;
      1616:data<=-16'd1623;
      1617:data<=-16'd2003;
      1618:data<=-16'd1795;
      1619:data<=-16'd1105;
      1620:data<=-16'd795;
      1621:data<=-16'd1480;
      1622:data<=-16'd1353;
      1623:data<=-16'd1221;
      1624:data<=-16'd1246;
      1625:data<=-16'd599;
      1626:data<=-16'd1199;
      1627:data<=-16'd923;
      1628:data<=16'd484;
      1629:data<=-16'd153;
      1630:data<=-16'd49;
      1631:data<=16'd693;
      1632:data<=16'd329;
      1633:data<=16'd970;
      1634:data<=16'd1151;
      1635:data<=16'd1830;
      1636:data<=16'd3509;
      1637:data<=16'd3062;
      1638:data<=16'd3624;
      1639:data<=16'd4469;
      1640:data<=16'd3682;
      1641:data<=16'd4658;
      1642:data<=16'd3833;
      1643:data<=16'd3177;
      1644:data<=16'd4693;
      1645:data<=16'd1513;
      1646:data<=16'd5406;
      1647:data<=16'd19247;
      1648:data<=16'd21967;
      1649:data<=16'd18762;
      1650:data<=16'd20392;
      1651:data<=16'd18619;
      1652:data<=16'd17547;
      1653:data<=16'd19547;
      1654:data<=16'd19032;
      1655:data<=16'd17823;
      1656:data<=16'd13106;
      1657:data<=16'd7498;
      1658:data<=16'd7729;
      1659:data<=16'd8066;
      1660:data<=16'd7600;
      1661:data<=16'd8522;
      1662:data<=16'd7556;
      1663:data<=16'd6828;
      1664:data<=16'd7050;
      1665:data<=16'd6877;
      1666:data<=16'd7406;
      1667:data<=16'd7124;
      1668:data<=16'd6760;
      1669:data<=16'd7275;
      1670:data<=16'd7579;
      1671:data<=16'd8094;
      1672:data<=16'd7577;
      1673:data<=16'd6902;
      1674:data<=16'd6968;
      1675:data<=16'd6213;
      1676:data<=16'd6542;
      1677:data<=16'd6479;
      1678:data<=16'd5265;
      1679:data<=16'd6217;
      1680:data<=16'd6037;
      1681:data<=16'd5092;
      1682:data<=16'd5641;
      1683:data<=16'd4485;
      1684:data<=16'd4943;
      1685:data<=16'd5829;
      1686:data<=16'd5160;
      1687:data<=16'd8519;
      1688:data<=16'd5072;
      1689:data<=-16'd8094;
      1690:data<=-16'd12108;
      1691:data<=-16'd9988;
      1692:data<=-16'd10910;
      1693:data<=-16'd9221;
      1694:data<=-16'd7950;
      1695:data<=-16'd8526;
      1696:data<=-16'd7873;
      1697:data<=-16'd8436;
      1698:data<=-16'd7887;
      1699:data<=-16'd6678;
      1700:data<=-16'd7530;
      1701:data<=-16'd7309;
      1702:data<=-16'd6402;
      1703:data<=-16'd4993;
      1704:data<=-16'd3773;
      1705:data<=-16'd4285;
      1706:data<=-16'd654;
      1707:data<=16'd4801;
      1708:data<=16'd4693;
      1709:data<=16'd3677;
      1710:data<=16'd4228;
      1711:data<=16'd4463;
      1712:data<=16'd4955;
      1713:data<=16'd4375;
      1714:data<=16'd3802;
      1715:data<=16'd3859;
      1716:data<=16'd3319;
      1717:data<=16'd3133;
      1718:data<=16'd2598;
      1719:data<=16'd3290;
      1720:data<=16'd5016;
      1721:data<=16'd3842;
      1722:data<=16'd3240;
      1723:data<=16'd4202;
      1724:data<=16'd4200;
      1725:data<=16'd4860;
      1726:data<=16'd3613;
      1727:data<=16'd2866;
      1728:data<=16'd3991;
      1729:data<=16'd432;
      1730:data<=16'd3212;
      1731:data<=16'd16108;
      1732:data<=16'd19925;
      1733:data<=16'd17280;
      1734:data<=16'd17858;
      1735:data<=16'd16039;
      1736:data<=16'd15082;
      1737:data<=16'd16264;
      1738:data<=16'd15515;
      1739:data<=16'd15763;
      1740:data<=16'd15477;
      1741:data<=16'd14310;
      1742:data<=16'd13861;
      1743:data<=16'd11967;
      1744:data<=16'd11583;
      1745:data<=16'd11828;
      1746:data<=16'd10261;
      1747:data<=16'd10373;
      1748:data<=16'd10055;
      1749:data<=16'd9370;
      1750:data<=16'd9814;
      1751:data<=16'd8140;
      1752:data<=16'd8134;
      1753:data<=16'd9386;
      1754:data<=16'd8470;
      1755:data<=16'd9427;
      1756:data<=16'd7010;
      1757:data<=16'd67;
      1758:data<=-16'd1509;
      1759:data<=-16'd758;
      1760:data<=-16'd1509;
      1761:data<=-16'd1568;
      1762:data<=-16'd2367;
      1763:data<=-16'd2140;
      1764:data<=-16'd1571;
      1765:data<=-16'd1906;
      1766:data<=-16'd1048;
      1767:data<=-16'd1739;
      1768:data<=-16'd2494;
      1769:data<=-16'd1717;
      1770:data<=-16'd1343;
      1771:data<=16'd1380;
      1772:data<=-16'd1478;
      1773:data<=-16'd13189;
      1774:data<=-16'd17805;
      1775:data<=-16'd15828;
      1776:data<=-16'd16205;
      1777:data<=-16'd15423;
      1778:data<=-16'd14933;
      1779:data<=-16'd14879;
      1780:data<=-16'd12983;
      1781:data<=-16'd13101;
      1782:data<=-16'd13277;
      1783:data<=-16'd11847;
      1784:data<=-16'd11544;
      1785:data<=-16'd11605;
      1786:data<=-16'd11306;
      1787:data<=-16'd9747;
      1788:data<=-16'd8804;
      1789:data<=-16'd9714;
      1790:data<=-16'd8495;
      1791:data<=-16'd7791;
      1792:data<=-16'd8809;
      1793:data<=-16'd7846;
      1794:data<=-16'd8064;
      1795:data<=-16'd8322;
      1796:data<=-16'd7062;
      1797:data<=-16'd7564;
      1798:data<=-16'd6605;
      1799:data<=-16'd5791;
      1800:data<=-16'd6942;
      1801:data<=-16'd5818;
      1802:data<=-16'd5927;
      1803:data<=-16'd5441;
      1804:data<=-16'd2890;
      1805:data<=-16'd4742;
      1806:data<=-16'd2634;
      1807:data<=16'd4494;
      1808:data<=16'd5195;
      1809:data<=16'd4560;
      1810:data<=16'd4569;
      1811:data<=16'd3388;
      1812:data<=16'd4303;
      1813:data<=16'd1770;
      1814:data<=16'd3318;
      1815:data<=16'd15484;
      1816:data<=16'd20528;
      1817:data<=16'd17983;
      1818:data<=16'd18017;
      1819:data<=16'd16728;
      1820:data<=16'd16543;
      1821:data<=16'd17097;
      1822:data<=16'd15091;
      1823:data<=16'd15502;
      1824:data<=16'd15103;
      1825:data<=16'd12891;
      1826:data<=16'd13505;
      1827:data<=16'd12878;
      1828:data<=16'd11488;
      1829:data<=16'd11470;
      1830:data<=16'd10087;
      1831:data<=16'd9221;
      1832:data<=16'd8704;
      1833:data<=16'd7843;
      1834:data<=16'd8153;
      1835:data<=16'd7812;
      1836:data<=16'd7949;
      1837:data<=16'd8495;
      1838:data<=16'd7483;
      1839:data<=16'd7588;
      1840:data<=16'd7444;
      1841:data<=16'd5792;
      1842:data<=16'd5227;
      1843:data<=16'd4678;
      1844:data<=16'd4513;
      1845:data<=16'd4508;
      1846:data<=16'd3630;
      1847:data<=16'd4144;
      1848:data<=16'd3959;
      1849:data<=16'd3207;
      1850:data<=16'd3824;
      1851:data<=16'd2423;
      1852:data<=16'd1817;
      1853:data<=16'd2429;
      1854:data<=16'd2011;
      1855:data<=16'd5375;
      1856:data<=16'd1325;
      1857:data<=-16'd16540;
      1858:data<=-16'd25575;
      1859:data<=-16'd22319;
      1860:data<=-16'd21713;
      1861:data<=-16'd21312;
      1862:data<=-16'd19725;
      1863:data<=-16'd19271;
      1864:data<=-16'd17799;
      1865:data<=-16'd17834;
      1866:data<=-16'd18469;
      1867:data<=-16'd17412;
      1868:data<=-16'd16747;
      1869:data<=-16'd15643;
      1870:data<=-16'd14542;
      1871:data<=-16'd14064;
      1872:data<=-16'd13047;
      1873:data<=-16'd12910;
      1874:data<=-16'd12736;
      1875:data<=-16'd12181;
      1876:data<=-16'd12643;
      1877:data<=-16'd12311;
      1878:data<=-16'd11621;
      1879:data<=-16'd11095;
      1880:data<=-16'd10226;
      1881:data<=-16'd10558;
      1882:data<=-16'd10238;
      1883:data<=-16'd9175;
      1884:data<=-16'd9286;
      1885:data<=-16'd8818;
      1886:data<=-16'd8998;
      1887:data<=-16'd9256;
      1888:data<=-16'd8106;
      1889:data<=-16'd9268;
      1890:data<=-16'd10025;
      1891:data<=-16'd8649;
      1892:data<=-16'd8903;
      1893:data<=-16'd7859;
      1894:data<=-16'd6857;
      1895:data<=-16'd7835;
      1896:data<=-16'd6928;
      1897:data<=-16'd8081;
      1898:data<=-16'd6830;
      1899:data<=16'd4431;
      1900:data<=16'd11724;
      1901:data<=16'd9776;
      1902:data<=16'd9118;
      1903:data<=16'd8793;
      1904:data<=16'd6435;
      1905:data<=16'd4435;
      1906:data<=16'd5494;
      1907:data<=16'd11395;
      1908:data<=16'd14402;
      1909:data<=16'd11941;
      1910:data<=16'd11411;
      1911:data<=16'd11420;
      1912:data<=16'd10308;
      1913:data<=16'd10557;
      1914:data<=16'd9647;
      1915:data<=16'd8143;
      1916:data<=16'd8423;
      1917:data<=16'd8846;
      1918:data<=16'd8366;
      1919:data<=16'd6758;
      1920:data<=16'd5103;
      1921:data<=16'd4243;
      1922:data<=16'd3712;
      1923:data<=16'd4081;
      1924:data<=16'd3976;
      1925:data<=16'd2916;
      1926:data<=16'd2769;
      1927:data<=16'd2591;
      1928:data<=16'd2212;
      1929:data<=16'd1927;
      1930:data<=16'd1328;
      1931:data<=16'd1964;
      1932:data<=16'd2108;
      1933:data<=16'd989;
      1934:data<=16'd1233;
      1935:data<=16'd1074;
      1936:data<=16'd368;
      1937:data<=-16'd284;
      1938:data<=-16'd2049;
      1939:data<=-16'd805;
      1940:data<=-16'd1128;
      1941:data<=-16'd11097;
      1942:data<=-16'd19478;
      1943:data<=-16'd18747;
      1944:data<=-16'd17338;
      1945:data<=-16'd16812;
      1946:data<=-16'd15343;
      1947:data<=-16'd14844;
      1948:data<=-16'd14530;
      1949:data<=-16'd14113;
      1950:data<=-16'd13896;
      1951:data<=-16'd13006;
      1952:data<=-16'd12334;
      1953:data<=-16'd13550;
      1954:data<=-16'd15147;
      1955:data<=-16'd13998;
      1956:data<=-16'd14187;
      1957:data<=-16'd19500;
      1958:data<=-16'd22522;
      1959:data<=-16'd20996;
      1960:data<=-16'd20312;
      1961:data<=-16'd19334;
      1962:data<=-16'd17881;
      1963:data<=-16'd17552;
      1964:data<=-16'd16451;
      1965:data<=-16'd15678;
      1966:data<=-16'd15622;
      1967:data<=-16'd15000;
      1968:data<=-16'd14418;
      1969:data<=-16'd13126;
      1970:data<=-16'd12806;
      1971:data<=-16'd13910;
      1972:data<=-16'd13174;
      1973:data<=-16'd12988;
      1974:data<=-16'd13696;
      1975:data<=-16'd12160;
      1976:data<=-16'd11455;
      1977:data<=-16'd11597;
      1978:data<=-16'd10524;
      1979:data<=-16'd10122;
      1980:data<=-16'd9451;
      1981:data<=-16'd9406;
      1982:data<=-16'd8577;
      1983:data<=-16'd36;
      1984:data<=16'd9781;
      1985:data<=16'd11097;
      1986:data<=16'd9078;
      1987:data<=16'd7829;
      1988:data<=16'd6208;
      1989:data<=16'd5735;
      1990:data<=16'd5908;
      1991:data<=16'd6017;
      1992:data<=16'd6361;
      1993:data<=16'd5830;
      1994:data<=16'd5524;
      1995:data<=16'd6250;
      1996:data<=16'd6332;
      1997:data<=16'd5926;
      1998:data<=16'd6078;
      1999:data<=16'd6172;
      2000:data<=16'd5466;
      2001:data<=16'd5115;
      2002:data<=16'd5891;
      2003:data<=16'd5862;
      2004:data<=16'd4470;
      2005:data<=16'd3130;
      2006:data<=16'd3501;
      2007:data<=16'd7779;
      2008:data<=16'd12437;
      2009:data<=16'd12375;
      2010:data<=16'd11077;
      2011:data<=16'd11104;
      2012:data<=16'd10698;
      2013:data<=16'd10417;
      2014:data<=16'd9592;
      2015:data<=16'd9250;
      2016:data<=16'd10514;
      2017:data<=16'd9615;
      2018:data<=16'd8592;
      2019:data<=16'd9570;
      2020:data<=16'd8055;
      2021:data<=16'd5974;
      2022:data<=16'd5483;
      2023:data<=16'd5403;
      2024:data<=16'd5673;
      2025:data<=-16'd832;
      2026:data<=-16'd11576;
      2027:data<=-16'd13069;
      2028:data<=-16'd10363;
      2029:data<=-16'd10727;
      2030:data<=-16'd9526;
      2031:data<=-16'd8853;
      2032:data<=-16'd9418;
      2033:data<=-16'd8598;
      2034:data<=-16'd8837;
      2035:data<=-16'd8249;
      2036:data<=-16'd6496;
      2037:data<=-16'd7409;
      2038:data<=-16'd8943;
      2039:data<=-16'd8918;
      2040:data<=-16'd8208;
      2041:data<=-16'd8062;
      2042:data<=-16'd8252;
      2043:data<=-16'd6895;
      2044:data<=-16'd6273;
      2045:data<=-16'd6821;
      2046:data<=-16'd5492;
      2047:data<=-16'd4575;
      2048:data<=-16'd4728;
      2049:data<=-16'd4402;
      2050:data<=-16'd4670;
      2051:data<=-16'd4338;
      2052:data<=-16'd3641;
      2053:data<=-16'd4026;
      2054:data<=-16'd4886;
      2055:data<=-16'd5222;
      2056:data<=-16'd4135;
      2057:data<=-16'd7116;
      2058:data<=-16'd13975;
      2059:data<=-16'd13937;
      2060:data<=-16'd11022;
      2061:data<=-16'd11418;
      2062:data<=-16'd10067;
      2063:data<=-16'd9966;
      2064:data<=-16'd10219;
      2065:data<=-16'd8169;
      2066:data<=-16'd9154;
      2067:data<=-16'd3868;
      2068:data<=16'd9086;
      2069:data<=16'd12498;
      2070:data<=16'd9703;
      2071:data<=16'd9204;
      2072:data<=16'd7332;
      2073:data<=16'd6326;
      2074:data<=16'd6423;
      2075:data<=16'd6153;
      2076:data<=16'd7189;
      2077:data<=16'd6684;
      2078:data<=16'd5727;
      2079:data<=16'd6613;
      2080:data<=16'd6839;
      2081:data<=16'd7031;
      2082:data<=16'd7736;
      2083:data<=16'd8049;
      2084:data<=16'd7837;
      2085:data<=16'd7366;
      2086:data<=16'd7743;
      2087:data<=16'd6579;
      2088:data<=16'd4372;
      2089:data<=16'd4689;
      2090:data<=16'd4507;
      2091:data<=16'd3896;
      2092:data<=16'd4757;
      2093:data<=16'd4338;
      2094:data<=16'd4504;
      2095:data<=16'd5247;
      2096:data<=16'd4416;
      2097:data<=16'd4168;
      2098:data<=16'd3718;
      2099:data<=16'd4332;
      2100:data<=16'd5738;
      2101:data<=16'd4129;
      2102:data<=16'd4297;
      2103:data<=16'd4884;
      2104:data<=16'd2362;
      2105:data<=16'd3022;
      2106:data<=16'd2546;
      2107:data<=16'd3133;
      2108:data<=16'd12046;
      2109:data<=16'd9324;
      2110:data<=-16'd5970;
      2111:data<=-16'd8599;
      2112:data<=-16'd5116;
      2113:data<=-16'd6546;
      2114:data<=-16'd5548;
      2115:data<=-16'd4780;
      2116:data<=-16'd5332;
      2117:data<=-16'd4115;
      2118:data<=-16'd3952;
      2119:data<=-16'd3592;
      2120:data<=-16'd3868;
      2121:data<=-16'd5965;
      2122:data<=-16'd5846;
      2123:data<=-16'd5245;
      2124:data<=-16'd5507;
      2125:data<=-16'd4757;
      2126:data<=-16'd4648;
      2127:data<=-16'd4432;
      2128:data<=-16'd3553;
      2129:data<=-16'd3507;
      2130:data<=-16'd3195;
      2131:data<=-16'd2908;
      2132:data<=-16'd3015;
      2133:data<=-16'd2881;
      2134:data<=-16'd2984;
      2135:data<=-16'd2414;
      2136:data<=-16'd1856;
      2137:data<=-16'd2634;
      2138:data<=-16'd3339;
      2139:data<=-16'd3381;
      2140:data<=-16'd2964;
      2141:data<=-16'd3180;
      2142:data<=-16'd3486;
      2143:data<=-16'd2017;
      2144:data<=-16'd1932;
      2145:data<=-16'd2402;
      2146:data<=-16'd638;
      2147:data<=-16'd1180;
      2148:data<=-16'd1239;
      2149:data<=16'd491;
      2150:data<=-16'd1885;
      2151:data<=16'd2645;
      2152:data<=16'd16415;
      2153:data<=16'd19919;
      2154:data<=16'd15391;
      2155:data<=16'd15541;
      2156:data<=16'd16026;
      2157:data<=16'd12942;
      2158:data<=16'd7632;
      2159:data<=16'd4589;
      2160:data<=16'd6185;
      2161:data<=16'd6214;
      2162:data<=16'd5250;
      2163:data<=16'd6159;
      2164:data<=16'd5655;
      2165:data<=16'd5940;
      2166:data<=16'd6731;
      2167:data<=16'd5651;
      2168:data<=16'd6169;
      2169:data<=16'd6640;
      2170:data<=16'd6478;
      2171:data<=16'd7979;
      2172:data<=16'd7780;
      2173:data<=16'd7030;
      2174:data<=16'd7398;
      2175:data<=16'd6717;
      2176:data<=16'd6963;
      2177:data<=16'd7239;
      2178:data<=16'd6463;
      2179:data<=16'd6663;
      2180:data<=16'd5977;
      2181:data<=16'd5400;
      2182:data<=16'd6182;
      2183:data<=16'd6238;
      2184:data<=16'd6686;
      2185:data<=16'd6449;
      2186:data<=16'd5397;
      2187:data<=16'd5899;
      2188:data<=16'd6287;
      2189:data<=16'd7239;
      2190:data<=16'd7354;
      2191:data<=16'd5953;
      2192:data<=16'd7885;
      2193:data<=16'd3779;
      2194:data<=-16'd9262;
      2195:data<=-16'd12577;
      2196:data<=-16'd8645;
      2197:data<=-16'd9958;
      2198:data<=-16'd9764;
      2199:data<=-16'd8258;
      2200:data<=-16'd9564;
      2201:data<=-16'd8787;
      2202:data<=-16'd7935;
      2203:data<=-16'd8390;
      2204:data<=-16'd6155;
      2205:data<=-16'd4266;
      2206:data<=-16'd5221;
      2207:data<=-16'd3727;
      2208:data<=16'd1820;
      2209:data<=16'd4657;
      2210:data<=16'd3486;
      2211:data<=16'd3621;
      2212:data<=16'd3899;
      2213:data<=16'd3263;
      2214:data<=16'd3504;
      2215:data<=16'd2370;
      2216:data<=16'd1676;
      2217:data<=16'd3018;
      2218:data<=16'd2564;
      2219:data<=16'd1747;
      2220:data<=16'd2323;
      2221:data<=16'd3068;
      2222:data<=16'd4225;
      2223:data<=16'd4610;
      2224:data<=16'd4689;
      2225:data<=16'd4223;
      2226:data<=16'd2552;
      2227:data<=16'd3277;
      2228:data<=16'd4032;
      2229:data<=16'd3142;
      2230:data<=16'd4466;
      2231:data<=16'd4040;
      2232:data<=16'd2517;
      2233:data<=16'd3190;
      2234:data<=16'd1594;
      2235:data<=16'd5921;
      2236:data<=16'd18484;
      2237:data<=16'd22213;
      2238:data<=16'd19252;
      2239:data<=16'd19970;
      2240:data<=16'd19397;
      2241:data<=16'd17834;
      2242:data<=16'd17699;
      2243:data<=16'd16660;
      2244:data<=16'd16231;
      2245:data<=16'd15641;
      2246:data<=16'd14060;
      2247:data<=16'd13499;
      2248:data<=16'd13320;
      2249:data<=16'd13382;
      2250:data<=16'd13379;
      2251:data<=16'd12684;
      2252:data<=16'd12358;
      2253:data<=16'd11731;
      2254:data<=16'd10887;
      2255:data<=16'd11394;
      2256:data<=16'd12455;
      2257:data<=16'd10812;
      2258:data<=16'd5277;
      2259:data<=16'd1674;
      2260:data<=16'd2243;
      2261:data<=16'd1970;
      2262:data<=16'd1588;
      2263:data<=16'd1739;
      2264:data<=16'd629;
      2265:data<=16'd842;
      2266:data<=16'd905;
      2267:data<=16'd420;
      2268:data<=16'd1698;
      2269:data<=16'd796;
      2270:data<=-16'd443;
      2271:data<=16'd829;
      2272:data<=16'd898;
      2273:data<=16'd1744;
      2274:data<=16'd1718;
      2275:data<=16'd62;
      2276:data<=16'd2460;
      2277:data<=-16'd1732;
      2278:data<=-16'd14929;
      2279:data<=-16'd18475;
      2280:data<=-16'd15317;
      2281:data<=-16'd15808;
      2282:data<=-16'd14536;
      2283:data<=-16'd13379;
      2284:data<=-16'd14286;
      2285:data<=-16'd13270;
      2286:data<=-16'd13174;
      2287:data<=-16'd13370;
      2288:data<=-16'd11039;
      2289:data<=-16'd9330;
      2290:data<=-16'd9329;
      2291:data<=-16'd9708;
      2292:data<=-16'd9483;
      2293:data<=-16'd8878;
      2294:data<=-16'd9145;
      2295:data<=-16'd9109;
      2296:data<=-16'd8375;
      2297:data<=-16'd7853;
      2298:data<=-16'd7588;
      2299:data<=-16'd8234;
      2300:data<=-16'd8337;
      2301:data<=-16'd7265;
      2302:data<=-16'd7595;
      2303:data<=-16'd8401;
      2304:data<=-16'd7115;
      2305:data<=-16'd5002;
      2306:data<=-16'd4628;
      2307:data<=-16'd3513;
      2308:data<=16'd1830;
      2309:data<=16'd5104;
      2310:data<=16'd3515;
      2311:data<=16'd4052;
      2312:data<=16'd4349;
      2313:data<=16'd2660;
      2314:data<=16'd3979;
      2315:data<=16'd3798;
      2316:data<=16'd2326;
      2317:data<=16'd3016;
      2318:data<=16'd1139;
      2319:data<=16'd4802;
      2320:data<=16'd16827;
      2321:data<=16'd20782;
      2322:data<=16'd18580;
      2323:data<=16'd19300;
      2324:data<=16'd18167;
      2325:data<=16'd17164;
      2326:data<=16'd17599;
      2327:data<=16'd16090;
      2328:data<=16'd15920;
      2329:data<=16'd15350;
      2330:data<=16'd13306;
      2331:data<=16'd13910;
      2332:data<=16'd13529;
      2333:data<=16'd11785;
      2334:data<=16'd12251;
      2335:data<=16'd11403;
      2336:data<=16'd9791;
      2337:data<=16'd10349;
      2338:data<=16'd10320;
      2339:data<=16'd9850;
      2340:data<=16'd10554;
      2341:data<=16'd10370;
      2342:data<=16'd9124;
      2343:data<=16'd8810;
      2344:data<=16'd8748;
      2345:data<=16'd7790;
      2346:data<=16'd7053;
      2347:data<=16'd6405;
      2348:data<=16'd5876;
      2349:data<=16'd5943;
      2350:data<=16'd4516;
      2351:data<=16'd3720;
      2352:data<=16'd5231;
      2353:data<=16'd4250;
      2354:data<=16'd2913;
      2355:data<=16'd3985;
      2356:data<=16'd3759;
      2357:data<=16'd3136;
      2358:data<=-16'd299;
      2359:data<=-16'd5524;
      2360:data<=-16'd4112;
      2361:data<=-16'd6837;
      2362:data<=-16'd19387;
      2363:data<=-16'd23813;
      2364:data<=-16'd20876;
      2365:data<=-16'd21120;
      2366:data<=-16'd20627;
      2367:data<=-16'd20148;
      2368:data<=-16'd20221;
      2369:data<=-16'd18738;
      2370:data<=-16'd18609;
      2371:data<=-16'd16897;
      2372:data<=-16'd13829;
      2373:data<=-16'd13641;
      2374:data<=-16'd13006;
      2375:data<=-16'd12683;
      2376:data<=-16'd13411;
      2377:data<=-16'd11771;
      2378:data<=-16'd11321;
      2379:data<=-16'd12287;
      2380:data<=-16'd11215;
      2381:data<=-16'd10375;
      2382:data<=-16'd10119;
      2383:data<=-16'd9919;
      2384:data<=-16'd10208;
      2385:data<=-16'd9840;
      2386:data<=-16'd9908;
      2387:data<=-16'd10272;
      2388:data<=-16'd9056;
      2389:data<=-16'd7235;
      2390:data<=-16'd6449;
      2391:data<=-16'd6557;
      2392:data<=-16'd5767;
      2393:data<=-16'd5143;
      2394:data<=-16'd5858;
      2395:data<=-16'd5206;
      2396:data<=-16'd4754;
      2397:data<=-16'd4963;
      2398:data<=-16'd3535;
      2399:data<=-16'd4385;
      2400:data<=-16'd5139;
      2401:data<=-16'd3571;
      2402:data<=-16'd5641;
      2403:data<=-16'd2513;
      2404:data<=16'd10047;
      2405:data<=16'd15652;
      2406:data<=16'd13571;
      2407:data<=16'd13676;
      2408:data<=16'd15415;
      2409:data<=16'd18080;
      2410:data<=16'd19073;
      2411:data<=16'd17461;
      2412:data<=16'd17074;
      2413:data<=16'd16322;
      2414:data<=16'd15191;
      2415:data<=16'd15336;
      2416:data<=16'd14675;
      2417:data<=16'd14037;
      2418:data<=16'd13668;
      2419:data<=16'd13124;
      2420:data<=16'd13104;
      2421:data<=16'd11809;
      2422:data<=16'd10554;
      2423:data<=16'd10314;
      2424:data<=16'd9391;
      2425:data<=16'd9395;
      2426:data<=16'd9163;
      2427:data<=16'd8005;
      2428:data<=16'd8155;
      2429:data<=16'd7424;
      2430:data<=16'd6824;
      2431:data<=16'd7535;
      2432:data<=16'd6067;
      2433:data<=16'd4713;
      2434:data<=16'd4698;
      2435:data<=16'd4100;
      2436:data<=16'd4473;
      2437:data<=16'd4103;
      2438:data<=16'd2408;
      2439:data<=16'd1146;
      2440:data<=-16'd123;
      2441:data<=16'd578;
      2442:data<=16'd719;
      2443:data<=-16'd902;
      2444:data<=16'd869;
      2445:data<=-16'd1941;
      2446:data<=-16'd13581;
      2447:data<=-16'd19646;
      2448:data<=-16'd17963;
      2449:data<=-16'd16772;
      2450:data<=-16'd16134;
      2451:data<=-16'd16204;
      2452:data<=-16'd16336;
      2453:data<=-16'd14879;
      2454:data<=-16'd14583;
      2455:data<=-16'd15875;
      2456:data<=-16'd15967;
      2457:data<=-16'd15023;
      2458:data<=-16'd16807;
      2459:data<=-16'd20864;
      2460:data<=-16'd21387;
      2461:data<=-16'd19628;
      2462:data<=-16'd19399;
      2463:data<=-16'd18544;
      2464:data<=-16'd17475;
      2465:data<=-16'd17094;
      2466:data<=-16'd16402;
      2467:data<=-16'd16759;
      2468:data<=-16'd16766;
      2469:data<=-16'd15575;
      2470:data<=-16'd15048;
      2471:data<=-16'd14728;
      2472:data<=-16'd15438;
      2473:data<=-16'd16035;
      2474:data<=-16'd14411;
      2475:data<=-16'd13797;
      2476:data<=-16'd13694;
      2477:data<=-16'd12372;
      2478:data<=-16'd12055;
      2479:data<=-16'd11327;
      2480:data<=-16'd10470;
      2481:data<=-16'd10370;
      2482:data<=-16'd8745;
      2483:data<=-16'd8404;
      2484:data<=-16'd9021;
      2485:data<=-16'd8437;
      2486:data<=-16'd9915;
      2487:data<=-16'd6717;
      2488:data<=16'd4247;
      2489:data<=16'd9209;
      2490:data<=16'd7245;
      2491:data<=16'd7244;
      2492:data<=16'd7222;
      2493:data<=16'd6733;
      2494:data<=16'd7544;
      2495:data<=16'd7450;
      2496:data<=16'd7115;
      2497:data<=16'd7348;
      2498:data<=16'd7162;
      2499:data<=16'd6590;
      2500:data<=16'd5789;
      2501:data<=16'd5597;
      2502:data<=16'd5976;
      2503:data<=16'd6112;
      2504:data<=16'd6132;
      2505:data<=16'd5463;
      2506:data<=16'd3964;
      2507:data<=16'd3072;
      2508:data<=16'd4998;
      2509:data<=16'd9083;
      2510:data<=16'd10320;
      2511:data<=16'd9019;
      2512:data<=16'd9132;
      2513:data<=16'd8710;
      2514:data<=16'd7720;
      2515:data<=16'd8025;
      2516:data<=16'd7476;
      2517:data<=16'd6843;
      2518:data<=16'd6798;
      2519:data<=16'd6065;
      2520:data<=16'd6184;
      2521:data<=16'd5747;
      2522:data<=16'd3903;
      2523:data<=16'd2986;
      2524:data<=16'd2196;
      2525:data<=16'd2378;
      2526:data<=16'd2984;
      2527:data<=16'd1996;
      2528:data<=16'd3327;
      2529:data<=16'd1842;
      2530:data<=-16'd8925;
      2531:data<=-16'd16154;
      2532:data<=-16'd14537;
      2533:data<=-16'd13949;
      2534:data<=-16'd14122;
      2535:data<=-16'd12907;
      2536:data<=-16'd12743;
      2537:data<=-16'd12105;
      2538:data<=-16'd11861;
      2539:data<=-16'd13076;
      2540:data<=-16'd13009;
      2541:data<=-16'd12031;
      2542:data<=-16'd11706;
      2543:data<=-16'd11817;
      2544:data<=-16'd11715;
      2545:data<=-16'd10921;
      2546:data<=-16'd10477;
      2547:data<=-16'd10425;
      2548:data<=-16'd9740;
      2549:data<=-16'd8933;
      2550:data<=-16'd8246;
      2551:data<=-16'd8040;
      2552:data<=-16'd8533;
      2553:data<=-16'd7967;
      2554:data<=-16'd6592;
      2555:data<=-16'd7319;
      2556:data<=-16'd8992;
      2557:data<=-16'd8150;
      2558:data<=-16'd8505;
      2559:data<=-16'd13157;
      2560:data<=-16'd14789;
      2561:data<=-16'd12355;
      2562:data<=-16'd12510;
      2563:data<=-16'd12002;
      2564:data<=-16'd9426;
      2565:data<=-16'd9383;
      2566:data<=-16'd9198;
      2567:data<=-16'd8737;
      2568:data<=-16'd9270;
      2569:data<=-16'd7859;
      2570:data<=-16'd7838;
      2571:data<=-16'd6331;
      2572:data<=16'd2984;
      2573:data<=16'd9608;
      2574:data<=16'd8872;
      2575:data<=16'd8962;
      2576:data<=16'd8884;
      2577:data<=16'd7865;
      2578:data<=16'd8539;
      2579:data<=16'd8432;
      2580:data<=16'd8205;
      2581:data<=16'd8395;
      2582:data<=16'd7283;
      2583:data<=16'd7348;
      2584:data<=16'd8275;
      2585:data<=16'd7665;
      2586:data<=16'd7359;
      2587:data<=16'd8147;
      2588:data<=16'd8082;
      2589:data<=16'd6440;
      2590:data<=16'd5283;
      2591:data<=16'd5457;
      2592:data<=16'd4842;
      2593:data<=16'd4416;
      2594:data<=16'd5321;
      2595:data<=16'd5190;
      2596:data<=16'd4534;
      2597:data<=16'd4720;
      2598:data<=16'd4916;
      2599:data<=16'd4899;
      2600:data<=16'd4487;
      2601:data<=16'd4391;
      2602:data<=16'd4569;
      2603:data<=16'd4170;
      2604:data<=16'd4607;
      2605:data<=16'd4452;
      2606:data<=16'd2217;
      2607:data<=16'd1162;
      2608:data<=16'd2493;
      2609:data<=16'd6103;
      2610:data<=16'd9209;
      2611:data<=16'd7909;
      2612:data<=16'd7641;
      2613:data<=16'd7363;
      2614:data<=-16'd2135;
      2615:data<=-16'd11550;
      2616:data<=-16'd11013;
      2617:data<=-16'd9019;
      2618:data<=-16'd9053;
      2619:data<=-16'd8513;
      2620:data<=-16'd8408;
      2621:data<=-16'd7962;
      2622:data<=-16'd7846;
      2623:data<=-16'd8693;
      2624:data<=-16'd8768;
      2625:data<=-16'd8786;
      2626:data<=-16'd8646;
      2627:data<=-16'd7993;
      2628:data<=-16'd7853;
      2629:data<=-16'd7529;
      2630:data<=-16'd7341;
      2631:data<=-16'd7247;
      2632:data<=-16'd6457;
      2633:data<=-16'd6387;
      2634:data<=-16'd6203;
      2635:data<=-16'd5125;
      2636:data<=-16'd4757;
      2637:data<=-16'd4384;
      2638:data<=-16'd4231;
      2639:data<=-16'd5086;
      2640:data<=-16'd5466;
      2641:data<=-16'd5266;
      2642:data<=-16'd4707;
      2643:data<=-16'd4422;
      2644:data<=-16'd4777;
      2645:data<=-16'd4102;
      2646:data<=-16'd3662;
      2647:data<=-16'd3829;
      2648:data<=-16'd2728;
      2649:data<=-16'd2500;
      2650:data<=-16'd2461;
      2651:data<=-16'd1230;
      2652:data<=-16'd1434;
      2653:data<=-16'd1093;
      2654:data<=-16'd883;
      2655:data<=-16'd1765;
      2656:data<=16'd5049;
      2657:data<=16'd15215;
      2658:data<=16'd14715;
      2659:data<=16'd9065;
      2660:data<=16'd7183;
      2661:data<=16'd6651;
      2662:data<=16'd6731;
      2663:data<=16'd7191;
      2664:data<=16'd6884;
      2665:data<=16'd6860;
      2666:data<=16'd6810;
      2667:data<=16'd6833;
      2668:data<=16'd7312;
      2669:data<=16'd7189;
      2670:data<=16'd7100;
      2671:data<=16'd7448;
      2672:data<=16'd6774;
      2673:data<=16'd5241;
      2674:data<=16'd4786;
      2675:data<=16'd5245;
      2676:data<=16'd4636;
      2677:data<=16'd3944;
      2678:data<=16'd4363;
      2679:data<=16'd4281;
      2680:data<=16'd4140;
      2681:data<=16'd4238;
      2682:data<=16'd3568;
      2683:data<=16'd3855;
      2684:data<=16'd4760;
      2685:data<=16'd4501;
      2686:data<=16'd4024;
      2687:data<=16'd3600;
      2688:data<=16'd4067;
      2689:data<=16'd4884;
      2690:data<=16'd3776;
      2691:data<=16'd3137;
      2692:data<=16'd3149;
      2693:data<=16'd2341;
      2694:data<=16'd3392;
      2695:data<=16'd3698;
      2696:data<=16'd3022;
      2697:data<=16'd4164;
      2698:data<=-16'd2020;
      2699:data<=-16'd13558;
      2700:data<=-16'd15312;
      2701:data<=-16'd12478;
      2702:data<=-16'd13118;
      2703:data<=-16'd12264;
      2704:data<=-16'd11483;
      2705:data<=-16'd11408;
      2706:data<=-16'd9075;
      2707:data<=-16'd8185;
      2708:data<=-16'd7447;
      2709:data<=-16'd3334;
      2710:data<=-16'd99;
      2711:data<=16'd65;
      2712:data<=-16'd487;
      2713:data<=-16'd385;
      2714:data<=-16'd8;
      2715:data<=-16'd150;
      2716:data<=-16'd282;
      2717:data<=-16'd293;
      2718:data<=-16'd103;
      2719:data<=16'd737;
      2720:data<=16'd785;
      2721:data<=16'd183;
      2722:data<=16'd928;
      2723:data<=16'd2626;
      2724:data<=16'd3463;
      2725:data<=16'd3046;
      2726:data<=16'd2910;
      2727:data<=16'd2978;
      2728:data<=16'd2776;
      2729:data<=16'd3592;
      2730:data<=16'd3334;
      2731:data<=16'd2366;
      2732:data<=16'd3879;
      2733:data<=16'd3929;
      2734:data<=16'd2775;
      2735:data<=16'd3762;
      2736:data<=16'd3239;
      2737:data<=16'd3521;
      2738:data<=16'd4047;
      2739:data<=16'd1710;
      2740:data<=16'd9128;
      2741:data<=16'd22615;
      2742:data<=16'd23581;
      2743:data<=16'd20635;
      2744:data<=16'd21778;
      2745:data<=16'd19657;
      2746:data<=16'd18553;
      2747:data<=16'd19478;
      2748:data<=16'd17829;
      2749:data<=16'd17168;
      2750:data<=16'd16833;
      2751:data<=16'd15609;
      2752:data<=16'd15656;
      2753:data<=16'd15182;
      2754:data<=16'd14548;
      2755:data<=16'd14584;
      2756:data<=16'd14568;
      2757:data<=16'd15456;
      2758:data<=16'd15035;
      2759:data<=16'd11664;
      2760:data<=16'd7987;
      2761:data<=16'd6119;
      2762:data<=16'd5973;
      2763:data<=16'd5702;
      2764:data<=16'd5392;
      2765:data<=16'd5489;
      2766:data<=16'd4816;
      2767:data<=16'd4742;
      2768:data<=16'd4907;
      2769:data<=16'd4585;
      2770:data<=16'd5051;
      2771:data<=16'd4073;
      2772:data<=16'd3662;
      2773:data<=16'd5523;
      2774:data<=16'd4519;
      2775:data<=16'd3591;
      2776:data<=16'd4258;
      2777:data<=16'd2778;
      2778:data<=16'd3344;
      2779:data<=16'd3227;
      2780:data<=16'd1703;
      2781:data<=16'd5083;
      2782:data<=16'd36;
      2783:data<=-16'd14433;
      2784:data<=-16'd16915;
      2785:data<=-16'd13082;
      2786:data<=-16'd14314;
      2787:data<=-16'd13843;
      2788:data<=-16'd13106;
      2789:data<=-16'd12555;
      2790:data<=-16'd9629;
      2791:data<=-16'd9477;
      2792:data<=-16'd9944;
      2793:data<=-16'd8640;
      2794:data<=-16'd8951;
      2795:data<=-16'd9100;
      2796:data<=-16'd9022;
      2797:data<=-16'd9289;
      2798:data<=-16'd8029;
      2799:data<=-16'd7403;
      2800:data<=-16'd7544;
      2801:data<=-16'd7016;
      2802:data<=-16'd6852;
      2803:data<=-16'd6253;
      2804:data<=-16'd5943;
      2805:data<=-16'd6575;
      2806:data<=-16'd5283;
      2807:data<=-16'd3310;
      2808:data<=-16'd3416;
      2809:data<=-16'd2052;
      2810:data<=16'd2200;
      2811:data<=16'd3365;
      2812:data<=16'd1738;
      2813:data<=16'd2902;
      2814:data<=16'd3034;
      2815:data<=16'd1172;
      2816:data<=16'd2722;
      2817:data<=16'd3219;
      2818:data<=16'd2023;
      2819:data<=16'd3403;
      2820:data<=16'd2331;
      2821:data<=16'd1471;
      2822:data<=16'd3266;
      2823:data<=16'd1780;
      2824:data<=16'd7291;
      2825:data<=16'd20638;
      2826:data<=16'd22704;
      2827:data<=16'd18824;
      2828:data<=16'd20189;
      2829:data<=16'd19358;
      2830:data<=16'd17520;
      2831:data<=16'd17609;
      2832:data<=16'd15923;
      2833:data<=16'd15611;
      2834:data<=16'd16060;
      2835:data<=16'd14208;
      2836:data<=16'd13662;
      2837:data<=16'd14049;
      2838:data<=16'd12857;
      2839:data<=16'd12046;
      2840:data<=16'd12795;
      2841:data<=16'd13374;
      2842:data<=16'd12545;
      2843:data<=16'd11938;
      2844:data<=16'd11668;
      2845:data<=16'd10411;
      2846:data<=16'd9917;
      2847:data<=16'd9919;
      2848:data<=16'd8795;
      2849:data<=16'd7785;
      2850:data<=16'd7379;
      2851:data<=16'd7750;
      2852:data<=16'd7902;
      2853:data<=16'd6830;
      2854:data<=16'd6398;
      2855:data<=16'd5664;
      2856:data<=16'd5092;
      2857:data<=16'd6948;
      2858:data<=16'd6801;
      2859:data<=16'd3516;
      2860:data<=16'd123;
      2861:data<=-16'd2384;
      2862:data<=-16'd1181;
      2863:data<=-16'd597;
      2864:data<=-16'd2576;
      2865:data<=-16'd472;
      2866:data<=-16'd4211;
      2867:data<=-16'd17297;
      2868:data<=-16'd20861;
      2869:data<=-16'd17227;
      2870:data<=-16'd17935;
      2871:data<=-16'd17302;
      2872:data<=-16'd16131;
      2873:data<=-16'd16101;
      2874:data<=-16'd13602;
      2875:data<=-16'd12841;
      2876:data<=-16'd13065;
      2877:data<=-16'd11573;
      2878:data<=-16'd12029;
      2879:data<=-16'd12721;
      2880:data<=-16'd12028;
      2881:data<=-16'd11582;
      2882:data<=-16'd10813;
      2883:data<=-16'd10756;
      2884:data<=-16'd11009;
      2885:data<=-16'd10440;
      2886:data<=-16'd10173;
      2887:data<=-16'd9761;
      2888:data<=-16'd9364;
      2889:data<=-16'd8525;
      2890:data<=-16'd6526;
      2891:data<=-16'd5671;
      2892:data<=-16'd5538;
      2893:data<=-16'd5303;
      2894:data<=-16'd5782;
      2895:data<=-16'd5603;
      2896:data<=-16'd5341;
      2897:data<=-16'd5195;
      2898:data<=-16'd4604;
      2899:data<=-16'd4566;
      2900:data<=-16'd3266;
      2901:data<=-16'd2763;
      2902:data<=-16'd4341;
      2903:data<=-16'd2934;
      2904:data<=-16'd2299;
      2905:data<=-16'd3406;
      2906:data<=-16'd1313;
      2907:data<=-16'd1685;
      2908:data<=16'd1967;
      2909:data<=16'd17053;
      2910:data<=16'd24808;
      2911:data<=16'd22013;
      2912:data<=16'd21914;
      2913:data<=16'd20621;
      2914:data<=16'd18724;
      2915:data<=16'd19638;
      2916:data<=16'd17764;
      2917:data<=16'd16281;
      2918:data<=16'd16366;
      2919:data<=16'd14751;
      2920:data<=16'd15151;
      2921:data<=16'd15409;
      2922:data<=16'd13509;
      2923:data<=16'd13823;
      2924:data<=16'd14737;
      2925:data<=16'd14396;
      2926:data<=16'd13653;
      2927:data<=16'd12533;
      2928:data<=16'd12422;
      2929:data<=16'd12155;
      2930:data<=16'd11010;
      2931:data<=16'd10269;
      2932:data<=16'd9147;
      2933:data<=16'd8830;
      2934:data<=16'd9015;
      2935:data<=16'd7586;
      2936:data<=16'd7201;
      2937:data<=16'd8084;
      2938:data<=16'd7212;
      2939:data<=16'd5883;
      2940:data<=16'd6379;
      2941:data<=16'd7351;
      2942:data<=16'd6384;
      2943:data<=16'd5298;
      2944:data<=16'd5429;
      2945:data<=16'd4610;
      2946:data<=16'd4287;
      2947:data<=16'd3809;
      2948:data<=16'd2719;
      2949:data<=16'd4461;
      2950:data<=-16'd217;
      2951:data<=-16'd13180;
      2952:data<=-16'd16725;
      2953:data<=-16'd13761;
      2954:data<=-16'd15106;
      2955:data<=-16'd14343;
      2956:data<=-16'd14043;
      2957:data<=-16'd15702;
      2958:data<=-16'd13076;
      2959:data<=-16'd14095;
      2960:data<=-16'd18968;
      2961:data<=-16'd18592;
      2962:data<=-16'd17814;
      2963:data<=-16'd18624;
      2964:data<=-16'd18036;
      2965:data<=-16'd18089;
      2966:data<=-16'd17303;
      2967:data<=-16'd16013;
      2968:data<=-16'd16263;
      2969:data<=-16'd15769;
      2970:data<=-16'd15244;
      2971:data<=-16'd15306;
      2972:data<=-16'd14389;
      2973:data<=-16'd14170;
      2974:data<=-16'd14980;
      2975:data<=-16'd14968;
      2976:data<=-16'd14222;
      2977:data<=-16'd13705;
      2978:data<=-16'd13778;
      2979:data<=-16'd14076;
      2980:data<=-16'd13837;
      2981:data<=-16'd12543;
      2982:data<=-16'd11661;
      2983:data<=-16'd11706;
      2984:data<=-16'd10640;
      2985:data<=-16'd9868;
      2986:data<=-16'd10052;
      2987:data<=-16'd9635;
      2988:data<=-16'd10499;
      2989:data<=-16'd10245;
      2990:data<=-16'd9342;
      2991:data<=-16'd12278;
      2992:data<=-16'd7553;
      2993:data<=16'd6035;
      2994:data<=16'd9307;
      2995:data<=16'd6417;
      2996:data<=16'd8291;
      2997:data<=16'd7465;
      2998:data<=16'd5632;
      2999:data<=16'd6526;
      3000:data<=16'd5971;
      3001:data<=16'd6219;
      3002:data<=16'd6440;
      3003:data<=16'd4927;
      3004:data<=16'd5025;
      3005:data<=16'd5131;
      3006:data<=16'd4980;
      3007:data<=16'd4611;
      3008:data<=16'd2364;
      3009:data<=16'd3401;
      3010:data<=16'd7421;
      3011:data<=16'd8322;
      3012:data<=16'd7752;
      3013:data<=16'd7532;
      3014:data<=16'd7269;
      3015:data<=16'd7315;
      3016:data<=16'd6763;
      3017:data<=16'd6520;
      3018:data<=16'd6485;
      3019:data<=16'd5658;
      3020:data<=16'd5430;
      3021:data<=16'd5589;
      3022:data<=16'd5275;
      3023:data<=16'd3967;
      3024:data<=16'd2303;
      3025:data<=16'd2111;
      3026:data<=16'd1477;
      3027:data<=16'd638;
      3028:data<=16'd1277;
      3029:data<=16'd996;
      3030:data<=16'd1199;
      3031:data<=16'd1063;
      3032:data<=-16'd567;
      3033:data<=16'd1516;
      3034:data<=-16'd1389;
      3035:data<=-16'd13946;
      3036:data<=-16'd18666;
      3037:data<=-16'd15911;
      3038:data<=-16'd16448;
      3039:data<=-16'd15338;
      3040:data<=-16'd14901;
      3041:data<=-16'd17138;
      3042:data<=-16'd15978;
      3043:data<=-16'd15291;
      3044:data<=-16'd15476;
      3045:data<=-16'd13775;
      3046:data<=-16'd14428;
      3047:data<=-16'd15132;
      3048:data<=-16'd13603;
      3049:data<=-16'd12728;
      3050:data<=-16'd11917;
      3051:data<=-16'd11670;
      3052:data<=-16'd11770;
      3053:data<=-16'd11207;
      3054:data<=-16'd11151;
      3055:data<=-16'd10419;
      3056:data<=-16'd10434;
      3057:data<=-16'd12037;
      3058:data<=-16'd11395;
      3059:data<=-16'd10828;
      3060:data<=-16'd13085;
      3061:data<=-16'd14650;
      3062:data<=-16'd14186;
      3063:data<=-16'd13402;
      3064:data<=-16'd13529;
      3065:data<=-16'd12930;
      3066:data<=-16'd11116;
      3067:data<=-16'd10551;
      3068:data<=-16'd9558;
      3069:data<=-16'd8555;
      3070:data<=-16'd9544;
      3071:data<=-16'd8868;
      3072:data<=-16'd7890;
      3073:data<=-16'd8200;
      3074:data<=-16'd8219;
      3075:data<=-16'd10480;
      3076:data<=-16'd7269;
      3077:data<=16'd4529;
      3078:data<=16'd8962;
      3079:data<=16'd6469;
      3080:data<=16'd7397;
      3081:data<=16'd7542;
      3082:data<=16'd7097;
      3083:data<=16'd7782;
      3084:data<=16'd6511;
      3085:data<=16'd6199;
      3086:data<=16'd6416;
      3087:data<=16'd5319;
      3088:data<=16'd5664;
      3089:data<=16'd5915;
      3090:data<=16'd4708;
      3091:data<=16'd3419;
      3092:data<=16'd2904;
      3093:data<=16'd3659;
      3094:data<=16'd3415;
      3095:data<=16'd2789;
      3096:data<=16'd3667;
      3097:data<=16'd3388;
      3098:data<=16'd2870;
      3099:data<=16'd3688;
      3100:data<=16'd3776;
      3101:data<=16'd3785;
      3102:data<=16'd3694;
      3103:data<=16'd2828;
      3104:data<=16'd2587;
      3105:data<=16'd3054;
      3106:data<=16'd3768;
      3107:data<=16'd2922;
      3108:data<=16'd537;
      3109:data<=16'd652;
      3110:data<=16'd3479;
      3111:data<=16'd6472;
      3112:data<=16'd7453;
      3113:data<=16'd6319;
      3114:data<=16'd6821;
      3115:data<=16'd7103;
      3116:data<=16'd5885;
      3117:data<=16'd7370;
      3118:data<=16'd4294;
      3119:data<=-16'd6276;
      3120:data<=-16'd10916;
      3121:data<=-16'd9147;
      3122:data<=-16'd9200;
      3123:data<=-16'd9687;
      3124:data<=-16'd10366;
      3125:data<=-16'd10721;
      3126:data<=-16'd8981;
      3127:data<=-16'd8551;
      3128:data<=-16'd8980;
      3129:data<=-16'd7682;
      3130:data<=-16'd6912;
      3131:data<=-16'd7392;
      3132:data<=-16'd7661;
      3133:data<=-16'd7142;
      3134:data<=-16'd6299;
      3135:data<=-16'd5965;
      3136:data<=-16'd5515;
      3137:data<=-16'd5281;
      3138:data<=-16'd5471;
      3139:data<=-16'd4672;
      3140:data<=-16'd4821;
      3141:data<=-16'd6528;
      3142:data<=-16'd6334;
      3143:data<=-16'd5318;
      3144:data<=-16'd5598;
      3145:data<=-16'd5486;
      3146:data<=-16'd5057;
      3147:data<=-16'd4805;
      3148:data<=-16'd4255;
      3149:data<=-16'd4134;
      3150:data<=-16'd4009;
      3151:data<=-16'd3416;
      3152:data<=-16'd2814;
      3153:data<=-16'd2096;
      3154:data<=-16'd1991;
      3155:data<=-16'd2229;
      3156:data<=-16'd2243;
      3157:data<=-16'd3043;
      3158:data<=-16'd3630;
      3159:data<=-16'd3745;
      3160:data<=-16'd2946;
      3161:data<=16'd1997;
      3162:data<=16'd6802;
      3163:data<=16'd6434;
      3164:data<=16'd5935;
      3165:data<=16'd6273;
      3166:data<=16'd5383;
      3167:data<=16'd6011;
      3168:data<=16'd6422;
      3169:data<=16'd5620;
      3170:data<=16'd5729;
      3171:data<=16'd4802;
      3172:data<=16'd4455;
      3173:data<=16'd5833;
      3174:data<=16'd4666;
      3175:data<=16'd2532;
      3176:data<=16'd2520;
      3177:data<=16'd3398;
      3178:data<=16'd4152;
      3179:data<=16'd3588;
      3180:data<=16'd2889;
      3181:data<=16'd3275;
      3182:data<=16'd3369;
      3183:data<=16'd4091;
      3184:data<=16'd4499;
      3185:data<=16'd3310;
      3186:data<=16'd3166;
      3187:data<=16'd3140;
      3188:data<=16'd2590;
      3189:data<=16'd3468;
      3190:data<=16'd3383;
      3191:data<=16'd1735;
      3192:data<=16'd784;
      3193:data<=16'd303;
      3194:data<=16'd438;
      3195:data<=16'd966;
      3196:data<=16'd1119;
      3197:data<=16'd1342;
      3198:data<=16'd1478;
      3199:data<=16'd1008;
      3200:data<=16'd664;
      3201:data<=16'd2073;
      3202:data<=16'd699;
      3203:data<=-16'd8455;
      3204:data<=-16'd15209;
      3205:data<=-16'd13459;
      3206:data<=-16'd12540;
      3207:data<=-16'd12636;
      3208:data<=-16'd11723;
      3209:data<=-16'd13429;
      3210:data<=-16'd11226;
      3211:data<=-16'd5043;
      3212:data<=-16'd3994;
      3213:data<=-16'd4485;
      3214:data<=-16'd3350;
      3215:data<=-16'd3782;
      3216:data<=-16'd3756;
      3217:data<=-16'd3057;
      3218:data<=-16'd3113;
      3219:data<=-16'd2813;
      3220:data<=-16'd2517;
      3221:data<=-16'd2046;
      3222:data<=-16'd1504;
      3223:data<=-16'd1850;
      3224:data<=-16'd2059;
      3225:data<=-16'd1792;
      3226:data<=-16'd1415;
      3227:data<=-16'd995;
      3228:data<=-16'd813;
      3229:data<=-16'd453;
      3230:data<=-16'd133;
      3231:data<=-16'd9;
      3232:data<=16'd161;
      3233:data<=-16'd103;
      3234:data<=16'd112;
      3235:data<=16'd1202;
      3236:data<=16'd1865;
      3237:data<=16'd2046;
      3238:data<=16'd1996;
      3239:data<=16'd1902;
      3240:data<=16'd2214;
      3241:data<=16'd3338;
      3242:data<=16'd4334;
      3243:data<=16'd2936;
      3244:data<=16'd4309;
      3245:data<=16'd13461;
      3246:data<=16'd19831;
      3247:data<=16'd18160;
      3248:data<=16'd17578;
      3249:data<=16'd18048;
      3250:data<=16'd16430;
      3251:data<=16'd16207;
      3252:data<=16'd15943;
      3253:data<=16'd14971;
      3254:data<=16'd15371;
      3255:data<=16'd15039;
      3256:data<=16'd14263;
      3257:data<=16'd14337;
      3258:data<=16'd14604;
      3259:data<=16'd15282;
      3260:data<=16'd13264;
      3261:data<=16'd8522;
      3262:data<=16'd7098;
      3263:data<=16'd7847;
      3264:data<=16'd6760;
      3265:data<=16'd6093;
      3266:data<=16'd6487;
      3267:data<=16'd6176;
      3268:data<=16'd5926;
      3269:data<=16'd6050;
      3270:data<=16'd5937;
      3271:data<=16'd5815;
      3272:data<=16'd5203;
      3273:data<=16'd4634;
      3274:data<=16'd6138;
      3275:data<=16'd7583;
      3276:data<=16'd6510;
      3277:data<=16'd6105;
      3278:data<=16'd6675;
      3279:data<=16'd5911;
      3280:data<=16'd5841;
      3281:data<=16'd6185;
      3282:data<=16'd5416;
      3283:data<=16'd4567;
      3284:data<=16'd3485;
      3285:data<=16'd4008;
      3286:data<=16'd3463;
      3287:data<=-16'd4284;
      3288:data<=-16'd11298;
      3289:data<=-16'd11311;
      3290:data<=-16'd11006;
      3291:data<=-16'd9876;
      3292:data<=-16'd7212;
      3293:data<=-16'd7473;
      3294:data<=-16'd7341;
      3295:data<=-16'd6040;
      3296:data<=-16'd6164;
      3297:data<=-16'd5451;
      3298:data<=-16'd4796;
      3299:data<=-16'd5148;
      3300:data<=-16'd5259;
      3301:data<=-16'd5406;
      3302:data<=-16'd4537;
      3303:data<=-16'd4043;
      3304:data<=-16'd4490;
      3305:data<=-16'd3932;
      3306:data<=-16'd4285;
      3307:data<=-16'd3530;
      3308:data<=-16'd970;
      3309:data<=-16'd1624;
      3310:data<=-16'd353;
      3311:data<=16'd5225;
      3312:data<=16'd6780;
      3313:data<=16'd5604;
      3314:data<=16'd5824;
      3315:data<=16'd5912;
      3316:data<=16'd5879;
      3317:data<=16'd5154;
      3318:data<=16'd4857;
      3319:data<=16'd5541;
      3320:data<=16'd5106;
      3321:data<=16'd5365;
      3322:data<=16'd5529;
      3323:data<=16'd4167;
      3324:data<=16'd4913;
      3325:data<=16'd6622;
      3326:data<=16'd6966;
      3327:data<=16'd6305;
      3328:data<=16'd6329;
      3329:data<=16'd12818;
      3330:data<=16'd21079;
      3331:data<=16'd21329;
      3332:data<=16'd19276;
      3333:data<=16'd19079;
      3334:data<=16'd17450;
      3335:data<=16'd16954;
      3336:data<=16'd17208;
      3337:data<=16'd15946;
      3338:data<=16'd15206;
      3339:data<=16'd14595;
      3340:data<=16'd14249;
      3341:data<=16'd15385;
      3342:data<=16'd16187;
      3343:data<=16'd15544;
      3344:data<=16'd14563;
      3345:data<=16'd14501;
      3346:data<=16'd14048;
      3347:data<=16'd12568;
      3348:data<=16'd12287;
      3349:data<=16'd11752;
      3350:data<=16'd10387;
      3351:data<=16'd10566;
      3352:data<=16'd10011;
      3353:data<=16'd8696;
      3354:data<=16'd8663;
      3355:data<=16'd8025;
      3356:data<=16'd7626;
      3357:data<=16'd7727;
      3358:data<=16'd8094;
      3359:data<=16'd10196;
      3360:data<=16'd8325;
      3361:data<=16'd2366;
      3362:data<=16'd720;
      3363:data<=16'd966;
      3364:data<=16'd290;
      3365:data<=16'd848;
      3366:data<=-16'd203;
      3367:data<=-16'd1465;
      3368:data<=-16'd1028;
      3369:data<=-16'd676;
      3370:data<=-16'd249;
      3371:data<=-16'd5900;
      3372:data<=-16'd16219;
      3373:data<=-16'd17628;
      3374:data<=-16'd13712;
      3375:data<=-16'd13230;
      3376:data<=-16'd12305;
      3377:data<=-16'd11800;
      3378:data<=-16'd12214;
      3379:data<=-16'd10505;
      3380:data<=-16'd10386;
      3381:data<=-16'd11257;
      3382:data<=-16'd10345;
      3383:data<=-16'd10536;
      3384:data<=-16'd10701;
      3385:data<=-16'd9633;
      3386:data<=-16'd9812;
      3387:data<=-16'd10108;
      3388:data<=-16'd9250;
      3389:data<=-16'd8727;
      3390:data<=-16'd8880;
      3391:data<=-16'd8056;
      3392:data<=-16'd6152;
      3393:data<=-16'd5723;
      3394:data<=-16'd6202;
      3395:data<=-16'd5595;
      3396:data<=-16'd5322;
      3397:data<=-16'd5648;
      3398:data<=-16'd5533;
      3399:data<=-16'd5057;
      3400:data<=-16'd4790;
      3401:data<=-16'd5143;
      3402:data<=-16'd4538;
      3403:data<=-16'd3747;
      3404:data<=-16'd4385;
      3405:data<=-16'd4135;
      3406:data<=-16'd4193;
      3407:data<=-16'd4419;
      3408:data<=-16'd1994;
      3409:data<=-16'd1227;
      3410:data<=-16'd343;
      3411:data<=16'd3660;
      3412:data<=16'd4651;
      3413:data<=16'd9236;
      3414:data<=16'd19705;
      3415:data<=16'd21203;
      3416:data<=16'd18102;
      3417:data<=16'd19186;
      3418:data<=16'd17672;
      3419:data<=16'd15904;
      3420:data<=16'd16063;
      3421:data<=16'd14377;
      3422:data<=16'd14257;
      3423:data<=16'd14430;
      3424:data<=16'd13294;
      3425:data<=16'd14348;
      3426:data<=16'd15051;
      3427:data<=16'd14142;
      3428:data<=16'd13098;
      3429:data<=16'd11819;
      3430:data<=16'd11491;
      3431:data<=16'd10963;
      3432:data<=16'd10276;
      3433:data<=16'd10147;
      3434:data<=16'd8749;
      3435:data<=16'd8269;
      3436:data<=16'd8573;
      3437:data<=16'd7530;
      3438:data<=16'd7418;
      3439:data<=16'd6620;
      3440:data<=16'd5313;
      3441:data<=16'd6774;
      3442:data<=16'd7868;
      3443:data<=16'd7567;
      3444:data<=16'd6843;
      3445:data<=16'd5521;
      3446:data<=16'd5498;
      3447:data<=16'd4990;
      3448:data<=16'd3987;
      3449:data<=16'd3903;
      3450:data<=16'd2446;
      3451:data<=16'd2262;
      3452:data<=16'd2312;
      3453:data<=16'd937;
      3454:data<=16'd3008;
      3455:data<=-16'd654;
      3456:data<=-16'd12463;
      3457:data<=-16'd15341;
      3458:data<=-16'd12166;
      3459:data<=-16'd12155;
      3460:data<=-16'd11749;
      3461:data<=-16'd14533;
      3462:data<=-16'd18107;
      3463:data<=-16'd16521;
      3464:data<=-16'd16257;
      3465:data<=-16'd17176;
      3466:data<=-16'd16183;
      3467:data<=-16'd16178;
      3468:data<=-16'd15749;
      3469:data<=-16'd15057;
      3470:data<=-16'd15015;
      3471:data<=-16'd14038;
      3472:data<=-16'd13747;
      3473:data<=-16'd13759;
      3474:data<=-16'd12897;
      3475:data<=-16'd11829;
      3476:data<=-16'd10508;
      3477:data<=-16'd10376;
      3478:data<=-16'd10255;
      3479:data<=-16'd9054;
      3480:data<=-16'd9050;
      3481:data<=-16'd8790;
      3482:data<=-16'd8328;
      3483:data<=-16'd8925;
      3484:data<=-16'd8117;
      3485:data<=-16'd7597;
      3486:data<=-16'd8375;
      3487:data<=-16'd8028;
      3488:data<=-16'd7451;
      3489:data<=-16'd6843;
      3490:data<=-16'd6680;
      3491:data<=-16'd6843;
      3492:data<=-16'd5927;
      3493:data<=-16'd6431;
      3494:data<=-16'd6310;
      3495:data<=-16'd5175;
      3496:data<=-16'd7412;
      3497:data<=-16'd3325;
      3498:data<=16'd8408;
      3499:data<=16'd11268;
      3500:data<=16'd8298;
      3501:data<=16'd8701;
      3502:data<=16'd7937;
      3503:data<=16'd7336;
      3504:data<=16'd7532;
      3505:data<=16'd5730;
      3506:data<=16'd5586;
      3507:data<=16'd6200;
      3508:data<=16'd5427;
      3509:data<=16'd4610;
      3510:data<=16'd3498;
      3511:data<=16'd5303;
      3512:data<=16'd9103;
      3513:data<=16'd9309;
      3514:data<=16'd8331;
      3515:data<=16'd8088;
      3516:data<=16'd7470;
      3517:data<=16'd7735;
      3518:data<=16'd7279;
      3519:data<=16'd6249;
      3520:data<=16'd6375;
      3521:data<=16'd5577;
      3522:data<=16'd4792;
      3523:data<=16'd5271;
      3524:data<=16'd4786;
      3525:data<=16'd3475;
      3526:data<=16'd2208;
      3527:data<=16'd1321;
      3528:data<=16'd1060;
      3529:data<=16'd425;
      3530:data<=-16'd170;
      3531:data<=-16'd109;
      3532:data<=-16'd112;
      3533:data<=-16'd649;
      3534:data<=-16'd1104;
      3535:data<=-16'd710;
      3536:data<=-16'd1433;
      3537:data<=-16'd1691;
      3538:data<=16'd619;
      3539:data<=-16'd3889;
      3540:data<=-16'd14778;
      3541:data<=-16'd17693;
      3542:data<=-16'd16167;
      3543:data<=-16'd17787;
      3544:data<=-16'd17327;
      3545:data<=-16'd16399;
      3546:data<=-16'd16688;
      3547:data<=-16'd15136;
      3548:data<=-16'd14844;
      3549:data<=-16'd15591;
      3550:data<=-16'd14962;
      3551:data<=-16'd14073;
      3552:data<=-16'd13022;
      3553:data<=-16'd13091;
      3554:data<=-16'd13142;
      3555:data<=-16'd12154;
      3556:data<=-16'd12281;
      3557:data<=-16'd11409;
      3558:data<=-16'd11317;
      3559:data<=-16'd13480;
      3560:data<=-16'd12627;
      3561:data<=-16'd13652;
      3562:data<=-16'd18384;
      3563:data<=-16'd18289;
      3564:data<=-16'd16826;
      3565:data<=-16'd17150;
      3566:data<=-16'd16060;
      3567:data<=-16'd16014;
      3568:data<=-16'd15591;
      3569:data<=-16'd14148;
      3570:data<=-16'd14002;
      3571:data<=-16'd12533;
      3572:data<=-16'd11641;
      3573:data<=-16'd12231;
      3574:data<=-16'd11245;
      3575:data<=-16'd11113;
      3576:data<=-16'd11919;
      3577:data<=-16'd12034;
      3578:data<=-16'd11112;
      3579:data<=-16'd9803;
      3580:data<=-16'd11110;
      3581:data<=-16'd7189;
      3582:data<=16'd4056;
      3583:data<=16'd7262;
      3584:data<=16'd5074;
      3585:data<=16'd6730;
      3586:data<=16'd6047;
      3587:data<=16'd5131;
      3588:data<=16'd6287;
      3589:data<=16'd5280;
      3590:data<=16'd5356;
      3591:data<=16'd5492;
      3592:data<=16'd3744;
      3593:data<=16'd3106;
      3594:data<=16'd2408;
      3595:data<=16'd2458;
      3596:data<=16'd3196;
      3597:data<=16'd2517;
      3598:data<=16'd2435;
      3599:data<=16'd2347;
      3600:data<=16'd2532;
      3601:data<=16'd3397;
      3602:data<=16'd2516;
      3603:data<=16'd2641;
      3604:data<=16'd3236;
      3605:data<=16'd2576;
      3606:data<=16'd3424;
      3607:data<=16'd2728;
      3608:data<=16'd1448;
      3609:data<=16'd1750;
      3610:data<=-16'd82;
      3611:data<=16'd1494;
      3612:data<=16'd6246;
      3613:data<=16'd6543;
      3614:data<=16'd6711;
      3615:data<=16'd6905;
      3616:data<=16'd5656;
      3617:data<=16'd6661;
      3618:data<=16'd6291;
      3619:data<=16'd5444;
      3620:data<=16'd5342;
      3621:data<=16'd4068;
      3622:data<=16'd6008;
      3623:data<=16'd3130;
      3624:data<=-16'd7809;
      3625:data<=-16'd11828;
      3626:data<=-16'd11435;
      3627:data<=-16'd12677;
      3628:data<=-16'd11129;
      3629:data<=-16'd11151;
      3630:data<=-16'd11497;
      3631:data<=-16'd9411;
      3632:data<=-16'd9691;
      3633:data<=-16'd9379;
      3634:data<=-16'd8311;
      3635:data<=-16'd8633;
      3636:data<=-16'd7565;
      3637:data<=-16'd7353;
      3638:data<=-16'd7213;
      3639:data<=-16'd6097;
      3640:data<=-16'd6578;
      3641:data<=-16'd5788;
      3642:data<=-16'd5664;
      3643:data<=-16'd7538;
      3644:data<=-16'd6896;
      3645:data<=-16'd6492;
      3646:data<=-16'd6572;
      3647:data<=-16'd5523;
      3648:data<=-16'd5557;
      3649:data<=-16'd4231;
      3650:data<=-16'd3457;
      3651:data<=-16'd4466;
      3652:data<=-16'd3441;
      3653:data<=-16'd3495;
      3654:data<=-16'd3412;
      3655:data<=-16'd2112;
      3656:data<=-16'd3403;
      3657:data<=-16'd2356;
      3658:data<=-16'd1633;
      3659:data<=-16'd4499;
      3660:data<=-16'd3421;
      3661:data<=-16'd4444;
      3662:data<=-16'd8752;
      3663:data<=-16'd8275;
      3664:data<=-16'd9317;
      3665:data<=-16'd6385;
      3666:data<=16'd5527;
      3667:data<=16'd9244;
      3668:data<=16'd6255;
      3669:data<=16'd7265;
      3670:data<=16'd7210;
      3671:data<=16'd6998;
      3672:data<=16'd7721;
      3673:data<=16'd6470;
      3674:data<=16'd6393;
      3675:data<=16'd6326;
      3676:data<=16'd4733;
      3677:data<=16'd3964;
      3678:data<=16'd3802;
      3679:data<=16'd4493;
      3680:data<=16'd4761;
      3681:data<=16'd4141;
      3682:data<=16'd4758;
      3683:data<=16'd4752;
      3684:data<=16'd4097;
      3685:data<=16'd4613;
      3686:data<=16'd4614;
      3687:data<=16'd4385;
      3688:data<=16'd4487;
      3689:data<=16'd4346;
      3690:data<=16'd4546;
      3691:data<=16'd4369;
      3692:data<=16'd3341;
      3693:data<=16'd1750;
      3694:data<=16'd1184;
      3695:data<=16'd2382;
      3696:data<=16'd1996;
      3697:data<=16'd1339;
      3698:data<=16'd2241;
      3699:data<=16'd1233;
      3700:data<=16'd1119;
      3701:data<=16'd2331;
      3702:data<=16'd1168;
      3703:data<=16'd1861;
      3704:data<=16'd2259;
      3705:data<=16'd681;
      3706:data<=16'd3096;
      3707:data<=16'd79;
      3708:data<=-16'd11088;
      3709:data<=-16'd15289;
      3710:data<=-16'd14540;
      3711:data<=-16'd13640;
      3712:data<=-16'd8407;
      3713:data<=-16'd5419;
      3714:data<=-16'd5865;
      3715:data<=-16'd4343;
      3716:data<=-16'd4102;
      3717:data<=-16'd4678;
      3718:data<=-16'd4225;
      3719:data<=-16'd4137;
      3720:data<=-16'd2980;
      3721:data<=-16'd2607;
      3722:data<=-16'd3542;
      3723:data<=-16'd2795;
      3724:data<=-16'd2261;
      3725:data<=-16'd2901;
      3726:data<=-16'd3477;
      3727:data<=-16'd4038;
      3728:data<=-16'd3911;
      3729:data<=-16'd3644;
      3730:data<=-16'd3210;
      3731:data<=-16'd2535;
      3732:data<=-16'd2599;
      3733:data<=-16'd1926;
      3734:data<=-16'd1231;
      3735:data<=-16'd1765;
      3736:data<=-16'd1606;
      3737:data<=-16'd1037;
      3738:data<=-16'd232;
      3739:data<=16'd224;
      3740:data<=-16'd337;
      3741:data<=16'd520;
      3742:data<=16'd197;
      3743:data<=-16'd1569;
      3744:data<=-16'd412;
      3745:data<=-16'd394;
      3746:data<=-16'd576;
      3747:data<=16'd1486;
      3748:data<=-16'd214;
      3749:data<=16'd2560;
      3750:data<=16'd13526;
      3751:data<=16'd16913;
      3752:data<=16'd14469;
      3753:data<=16'd15192;
      3754:data<=16'd14906;
      3755:data<=16'd14357;
      3756:data<=16'd14327;
      3757:data<=16'd13082;
      3758:data<=16'd12924;
      3759:data<=16'd12903;
      3760:data<=16'd12924;
      3761:data<=16'd11790;
      3762:data<=16'd7268;
      3763:data<=16'd4845;
      3764:data<=16'd5148;
      3765:data<=16'd4661;
      3766:data<=16'd5233;
      3767:data<=16'd5266;
      3768:data<=16'd4538;
      3769:data<=16'd5274;
      3770:data<=16'd5045;
      3771:data<=16'd4620;
      3772:data<=16'd5406;
      3773:data<=16'd5547;
      3774:data<=16'd5153;
      3775:data<=16'd4799;
      3776:data<=16'd5559;
      3777:data<=16'd6619;
      3778:data<=16'd6611;
      3779:data<=16'd7181;
      3780:data<=16'd6633;
      3781:data<=16'd5624;
      3782:data<=16'd6677;
      3783:data<=16'd5838;
      3784:data<=16'd4942;
      3785:data<=16'd6100;
      3786:data<=16'd5230;
      3787:data<=16'd5365;
      3788:data<=16'd5465;
      3789:data<=16'd3554;
      3790:data<=16'd5532;
      3791:data<=16'd3174;
      3792:data<=-16'd7154;
      3793:data<=-16'd10155;
      3794:data<=-16'd7263;
      3795:data<=-16'd7492;
      3796:data<=-16'd7028;
      3797:data<=-16'd6040;
      3798:data<=-16'd6261;
      3799:data<=-16'd5985;
      3800:data<=-16'd5747;
      3801:data<=-16'd5459;
      3802:data<=-16'd5379;
      3803:data<=-16'd4861;
      3804:data<=-16'd3738;
      3805:data<=-16'd4140;
      3806:data<=-16'd3988;
      3807:data<=-16'd3016;
      3808:data<=-16'd3610;
      3809:data<=-16'd2934;
      3810:data<=-16'd987;
      3811:data<=16'd365;
      3812:data<=16'd3207;
      3813:data<=16'd6305;
      3814:data<=16'd7083;
      3815:data<=16'd6276;
      3816:data<=16'd5858;
      3817:data<=16'd6467;
      3818:data<=16'd5994;
      3819:data<=16'd5184;
      3820:data<=16'd5808;
      3821:data<=16'd5747;
      3822:data<=16'd5251;
      3823:data<=16'd5080;
      3824:data<=16'd4670;
      3825:data<=16'd5510;
      3826:data<=16'd6575;
      3827:data<=16'd7341;
      3828:data<=16'd8147;
      3829:data<=16'd7003;
      3830:data<=16'd7292;
      3831:data<=16'd8827;
      3832:data<=16'd6378;
      3833:data<=16'd8155;
      3834:data<=16'd17779;
      3835:data<=16'd22306;
      3836:data<=16'd20465;
      3837:data<=16'd20005;
      3838:data<=16'd19600;
      3839:data<=16'd18289;
      3840:data<=16'd17676;
      3841:data<=16'd16918;
      3842:data<=16'd16463;
      3843:data<=16'd16932;
      3844:data<=16'd17317;
      3845:data<=16'd17006;
      3846:data<=16'd16180;
      3847:data<=16'd15320;
      3848:data<=16'd14737;
      3849:data<=16'd14721;
      3850:data<=16'd14715;
      3851:data<=16'd13608;
      3852:data<=16'd12466;
      3853:data<=16'd12496;
      3854:data<=16'd12366;
      3855:data<=16'd11341;
      3856:data<=16'd10417;
      3857:data<=16'd10038;
      3858:data<=16'd9730;
      3859:data<=16'd9652;
      3860:data<=16'd10461;
      3861:data<=16'd10275;
      3862:data<=16'd7037;
      3863:data<=16'd3582;
      3864:data<=16'd2591;
      3865:data<=16'd2581;
      3866:data<=16'd2311;
      3867:data<=16'd1592;
      3868:data<=16'd751;
      3869:data<=16'd522;
      3870:data<=16'd593;
      3871:data<=16'd914;
      3872:data<=16'd379;
      3873:data<=-16'd1037;
      3874:data<=-16'd167;
      3875:data<=-16'd1583;
      3876:data<=-16'd10072;
      3877:data<=-16'd15443;
      3878:data<=-16'd13502;
      3879:data<=-16'd12792;
      3880:data<=-16'd13032;
      3881:data<=-16'd11793;
      3882:data<=-16'd11843;
      3883:data<=-16'd11659;
      3884:data<=-16'd10796;
      3885:data<=-16'd11048;
      3886:data<=-16'd11273;
      3887:data<=-16'd10980;
      3888:data<=-16'd10019;
      3889:data<=-16'd9091;
      3890:data<=-16'd9659;
      3891:data<=-16'd10190;
      3892:data<=-16'd9468;
      3893:data<=-16'd7829;
      3894:data<=-16'd6299;
      3895:data<=-16'd6346;
      3896:data<=-16'd6170;
      3897:data<=-16'd5016;
      3898:data<=-16'd5080;
      3899:data<=-16'd5507;
      3900:data<=-16'd5112;
      3901:data<=-16'd4601;
      3902:data<=-16'd4464;
      3903:data<=-16'd4802;
      3904:data<=-16'd4984;
      3905:data<=-16'd5210;
      3906:data<=-16'd4868;
      3907:data<=-16'd4005;
      3908:data<=-16'd4834;
      3909:data<=-16'd4297;
      3910:data<=-16'd1841;
      3911:data<=-16'd1833;
      3912:data<=16'd331;
      3913:data<=16'd5066;
      3914:data<=16'd5894;
      3915:data<=16'd5679;
      3916:data<=16'd4943;
      3917:data<=16'd5436;
      3918:data<=16'd13919;
      3919:data<=16'd20539;
      3920:data<=16'd18665;
      3921:data<=16'd17535;
      3922:data<=16'd16607;
      3923:data<=16'd14662;
      3924:data<=16'd15127;
      3925:data<=16'd14440;
      3926:data<=16'd13978;
      3927:data<=16'd15562;
      3928:data<=16'd15341;
      3929:data<=16'd14706;
      3930:data<=16'd14052;
      3931:data<=16'd12518;
      3932:data<=16'd12173;
      3933:data<=16'd11705;
      3934:data<=16'd10903;
      3935:data<=16'd10469;
      3936:data<=16'd9494;
      3937:data<=16'd9580;
      3938:data<=16'd9338;
      3939:data<=16'd7467;
      3940:data<=16'd7144;
      3941:data<=16'd7492;
      3942:data<=16'd6912;
      3943:data<=16'd6993;
      3944:data<=16'd7750;
      3945:data<=16'd8132;
      3946:data<=16'd7286;
      3947:data<=16'd6458;
      3948:data<=16'd6448;
      3949:data<=16'd5521;
      3950:data<=16'd4933;
      3951:data<=16'd4734;
      3952:data<=16'd3119;
      3953:data<=16'd2356;
      3954:data<=16'd2511;
      3955:data<=16'd2247;
      3956:data<=16'd1686;
      3957:data<=16'd311;
      3958:data<=16'd984;
      3959:data<=16'd702;
      3960:data<=-16'd6448;
      3961:data<=-16'd12493;
      3962:data<=-16'd14198;
      3963:data<=-16'd17794;
      3964:data<=-16'd19105;
      3965:data<=-16'd17280;
      3966:data<=-16'd17640;
      3967:data<=-16'd17300;
      3968:data<=-16'd16137;
      3969:data<=-16'd16563;
      3970:data<=-16'd16536;
      3971:data<=-16'd16501;
      3972:data<=-16'd16126;
      3973:data<=-16'd14630;
      3974:data<=-16'd14440;
      3975:data<=-16'd14741;
      3976:data<=-16'd13769;
      3977:data<=-16'd12270;
      3978:data<=-16'd11030;
      3979:data<=-16'd10994;
      3980:data<=-16'd11133;
      3981:data<=-16'd10302;
      3982:data<=-16'd9928;
      3983:data<=-16'd10135;
      3984:data<=-16'd9982;
      3985:data<=-16'd9364;
      3986:data<=-16'd8802;
      3987:data<=-16'd8987;
      3988:data<=-16'd9250;
      3989:data<=-16'd9194;
      3990:data<=-16'd8848;
      3991:data<=-16'd8226;
      3992:data<=-16'd8193;
      3993:data<=-16'd7339;
      3994:data<=-16'd5454;
      3995:data<=-16'd5201;
      3996:data<=-16'd5137;
      3997:data<=-16'd4704;
      3998:data<=-16'd5113;
      3999:data<=-16'd4196;
      4000:data<=-16'd4147;
      4001:data<=-16'd4256;
      4002:data<=16'd3016;
      4003:data<=16'd11585;
      4004:data<=16'd11762;
      4005:data<=16'd9580;
      4006:data<=16'd9747;
      4007:data<=16'd8916;
      4008:data<=16'd7724;
      4009:data<=16'd8396;
      4010:data<=16'd8951;
      4011:data<=16'd8294;
      4012:data<=16'd10363;
      4013:data<=16'd14439;
      4014:data<=16'd14433;
      4015:data<=16'd12739;
      4016:data<=16'd12819;
      4017:data<=16'd12029;
      4018:data<=16'd11721;
      4019:data<=16'd11715;
      4020:data<=16'd10170;
      4021:data<=16'd10580;
      4022:data<=16'd10939;
      4023:data<=16'd8625;
      4024:data<=16'd8152;
      4025:data<=16'd8862;
      4026:data<=16'd8382;
      4027:data<=16'd8022;
      4028:data<=16'd7089;
      4029:data<=16'd6335;
      4030:data<=16'd6297;
      4031:data<=16'd5574;
      4032:data<=16'd4833;
      4033:data<=16'd3999;
      4034:data<=16'd3574;
      4035:data<=16'd3818;
      4036:data<=16'd2883;
      4037:data<=16'd2279;
      4038:data<=16'd2206;
      4039:data<=16'd1351;
      4040:data<=16'd1292;
      4041:data<=16'd396;
      4042:data<=-16'd264;
      4043:data<=16'd12;
      4044:data<=-16'd7009;
      4045:data<=-16'd16882;
      4046:data<=-16'd17823;
      4047:data<=-16'd15945;
      4048:data<=-16'd16666;
      4049:data<=-16'd16108;
      4050:data<=-16'd15564;
      4051:data<=-16'd15643;
      4052:data<=-16'd14971;
      4053:data<=-16'd14704;
      4054:data<=-16'd14784;
      4055:data<=-16'd14651;
      4056:data<=-16'd14114;
      4057:data<=-16'd13529;
      4058:data<=-16'd13054;
      4059:data<=-16'd12719;
      4060:data<=-16'd13640;
      4061:data<=-16'd13940;
      4062:data<=-16'd14490;
      4063:data<=-16'd18615;
      4064:data<=-16'd20416;
      4065:data<=-16'd18565;
      4066:data<=-16'd18909;
      4067:data<=-16'd18674;
      4068:data<=-16'd17725;
      4069:data<=-16'd17744;
      4070:data<=-16'd15575;
      4071:data<=-16'd15154;
      4072:data<=-16'd16278;
      4073:data<=-16'd14545;
      4074:data<=-16'd14270;
      4075:data<=-16'd14319;
      4076:data<=-16'd13490;
      4077:data<=-16'd15391;
      4078:data<=-16'd15258;
      4079:data<=-16'd13332;
      4080:data<=-16'd13335;
      4081:data<=-16'd12577;
      4082:data<=-16'd12478;
      4083:data<=-16'd11433;
      4084:data<=-16'd9632;
      4085:data<=-16'd11265;
      4086:data<=-16'd6032;
      4087:data<=16'd5145;
      4088:data<=16'd6586;
      4089:data<=16'd4541;
      4090:data<=16'd5888;
      4091:data<=16'd4864;
      4092:data<=16'd4640;
      4093:data<=16'd5121;
      4094:data<=16'd3051;
      4095:data<=16'd2684;
      4096:data<=16'd3353;
      4097:data<=16'd2869;
      4098:data<=16'd2675;
      4099:data<=16'd2165;
      4100:data<=16'd1595;
      4101:data<=16'd1668;
      4102:data<=16'd2082;
      4103:data<=16'd2296;
      4104:data<=16'd1770;
      4105:data<=16'd1788;
      4106:data<=16'd1977;
      4107:data<=16'd1439;
      4108:data<=16'd1814;
      4109:data<=16'd2493;
      4110:data<=16'd1651;
      4111:data<=-16'd174;
      4112:data<=16'd388;
      4113:data<=16'd4731;
      4114:data<=16'd7074;
      4115:data<=16'd6008;
      4116:data<=16'd5785;
      4117:data<=16'd5259;
      4118:data<=16'd5116;
      4119:data<=16'd5993;
      4120:data<=16'd4813;
      4121:data<=16'd4369;
      4122:data<=16'd4599;
      4123:data<=16'd3583;
      4124:data<=16'd4469;
      4125:data<=16'd3609;
      4126:data<=16'd1956;
      4127:data<=16'd4012;
      4128:data<=-16'd1363;
      4129:data<=-16'd12994;
      4130:data<=-16'd15001;
      4131:data<=-16'd12381;
      4132:data<=-16'd13226;
      4133:data<=-16'd12921;
      4134:data<=-16'd12232;
      4135:data<=-16'd12613;
      4136:data<=-16'd11737;
      4137:data<=-16'd10571;
      4138:data<=-16'd10217;
      4139:data<=-16'd10310;
      4140:data<=-16'd9969;
      4141:data<=-16'd8851;
      4142:data<=-16'd8000;
      4143:data<=-16'd8084;
      4144:data<=-16'd9163;
      4145:data<=-16'd9432;
      4146:data<=-16'd8232;
      4147:data<=-16'd8232;
      4148:data<=-16'd8661;
      4149:data<=-16'd7968;
      4150:data<=-16'd7787;
      4151:data<=-16'd7835;
      4152:data<=-16'd7567;
      4153:data<=-16'd7103;
      4154:data<=-16'd6320;
      4155:data<=-16'd6159;
      4156:data<=-16'd5786;
      4157:data<=-16'd5356;
      4158:data<=-16'd5383;
      4159:data<=-16'd4164;
      4160:data<=-16'd4258;
      4161:data<=-16'd5735;
      4162:data<=-16'd5861;
      4163:data<=-16'd8686;
      4164:data<=-16'd11547;
      4165:data<=-16'd10169;
      4166:data<=-16'd10272;
      4167:data<=-16'd9621;
      4168:data<=-16'd7841;
      4169:data<=-16'd10040;
      4170:data<=-16'd4946;
      4171:data<=16'd7415;
      4172:data<=16'd10182;
      4173:data<=16'd7762;
      4174:data<=16'd8419;
      4175:data<=16'd8002;
      4176:data<=16'd7685;
      4177:data<=16'd7507;
      4178:data<=16'd5938;
      4179:data<=16'd5486;
      4180:data<=16'd5332;
      4181:data<=16'd5385;
      4182:data<=16'd5905;
      4183:data<=16'd5375;
      4184:data<=16'd5172;
      4185:data<=16'd5482;
      4186:data<=16'd5915;
      4187:data<=16'd6052;
      4188:data<=16'd5004;
      4189:data<=16'd5658;
      4190:data<=16'd6452;
      4191:data<=16'd4840;
      4192:data<=16'd5280;
      4193:data<=16'd5982;
      4194:data<=16'd4143;
      4195:data<=16'd3439;
      4196:data<=16'd2857;
      4197:data<=16'd2390;
      4198:data<=16'd3565;
      4199:data<=16'd3750;
      4200:data<=16'd3721;
      4201:data<=16'd3691;
      4202:data<=16'd3303;
      4203:data<=16'd4344;
      4204:data<=16'd4106;
      4205:data<=16'd2981;
      4206:data<=16'd3042;
      4207:data<=16'd2500;
      4208:data<=16'd3209;
      4209:data<=16'd3240;
      4210:data<=16'd1703;
      4211:data<=16'd2737;
      4212:data<=-16'd1548;
      4213:data<=-16'd10261;
      4214:data<=-16'd9317;
      4215:data<=-16'd5708;
      4216:data<=-16'd7221;
      4217:data<=-16'd6420;
      4218:data<=-16'd5221;
      4219:data<=-16'd5799;
      4220:data<=-16'd4754;
      4221:data<=-16'd4502;
      4222:data<=-16'd4905;
      4223:data<=-16'd4155;
      4224:data<=-16'd3697;
      4225:data<=-16'd3294;
      4226:data<=-16'd2569;
      4227:data<=-16'd2535;
      4228:data<=-16'd3908;
      4229:data<=-16'd4534;
      4230:data<=-16'd3228;
      4231:data<=-16'd3251;
      4232:data<=-16'd3368;
      4233:data<=-16'd2173;
      4234:data<=-16'd2905;
      4235:data<=-16'd3148;
      4236:data<=-16'd1908;
      4237:data<=-16'd1847;
      4238:data<=-16'd1061;
      4239:data<=-16'd726;
      4240:data<=-16'd1566;
      4241:data<=-16'd1080;
      4242:data<=-16'd828;
      4243:data<=-16'd443;
      4244:data<=-16'd569;
      4245:data<=-16'd2391;
      4246:data<=-16'd1700;
      4247:data<=-16'd667;
      4248:data<=-16'd1121;
      4249:data<=-16'd68;
      4250:data<=-16'd588;
      4251:data<=-16'd337;
      4252:data<=16'd1184;
      4253:data<=-16'd1249;
      4254:data<=16'd2975;
      4255:data<=16'd14804;
      4256:data<=16'd17776;
      4257:data<=16'd15267;
      4258:data<=16'd15647;
      4259:data<=16'd15426;
      4260:data<=16'd14386;
      4261:data<=16'd13101;
      4262:data<=16'd12264;
      4263:data<=16'd10540;
      4264:data<=16'd5862;
      4265:data<=16'd4670;
      4266:data<=16'd6335;
      4267:data<=16'd5054;
      4268:data<=16'd4681;
      4269:data<=16'd4999;
      4270:data<=16'd4514;
      4271:data<=16'd5404;
      4272:data<=16'd4937;
      4273:data<=16'd4364;
      4274:data<=16'd4828;
      4275:data<=16'd4067;
      4276:data<=16'd5013;
      4277:data<=16'd5002;
      4278:data<=16'd1927;
      4279:data<=16'd1638;
      4280:data<=16'd2299;
      4281:data<=16'd1950;
      4282:data<=16'd2960;
      4283:data<=16'd3180;
      4284:data<=16'd2954;
      4285:data<=16'd2937;
      4286:data<=16'd2616;
      4287:data<=16'd3146;
      4288:data<=16'd2487;
      4289:data<=16'd1927;
      4290:data<=16'd2620;
      4291:data<=16'd1765;
      4292:data<=16'd2035;
      4293:data<=16'd2099;
      4294:data<=16'd1083;
      4295:data<=16'd3516;
      4296:data<=-16'd58;
      4297:data<=-16'd11238;
      4298:data<=-16'd14002;
      4299:data<=-16'd11112;
      4300:data<=-16'd11370;
      4301:data<=-16'd10809;
      4302:data<=-16'd10173;
      4303:data<=-16'd10389;
      4304:data<=-16'd9711;
      4305:data<=-16'd9635;
      4306:data<=-16'd9036;
      4307:data<=-16'd7940;
      4308:data<=-16'd7750;
      4309:data<=-16'd7241;
      4310:data<=-16'd6017;
      4311:data<=-16'd4660;
      4312:data<=-16'd4335;
      4313:data<=-16'd2370;
      4314:data<=16'd2863;
      4315:data<=16'd4484;
      4316:data<=16'd3242;
      4317:data<=16'd4338;
      4318:data<=16'd3897;
      4319:data<=16'd3210;
      4320:data<=16'd4385;
      4321:data<=16'd3635;
      4322:data<=16'd3560;
      4323:data<=16'd4473;
      4324:data<=16'd3808;
      4325:data<=16'd3830;
      4326:data<=16'd3714;
      4327:data<=16'd4396;
      4328:data<=16'd6802;
      4329:data<=16'd6946;
      4330:data<=16'd6707;
      4331:data<=16'd7147;
      4332:data<=16'd6745;
      4333:data<=16'd7494;
      4334:data<=16'd7006;
      4335:data<=16'd6058;
      4336:data<=16'd6361;
      4337:data<=16'd4240;
      4338:data<=16'd7841;
      4339:data<=16'd19086;
      4340:data<=16'd22551;
      4341:data<=16'd19845;
      4342:data<=16'd19980;
      4343:data<=16'd19334;
      4344:data<=16'd18880;
      4345:data<=16'd20131;
      4346:data<=16'd19579;
      4347:data<=16'd18425;
      4348:data<=16'd17794;
      4349:data<=16'd17238;
      4350:data<=16'd16968;
      4351:data<=16'd16196;
      4352:data<=16'd15258;
      4353:data<=16'd14545;
      4354:data<=16'd14272;
      4355:data<=16'd14299;
      4356:data<=16'd13468;
      4357:data<=16'd12825;
      4358:data<=16'd12798;
      4359:data<=16'd12129;
      4360:data<=16'd11559;
      4361:data<=16'd12175;
      4362:data<=16'd13308;
      4363:data<=16'd11085;
      4364:data<=16'd5615;
      4365:data<=16'd4111;
      4366:data<=16'd5515;
      4367:data<=16'd4871;
      4368:data<=16'd4739;
      4369:data<=16'd4578;
      4370:data<=16'd3695;
      4371:data<=16'd4262;
      4372:data<=16'd3833;
      4373:data<=16'd3107;
      4374:data<=16'd2934;
      4375:data<=16'd1579;
      4376:data<=16'd2130;
      4377:data<=16'd2403;
      4378:data<=16'd1485;
      4379:data<=16'd4285;
      4380:data<=16'd1510;
      4381:data<=-16'd9785;
      4382:data<=-16'd13890;
      4383:data<=-16'd11236;
      4384:data<=-16'd11336;
      4385:data<=-16'd11395;
      4386:data<=-16'd10487;
      4387:data<=-16'd10489;
      4388:data<=-16'd10445;
      4389:data<=-16'd10317;
      4390:data<=-16'd9793;
      4391:data<=-16'd9464;
      4392:data<=-16'd9494;
      4393:data<=-16'd8804;
      4394:data<=-16'd7837;
      4395:data<=-16'd6369;
      4396:data<=-16'd5551;
      4397:data<=-16'd6240;
      4398:data<=-16'd5623;
      4399:data<=-16'd4602;
      4400:data<=-16'd4965;
      4401:data<=-16'd4893;
      4402:data<=-16'd4939;
      4403:data<=-16'd5285;
      4404:data<=-16'd4951;
      4405:data<=-16'd4737;
      4406:data<=-16'd4338;
      4407:data<=-16'd4073;
      4408:data<=-16'd4279;
      4409:data<=-16'd4234;
      4410:data<=-16'd4214;
      4411:data<=-16'd3453;
      4412:data<=-16'd2528;
      4413:data<=-16'd789;
      4414:data<=16'd3788;
      4415:data<=16'd5735;
      4416:data<=16'd4645;
      4417:data<=16'd5771;
      4418:data<=16'd4939;
      4419:data<=16'd3962;
      4420:data<=16'd5533;
      4421:data<=16'd2964;
      4422:data<=16'd5304;
      4423:data<=16'd16971;
      4424:data<=16'd21123;
      4425:data<=16'd18662;
      4426:data<=16'd18644;
      4427:data<=16'd17666;
      4428:data<=16'd17723;
      4429:data<=16'd18760;
      4430:data<=16'd17638;
      4431:data<=16'd17153;
      4432:data<=16'd15729;
      4433:data<=16'd14122;
      4434:data<=16'd14744;
      4435:data<=16'd13620;
      4436:data<=16'd12055;
      4437:data<=16'd11712;
      4438:data<=16'd10909;
      4439:data<=16'd11159;
      4440:data<=16'd10602;
      4441:data<=16'd9327;
      4442:data<=16'd9599;
      4443:data<=16'd8777;
      4444:data<=16'd8719;
      4445:data<=16'd10108;
      4446:data<=16'd9368;
      4447:data<=16'd8860;
      4448:data<=16'd8540;
      4449:data<=16'd6998;
      4450:data<=16'd6623;
      4451:data<=16'd6216;
      4452:data<=16'd5833;
      4453:data<=16'd6102;
      4454:data<=16'd5385;
      4455:data<=16'd5043;
      4456:data<=16'd4291;
      4457:data<=16'd3022;
      4458:data<=16'd3110;
      4459:data<=16'd2231;
      4460:data<=16'd1551;
      4461:data<=16'd2229;
      4462:data<=16'd2805;
      4463:data<=16'd3892;
      4464:data<=-16'd1823;
      4465:data<=-16'd14436;
      4466:data<=-16'd19194;
      4467:data<=-16'd17141;
      4468:data<=-16'd16923;
      4469:data<=-16'd16337;
      4470:data<=-16'd15978;
      4471:data<=-16'd16495;
      4472:data<=-16'd16104;
      4473:data<=-16'd15770;
      4474:data<=-16'd14678;
      4475:data<=-16'd14045;
      4476:data<=-16'd14619;
      4477:data<=-16'd13832;
      4478:data<=-16'd12622;
      4479:data<=-16'd11217;
      4480:data<=-16'd10073;
      4481:data<=-16'd10783;
      4482:data<=-16'd10480;
      4483:data<=-16'd9693;
      4484:data<=-16'd10383;
      4485:data<=-16'd10082;
      4486:data<=-16'd9315;
      4487:data<=-16'd9009;
      4488:data<=-16'd8790;
      4489:data<=-16'd8992;
      4490:data<=-16'd8320;
      4491:data<=-16'd7683;
      4492:data<=-16'd7514;
      4493:data<=-16'd7112;
      4494:data<=-16'd7708;
      4495:data<=-16'd6670;
      4496:data<=-16'd4540;
      4497:data<=-16'd4773;
      4498:data<=-16'd4306;
      4499:data<=-16'd4190;
      4500:data<=-16'd5224;
      4501:data<=-16'd3899;
      4502:data<=-16'd4278;
      4503:data<=-16'd5203;
      4504:data<=-16'd3744;
      4505:data<=-16'd5362;
      4506:data<=-16'd3028;
      4507:data<=16'd7533;
      4508:data<=16'd12666;
      4509:data<=16'd11015;
      4510:data<=16'd10478;
      4511:data<=16'd10856;
      4512:data<=16'd11629;
      4513:data<=16'd12536;
      4514:data<=16'd14113;
      4515:data<=16'd15746;
      4516:data<=16'd14230;
      4517:data<=16'd12478;
      4518:data<=16'd12333;
      4519:data<=16'd11314;
      4520:data<=16'd10839;
      4521:data<=16'd10716;
      4522:data<=16'd10019;
      4523:data<=16'd9568;
      4524:data<=16'd8437;
      4525:data<=16'd8310;
      4526:data<=16'd8813;
      4527:data<=16'd7421;
      4528:data<=16'd7582;
      4529:data<=16'd9163;
      4530:data<=16'd8419;
      4531:data<=16'd7365;
      4532:data<=16'd7075;
      4533:data<=16'd6285;
      4534:data<=16'd5275;
      4535:data<=16'd4742;
      4536:data<=16'd5031;
      4537:data<=16'd4514;
      4538:data<=16'd3519;
      4539:data<=16'd3526;
      4540:data<=16'd2613;
      4541:data<=16'd1921;
      4542:data<=16'd2209;
      4543:data<=16'd892;
      4544:data<=16'd934;
      4545:data<=16'd2396;
      4546:data<=16'd1945;
      4547:data<=16'd2789;
      4548:data<=16'd926;
      4549:data<=-16'd8661;
      4550:data<=-16'd15138;
      4551:data<=-16'd14152;
      4552:data<=-16'd13720;
      4553:data<=-16'd13831;
      4554:data<=-16'd12690;
      4555:data<=-16'd12780;
      4556:data<=-16'd13336;
      4557:data<=-16'd13305;
      4558:data<=-16'd12731;
      4559:data<=-16'd11521;
      4560:data<=-16'd11194;
      4561:data<=-16'd11632;
      4562:data<=-16'd11063;
      4563:data<=-16'd10610;
      4564:data<=-16'd12460;
      4565:data<=-16'd14822;
      4566:data<=-16'd14619;
      4567:data<=-16'd13829;
      4568:data<=-16'd14345;
      4569:data<=-16'd13888;
      4570:data<=-16'd13173;
      4571:data<=-16'd13338;
      4572:data<=-16'd12354;
      4573:data<=-16'd11403;
      4574:data<=-16'd11862;
      4575:data<=-16'd11952;
      4576:data<=-16'd11112;
      4577:data<=-16'd10226;
      4578:data<=-16'd10995;
      4579:data<=-16'd12609;
      4580:data<=-16'd12289;
      4581:data<=-16'd11600;
      4582:data<=-16'd11420;
      4583:data<=-16'd10590;
      4584:data<=-16'd10199;
      4585:data<=-16'd9502;
      4586:data<=-16'd8889;
      4587:data<=-16'd9000;
      4588:data<=-16'd7856;
      4589:data<=-16'd8234;
      4590:data<=-16'd7228;
      4591:data<=16'd1814;
      4592:data<=16'd9048;
      4593:data<=16'd8410;
      4594:data<=16'd7967;
      4595:data<=16'd7116;
      4596:data<=16'd4631;
      4597:data<=16'd4593;
      4598:data<=16'd5039;
      4599:data<=16'd4887;
      4600:data<=16'd4484;
      4601:data<=16'd3381;
      4602:data<=16'd3677;
      4603:data<=16'd3856;
      4604:data<=16'd2689;
      4605:data<=16'd2491;
      4606:data<=16'd2487;
      4607:data<=16'd2288;
      4608:data<=16'd2244;
      4609:data<=16'd1867;
      4610:data<=16'd2273;
      4611:data<=16'd2159;
      4612:data<=16'd538;
      4613:data<=-16'd173;
      4614:data<=16'd870;
      4615:data<=16'd2999;
      4616:data<=16'd4071;
      4617:data<=16'd2984;
      4618:data<=16'd2341;
      4619:data<=16'd2698;
      4620:data<=16'd2996;
      4621:data<=16'd2999;
      4622:data<=16'd2397;
      4623:data<=16'd2306;
      4624:data<=16'd2416;
      4625:data<=16'd2187;
      4626:data<=16'd2370;
      4627:data<=16'd1521;
      4628:data<=16'd546;
      4629:data<=16'd120;
      4630:data<=-16'd1331;
      4631:data<=-16'd456;
      4632:data<=-16'd602;
      4633:data<=-16'd9222;
      4634:data<=-16'd17459;
      4635:data<=-16'd17443;
      4636:data<=-16'd15828;
      4637:data<=-16'd15503;
      4638:data<=-16'd14636;
      4639:data<=-16'd14046;
      4640:data<=-16'd14045;
      4641:data<=-16'd13919;
      4642:data<=-16'd12900;
      4643:data<=-16'd11583;
      4644:data<=-16'd11004;
      4645:data<=-16'd11254;
      4646:data<=-16'd12325;
      4647:data<=-16'd12411;
      4648:data<=-16'd11104;
      4649:data<=-16'd10640;
      4650:data<=-16'd10451;
      4651:data<=-16'd10143;
      4652:data<=-16'd10460;
      4653:data<=-16'd9814;
      4654:data<=-16'd8522;
      4655:data<=-16'd8316;
      4656:data<=-16'd8398;
      4657:data<=-16'd7662;
      4658:data<=-16'd6743;
      4659:data<=-16'd6542;
      4660:data<=-16'd5871;
      4661:data<=-16'd5265;
      4662:data<=-16'd6561;
      4663:data<=-16'd7188;
      4664:data<=-16'd7852;
      4665:data<=-16'd10947;
      4666:data<=-16'd11546;
      4667:data<=-16'd10099;
      4668:data<=-16'd10288;
      4669:data<=-16'd8601;
      4670:data<=-16'd7297;
      4671:data<=-16'd8308;
      4672:data<=-16'd6899;
      4673:data<=-16'd6810;
      4674:data<=-16'd7042;
      4675:data<=16'd1055;
      4676:data<=16'd9893;
      4677:data<=16'd10878;
      4678:data<=16'd9586;
      4679:data<=16'd8508;
      4680:data<=16'd7150;
      4681:data<=16'd7009;
      4682:data<=16'd7134;
      4683:data<=16'd7427;
      4684:data<=16'd7363;
      4685:data<=16'd5962;
      4686:data<=16'd5632;
      4687:data<=16'd6457;
      4688:data<=16'd6461;
      4689:data<=16'd5970;
      4690:data<=16'd5301;
      4691:data<=16'd5278;
      4692:data<=16'd5771;
      4693:data<=16'd5682;
      4694:data<=16'd6158;
      4695:data<=16'd5651;
      4696:data<=16'd3043;
      4697:data<=16'd2475;
      4698:data<=16'd3228;
      4699:data<=16'd2514;
      4700:data<=16'd2517;
      4701:data<=16'd2576;
      4702:data<=16'd1865;
      4703:data<=16'd2270;
      4704:data<=16'd2485;
      4705:data<=16'd2282;
      4706:data<=16'd2514;
      4707:data<=16'd2212;
      4708:data<=16'd2384;
      4709:data<=16'd2820;
      4710:data<=16'd2464;
      4711:data<=16'd2458;
      4712:data<=16'd2085;
      4713:data<=16'd858;
      4714:data<=16'd936;
      4715:data<=16'd4109;
      4716:data<=16'd6513;
      4717:data<=-16'd129;
      4718:data<=-16'd10634;
      4719:data<=-16'd12533;
      4720:data<=-16'd10296;
      4721:data<=-16'd10126;
      4722:data<=-16'd8909;
      4723:data<=-16'd8495;
      4724:data<=-16'd9092;
      4725:data<=-16'd8150;
      4726:data<=-16'd7714;
      4727:data<=-16'd7100;
      4728:data<=-16'd6475;
      4729:data<=-16'd7753;
      4730:data<=-16'd8150;
      4731:data<=-16'd7221;
      4732:data<=-16'd6626;
      4733:data<=-16'd6263;
      4734:data<=-16'd6269;
      4735:data<=-16'd5777;
      4736:data<=-16'd5653;
      4737:data<=-16'd5982;
      4738:data<=-16'd4642;
      4739:data<=-16'd3983;
      4740:data<=-16'd4302;
      4741:data<=-16'd3181;
      4742:data<=-16'd2769;
      4743:data<=-16'd2823;
      4744:data<=-16'd2052;
      4745:data<=-16'd2376;
      4746:data<=-16'd3406;
      4747:data<=-16'd4012;
      4748:data<=-16'd3662;
      4749:data<=-16'd2813;
      4750:data<=-16'd2828;
      4751:data<=-16'd2505;
      4752:data<=-16'd2127;
      4753:data<=-16'd2065;
      4754:data<=-16'd1172;
      4755:data<=-16'd1081;
      4756:data<=-16'd315;
      4757:data<=16'd118;
      4758:data<=-16'd2205;
      4759:data<=16'd3360;
      4760:data<=16'd15641;
      4761:data<=16'd17631;
      4762:data<=16'd13490;
      4763:data<=16'd12730;
      4764:data<=16'd10566;
      4765:data<=16'd7903;
      4766:data<=16'd7256;
      4767:data<=16'd6695;
      4768:data<=16'd6878;
      4769:data<=16'd6907;
      4770:data<=16'd6801;
      4771:data<=16'd7301;
      4772:data<=16'd6710;
      4773:data<=16'd6152;
      4774:data<=16'd6255;
      4775:data<=16'd5941;
      4776:data<=16'd5821;
      4777:data<=16'd5950;
      4778:data<=16'd6202;
      4779:data<=16'd5215;
      4780:data<=16'd2972;
      4781:data<=16'd2610;
      4782:data<=16'd3062;
      4783:data<=16'd2917;
      4784:data<=16'd3239;
      4785:data<=16'd2690;
      4786:data<=16'd2332;
      4787:data<=16'd3077;
      4788:data<=16'd3157;
      4789:data<=16'd3385;
      4790:data<=16'd3328;
      4791:data<=16'd3075;
      4792:data<=16'd3529;
      4793:data<=16'd2955;
      4794:data<=16'd3306;
      4795:data<=16'd3498;
      4796:data<=16'd693;
      4797:data<=16'd191;
      4798:data<=16'd605;
      4799:data<=16'd33;
      4800:data<=16'd2576;
      4801:data<=-16'd2008;
      4802:data<=-16'd14340;
      4803:data<=-16'd16903;
      4804:data<=-16'd13694;
      4805:data<=-16'd14048;
      4806:data<=-16'd12956;
      4807:data<=-16'd11973;
      4808:data<=-16'd11794;
      4809:data<=-16'd10358;
      4810:data<=-16'd10722;
      4811:data<=-16'd10208;
      4812:data<=-16'd9333;
      4813:data<=-16'd11470;
      4814:data<=-16'd10279;
      4815:data<=-16'd5961;
      4816:data<=-16'd4689;
      4817:data<=-16'd4325;
      4818:data<=-16'd3620;
      4819:data<=-16'd3779;
      4820:data<=-16'd3665;
      4821:data<=-16'd3142;
      4822:data<=-16'd2543;
      4823:data<=-16'd2134;
      4824:data<=-16'd1785;
      4825:data<=-16'd1475;
      4826:data<=-16'd1580;
      4827:data<=-16'd1036;
      4828:data<=-16'd490;
      4829:data<=-16'd726;
      4830:data<=-16'd340;
      4831:data<=-16'd129;
      4832:data<=-16'd127;
      4833:data<=16'd411;
      4834:data<=16'd317;
      4835:data<=16'd338;
      4836:data<=16'd350;
      4837:data<=16'd599;
      4838:data<=16'd2044;
      4839:data<=16'd1691;
      4840:data<=16'd1559;
      4841:data<=16'd2760;
      4842:data<=16'd1206;
      4843:data<=16'd5421;
      4844:data<=16'd16732;
      4845:data<=16'd19866;
      4846:data<=16'd17885;
      4847:data<=16'd19321;
      4848:data<=16'd18873;
      4849:data<=16'd17681;
      4850:data<=16'd17673;
      4851:data<=16'd16728;
      4852:data<=16'd16910;
      4853:data<=16'd16434;
      4854:data<=16'd15394;
      4855:data<=16'd16211;
      4856:data<=16'd15174;
      4857:data<=16'd13333;
      4858:data<=16'd13429;
      4859:data<=16'd13294;
      4860:data<=16'd13130;
      4861:data<=16'd12411;
      4862:data<=16'd11690;
      4863:data<=16'd12821;
      4864:data<=16'd12126;
      4865:data<=16'd9332;
      4866:data<=16'd7952;
      4867:data<=16'd7413;
      4868:data<=16'd7150;
      4869:data<=16'd6764;
      4870:data<=16'd6244;
      4871:data<=16'd6390;
      4872:data<=16'd6100;
      4873:data<=16'd5724;
      4874:data<=16'd5532;
      4875:data<=16'd5104;
      4876:data<=16'd5336;
      4877:data<=16'd4831;
      4878:data<=16'd4259;
      4879:data<=16'd5175;
      4880:data<=16'd5456;
      4881:data<=16'd5796;
      4882:data<=16'd5454;
      4883:data<=16'd4438;
      4884:data<=16'd6281;
      4885:data<=16'd2479;
      4886:data<=-16'd9283;
      4887:data<=-16'd13186;
      4888:data<=-16'd10207;
      4889:data<=-16'd10596;
      4890:data<=-16'd10217;
      4891:data<=-16'd8924;
      4892:data<=-16'd9401;
      4893:data<=-16'd8718;
      4894:data<=-16'd8355;
      4895:data<=-16'd8595;
      4896:data<=-16'd7429;
      4897:data<=-16'd6473;
      4898:data<=-16'd5594;
      4899:data<=-16'd4645;
      4900:data<=-16'd4695;
      4901:data<=-16'd4730;
      4902:data<=-16'd4687;
      4903:data<=-16'd4726;
      4904:data<=-16'd4225;
      4905:data<=-16'd3824;
      4906:data<=-16'd3847;
      4907:data<=-16'd3833;
      4908:data<=-16'd3453;
      4909:data<=-16'd2822;
      4910:data<=-16'd2543;
      4911:data<=-16'd2572;
      4912:data<=-16'd2171;
      4913:data<=-16'd961;
      4914:data<=16'd488;
      4915:data<=16'd2311;
      4916:data<=16'd4329;
      4917:data<=16'd4259;
      4918:data<=16'd3676;
      4919:data<=16'd4696;
      4920:data<=16'd4099;
      4921:data<=16'd3436;
      4922:data<=16'd4549;
      4923:data<=16'd3847;
      4924:data<=16'd4220;
      4925:data<=16'd4927;
      4926:data<=16'd2399;
      4927:data<=16'd7104;
      4928:data<=16'd18099;
      4929:data<=16'd20800;
      4930:data<=16'd19378;
      4931:data<=16'd20084;
      4932:data<=16'd19139;
      4933:data<=16'd18668;
      4934:data<=16'd18172;
      4935:data<=16'd16146;
      4936:data<=16'd16261;
      4937:data<=16'd16161;
      4938:data<=16'd14694;
      4939:data<=16'd14572;
      4940:data<=16'd13728;
      4941:data<=16'd12445;
      4942:data<=16'd12243;
      4943:data<=16'd11671;
      4944:data<=16'd11185;
      4945:data<=16'd10813;
      4946:data<=16'd10619;
      4947:data<=16'd11259;
      4948:data<=16'd11291;
      4949:data<=16'd10856;
      4950:data<=16'd10314;
      4951:data<=16'd9433;
      4952:data<=16'd9312;
      4953:data<=16'd8728;
      4954:data<=16'd7506;
      4955:data<=16'd7339;
      4956:data<=16'd7157;
      4957:data<=16'd6949;
      4958:data<=16'd6889;
      4959:data<=16'd6147;
      4960:data<=16'd5598;
      4961:data<=16'd4807;
      4962:data<=16'd4413;
      4963:data<=16'd5348;
      4964:data<=16'd5171;
      4965:data<=16'd3697;
      4966:data<=16'd1271;
      4967:data<=-16'd279;
      4968:data<=16'd1254;
      4969:data<=-16'd2849;
      4970:data<=-16'd13515;
      4971:data<=-16'd17004;
      4972:data<=-16'd15117;
      4973:data<=-16'd15426;
      4974:data<=-16'd14434;
      4975:data<=-16'd13565;
      4976:data<=-16'd13893;
      4977:data<=-16'd13073;
      4978:data<=-16'd13576;
      4979:data<=-16'd13289;
      4980:data<=-16'd10945;
      4981:data<=-16'd10707;
      4982:data<=-16'd10866;
      4983:data<=-16'd9985;
      4984:data<=-16'd9577;
      4985:data<=-16'd8965;
      4986:data<=-16'd9044;
      4987:data<=-16'd9418;
      4988:data<=-16'd8757;
      4989:data<=-16'd8302;
      4990:data<=-16'd7934;
      4991:data<=-16'd7844;
      4992:data<=-16'd8290;
      4993:data<=-16'd7753;
      4994:data<=-16'd7009;
      4995:data<=-16'd6957;
      4996:data<=-16'd6391;
      4997:data<=-16'd4902;
      4998:data<=-16'd3877;
      4999:data<=-16'd4235;
      5000:data<=-16'd4258;
      5001:data<=-16'd4073;
      5002:data<=-16'd4504;
      5003:data<=-16'd3653;
      5004:data<=-16'd3454;
      5005:data<=-16'd4243;
      5006:data<=-16'd3046;
      5007:data<=-16'd3080;
      5008:data<=-16'd3533;
      5009:data<=-16'd2243;
      5010:data<=-16'd3348;
      5011:data<=-16'd53;
      5012:data<=16'd10519;
      5013:data<=16'd14643;
      5014:data<=16'd13279;
      5015:data<=16'd15524;
      5016:data<=16'd17132;
      5017:data<=16'd16425;
      5018:data<=16'd15960;
      5019:data<=16'd15214;
      5020:data<=16'd14710;
      5021:data<=16'd13899;
      5022:data<=16'd12859;
      5023:data<=16'd12698;
      5024:data<=16'd12267;
      5025:data<=16'd11391;
      5026:data<=16'd10557;
      5027:data<=16'd9928;
      5028:data<=16'd9714;
      5029:data<=16'd9643;
      5030:data<=16'd10241;
      5031:data<=16'd10507;
      5032:data<=16'd9747;
      5033:data<=16'd9517;
      5034:data<=16'd9098;
      5035:data<=16'd8349;
      5036:data<=16'd7773;
      5037:data<=16'd6601;
      5038:data<=16'd6440;
      5039:data<=16'd6191;
      5040:data<=16'd4598;
      5041:data<=16'd4717;
      5042:data<=16'd5002;
      5043:data<=16'd4452;
      5044:data<=16'd4411;
      5045:data<=16'd2702;
      5046:data<=16'd2826;
      5047:data<=16'd5585;
      5048:data<=16'd4881;
      5049:data<=16'd3900;
      5050:data<=16'd3903;
      5051:data<=16'd2481;
      5052:data<=16'd3519;
      5053:data<=16'd387;
      5054:data<=-16'd10266;
      5055:data<=-16'd14584;
      5056:data<=-16'd12683;
      5057:data<=-16'd13123;
      5058:data<=-16'd12759;
      5059:data<=-16'd12105;
      5060:data<=-16'd12719;
      5061:data<=-16'd12019;
      5062:data<=-16'd12132;
      5063:data<=-16'd11506;
      5064:data<=-16'd8501;
      5065:data<=-16'd9404;
      5066:data<=-16'd12906;
      5067:data<=-16'd12690;
      5068:data<=-16'd11705;
      5069:data<=-16'd12261;
      5070:data<=-16'd11752;
      5071:data<=-16'd11194;
      5072:data<=-16'd11347;
      5073:data<=-16'd10596;
      5074:data<=-16'd10228;
      5075:data<=-16'd10611;
      5076:data<=-16'd10069;
      5077:data<=-16'd9570;
      5078:data<=-16'd9241;
      5079:data<=-16'd8146;
      5080:data<=-16'd7413;
      5081:data<=-16'd6523;
      5082:data<=-16'd5374;
      5083:data<=-16'd5498;
      5084:data<=-16'd5441;
      5085:data<=-16'd5115;
      5086:data<=-16'd5365;
      5087:data<=-16'd4560;
      5088:data<=-16'd4369;
      5089:data<=-16'd4980;
      5090:data<=-16'd4023;
      5091:data<=-16'd4399;
      5092:data<=-16'd4974;
      5093:data<=-16'd3548;
      5094:data<=-16'd4303;
      5095:data<=-16'd1292;
      5096:data<=16'd9066;
      5097:data<=16'd13383;
      5098:data<=16'd11094;
      5099:data<=16'd11459;
      5100:data<=16'd11132;
      5101:data<=16'd9828;
      5102:data<=16'd10181;
      5103:data<=16'd9244;
      5104:data<=16'd8721;
      5105:data<=16'd8778;
      5106:data<=16'd7445;
      5107:data<=16'd7555;
      5108:data<=16'd7782;
      5109:data<=16'd6664;
      5110:data<=16'd6510;
      5111:data<=16'd6328;
      5112:data<=16'd6287;
      5113:data<=16'd6011;
      5114:data<=16'd4050;
      5115:data<=16'd4469;
      5116:data<=16'd7071;
      5117:data<=16'd7191;
      5118:data<=16'd6457;
      5119:data<=16'd6522;
      5120:data<=16'd5894;
      5121:data<=16'd4769;
      5122:data<=16'd4255;
      5123:data<=16'd4314;
      5124:data<=16'd3845;
      5125:data<=16'd3642;
      5126:data<=16'd4114;
      5127:data<=16'd3535;
      5128:data<=16'd2937;
      5129:data<=16'd2801;
      5130:data<=16'd1768;
      5131:data<=16'd587;
      5132:data<=-16'd318;
      5133:data<=-16'd99;
      5134:data<=16'd127;
      5135:data<=-16'd1090;
      5136:data<=-16'd409;
      5137:data<=-16'd2969;
      5138:data<=-16'd13177;
      5139:data<=-16'd18167;
      5140:data<=-16'd15770;
      5141:data<=-16'd15846;
      5142:data<=-16'd15676;
      5143:data<=-16'd14175;
      5144:data<=-16'd14255;
      5145:data<=-16'd13490;
      5146:data<=-16'd13603;
      5147:data<=-16'd14707;
      5148:data<=-16'd14245;
      5149:data<=-16'd14225;
      5150:data<=-16'd14010;
      5151:data<=-16'd13215;
      5152:data<=-16'd13204;
      5153:data<=-16'd12404;
      5154:data<=-16'd11755;
      5155:data<=-16'd11776;
      5156:data<=-16'd11097;
      5157:data<=-16'd10730;
      5158:data<=-16'd10161;
      5159:data<=-16'd9409;
      5160:data<=-16'd9313;
      5161:data<=-16'd8605;
      5162:data<=-16'd8147;
      5163:data<=-16'd8326;
      5164:data<=-16'd8502;
      5165:data<=-16'd10084;
      5166:data<=-16'd12296;
      5167:data<=-16'd13335;
      5168:data<=-16'd12977;
      5169:data<=-16'd12211;
      5170:data<=-16'd12093;
      5171:data<=-16'd11436;
      5172:data<=-16'd11016;
      5173:data<=-16'd11009;
      5174:data<=-16'd9313;
      5175:data<=-16'd9000;
      5176:data<=-16'd9420;
      5177:data<=-16'd7905;
      5178:data<=-16'd8428;
      5179:data<=-16'd5526;
      5180:data<=16'd3935;
      5181:data<=16'd7491;
      5182:data<=16'd5538;
      5183:data<=16'd5905;
      5184:data<=16'd5653;
      5185:data<=16'd5263;
      5186:data<=16'd5629;
      5187:data<=16'd5022;
      5188:data<=16'd5418;
      5189:data<=16'd5272;
      5190:data<=16'd4402;
      5191:data<=16'd5072;
      5192:data<=16'd5004;
      5193:data<=16'd4585;
      5194:data<=16'd4573;
      5195:data<=16'd3739;
      5196:data<=16'd3638;
      5197:data<=16'd3215;
      5198:data<=16'd1888;
      5199:data<=16'd1616;
      5200:data<=16'd1216;
      5201:data<=16'd876;
      5202:data<=16'd996;
      5203:data<=16'd517;
      5204:data<=16'd641;
      5205:data<=16'd593;
      5206:data<=16'd12;
      5207:data<=16'd262;
      5208:data<=16'd44;
      5209:data<=16'd170;
      5210:data<=16'd957;
      5211:data<=16'd608;
      5212:data<=16'd631;
      5213:data<=16'd56;
      5214:data<=-16'd1680;
      5215:data<=-16'd816;
      5216:data<=16'd1445;
      5217:data<=16'd2743;
      5218:data<=16'd3004;
      5219:data<=16'd2217;
      5220:data<=16'd2898;
      5221:data<=16'd967;
      5222:data<=-16'd7835;
      5223:data<=-16'd13728;
      5224:data<=-16'd12959;
      5225:data<=-16'd12369;
      5226:data<=-16'd11561;
      5227:data<=-16'd10548;
      5228:data<=-16'd11077;
      5229:data<=-16'd10326;
      5230:data<=-16'd10069;
      5231:data<=-16'd11693;
      5232:data<=-16'd11802;
      5233:data<=-16'd11462;
      5234:data<=-16'd11543;
      5235:data<=-16'd10458;
      5236:data<=-16'd9605;
      5237:data<=-16'd9359;
      5238:data<=-16'd8904;
      5239:data<=-16'd8329;
      5240:data<=-16'd7365;
      5241:data<=-16'd6931;
      5242:data<=-16'd6855;
      5243:data<=-16'd5953;
      5244:data<=-16'd5288;
      5245:data<=-16'd4875;
      5246:data<=-16'd4432;
      5247:data<=-16'd5213;
      5248:data<=-16'd6070;
      5249:data<=-16'd5829;
      5250:data<=-16'd5752;
      5251:data<=-16'd5958;
      5252:data<=-16'd5717;
      5253:data<=-16'd5172;
      5254:data<=-16'd4385;
      5255:data<=-16'd3447;
      5256:data<=-16'd3298;
      5257:data<=-16'd3607;
      5258:data<=-16'd2754;
      5259:data<=-16'd2137;
      5260:data<=-16'd2485;
      5261:data<=-16'd2015;
      5262:data<=-16'd2485;
      5263:data<=-16'd1315;
      5264:data<=16'd6525;
      5265:data<=16'd12023;
      5266:data<=16'd8974;
      5267:data<=16'd6457;
      5268:data<=16'd6757;
      5269:data<=16'd6279;
      5270:data<=16'd6501;
      5271:data<=16'd6552;
      5272:data<=16'd5968;
      5273:data<=16'd6217;
      5274:data<=16'd6120;
      5275:data<=16'd6065;
      5276:data<=16'd6261;
      5277:data<=16'd5576;
      5278:data<=16'd5319;
      5279:data<=16'd5454;
      5280:data<=16'd4479;
      5281:data<=16'd3034;
      5282:data<=16'd2532;
      5283:data<=16'd2813;
      5284:data<=16'd2279;
      5285:data<=16'd1645;
      5286:data<=16'd2123;
      5287:data<=16'd2281;
      5288:data<=16'd2420;
      5289:data<=16'd2722;
      5290:data<=16'd2030;
      5291:data<=16'd1894;
      5292:data<=16'd2396;
      5293:data<=16'd2405;
      5294:data<=16'd2638;
      5295:data<=16'd2578;
      5296:data<=16'd2241;
      5297:data<=16'd1415;
      5298:data<=-16'd291;
      5299:data<=-16'd557;
      5300:data<=-16'd211;
      5301:data<=-16'd491;
      5302:data<=16'd85;
      5303:data<=-16'd2;
      5304:data<=16'd165;
      5305:data<=-16'd667;
      5306:data<=-16'd8194;
      5307:data<=-16'd15057;
      5308:data<=-16'd14524;
      5309:data<=-16'd13946;
      5310:data<=-16'd14029;
      5311:data<=-16'd12631;
      5312:data<=-16'd12489;
      5313:data<=-16'd11506;
      5314:data<=-16'd11075;
      5315:data<=-16'd12742;
      5316:data<=-16'd10765;
      5317:data<=-16'd7194;
      5318:data<=-16'd6719;
      5319:data<=-16'd6228;
      5320:data<=-16'd5090;
      5321:data<=-16'd4849;
      5322:data<=-16'd4617;
      5323:data<=-16'd4065;
      5324:data<=-16'd3524;
      5325:data<=-16'd3189;
      5326:data<=-16'd2400;
      5327:data<=-16'd1850;
      5328:data<=-16'd2378;
      5329:data<=-16'd1888;
      5330:data<=-16'd1676;
      5331:data<=-16'd3322;
      5332:data<=-16'd3351;
      5333:data<=-16'd2464;
      5334:data<=-16'd2796;
      5335:data<=-16'd2460;
      5336:data<=-16'd2005;
      5337:data<=-16'd1911;
      5338:data<=-16'd1354;
      5339:data<=-16'd1004;
      5340:data<=-16'd652;
      5341:data<=-16'd731;
      5342:data<=-16'd622;
      5343:data<=16'd317;
      5344:data<=-16'd91;
      5345:data<=16'd12;
      5346:data<=16'd886;
      5347:data<=16'd741;
      5348:data<=16'd6018;
      5349:data<=16'd14098;
      5350:data<=16'd14613;
      5351:data<=16'd12951;
      5352:data<=16'd13637;
      5353:data<=16'd12748;
      5354:data<=16'd12684;
      5355:data<=16'd12951;
      5356:data<=16'd11753;
      5357:data<=16'd11993;
      5358:data<=16'd11796;
      5359:data<=16'd10916;
      5360:data<=16'd11295;
      5361:data<=16'd10658;
      5362:data<=16'd9828;
      5363:data<=16'd9565;
      5364:data<=16'd9135;
      5365:data<=16'd9577;
      5366:data<=16'd7733;
      5367:data<=16'd3753;
      5368:data<=16'd2743;
      5369:data<=16'd3074;
      5370:data<=16'd2666;
      5371:data<=16'd2839;
      5372:data<=16'd3063;
      5373:data<=16'd2958;
      5374:data<=16'd2473;
      5375:data<=16'd2232;
      5376:data<=16'd2344;
      5377:data<=16'd1891;
      5378:data<=16'd2291;
      5379:data<=16'd2773;
      5380:data<=16'd2385;
      5381:data<=16'd3518;
      5382:data<=16'd4538;
      5383:data<=16'd4352;
      5384:data<=16'd4347;
      5385:data<=16'd3753;
      5386:data<=16'd4005;
      5387:data<=16'd4121;
      5388:data<=16'd3585;
      5389:data<=16'd4408;
      5390:data<=-16'd1108;
      5391:data<=-16'd11385;
      5392:data<=-16'd12895;
      5393:data<=-16'd10701;
      5394:data<=-16'd11233;
      5395:data<=-16'd10050;
      5396:data<=-16'd9911;
      5397:data<=-16'd9514;
      5398:data<=-16'd6510;
      5399:data<=-16'd6132;
      5400:data<=-16'd5953;
      5401:data<=-16'd4690;
      5402:data<=-16'd5362;
      5403:data<=-16'd4855;
      5404:data<=-16'd3817;
      5405:data<=-16'd4027;
      5406:data<=-16'd3847;
      5407:data<=-16'd3905;
      5408:data<=-16'd3315;
      5409:data<=-16'd2616;
      5410:data<=-16'd2657;
      5411:data<=-16'd1792;
      5412:data<=-16'd1980;
      5413:data<=-16'd2044;
      5414:data<=-16'd320;
      5415:data<=16'd197;
      5416:data<=16'd2231;
      5417:data<=16'd5691;
      5418:data<=16'd6002;
      5419:data<=16'd5742;
      5420:data<=16'd5705;
      5421:data<=16'd5092;
      5422:data<=16'd5492;
      5423:data<=16'd5442;
      5424:data<=16'd5168;
      5425:data<=16'd4943;
      5426:data<=16'd4748;
      5427:data<=16'd5647;
      5428:data<=16'd5103;
      5429:data<=16'd5109;
      5430:data<=16'd5811;
      5431:data<=16'd4062;
      5432:data<=16'd10091;
      5433:data<=16'd21779;
      5434:data<=16'd22786;
      5435:data<=16'd19951;
      5436:data<=16'd20663;
      5437:data<=16'd18921;
      5438:data<=16'd17996;
      5439:data<=16'd18266;
      5440:data<=16'd16977;
      5441:data<=16'd16898;
      5442:data<=16'd16087;
      5443:data<=16'd15083;
      5444:data<=16'd15514;
      5445:data<=16'd14451;
      5446:data<=16'd13582;
      5447:data<=16'd13641;
      5448:data<=16'd13570;
      5449:data<=16'd14239;
      5450:data<=16'd13937;
      5451:data<=16'd13085;
      5452:data<=16'd12075;
      5453:data<=16'd10513;
      5454:data<=16'd10683;
      5455:data<=16'd10284;
      5456:data<=16'd9195;
      5457:data<=16'd9919;
      5458:data<=16'd9095;
      5459:data<=16'd8191;
      5460:data<=16'd8561;
      5461:data<=16'd7380;
      5462:data<=16'd7354;
      5463:data<=16'd7186;
      5464:data<=16'd6463;
      5465:data<=16'd8501;
      5466:data<=16'd7194;
      5467:data<=16'd3248;
      5468:data<=16'd2740;
      5469:data<=16'd2182;
      5470:data<=16'd2080;
      5471:data<=16'd1908;
      5472:data<=16'd640;
      5473:data<=16'd2400;
      5474:data<=-16'd2024;
      5475:data<=-16'd13505;
      5476:data<=-16'd16123;
      5477:data<=-16'd13843;
      5478:data<=-16'd14126;
      5479:data<=-16'd12668;
      5480:data<=-16'd12340;
      5481:data<=-16'd12123;
      5482:data<=-16'd9442;
      5483:data<=-16'd9063;
      5484:data<=-16'd9265;
      5485:data<=-16'd8883;
      5486:data<=-16'd9589;
      5487:data<=-16'd8590;
      5488:data<=-16'd7110;
      5489:data<=-16'd6840;
      5490:data<=-16'd6922;
      5491:data<=-16'd7642;
      5492:data<=-16'd7112;
      5493:data<=-16'd5985;
      5494:data<=-16'd5955;
      5495:data<=-16'd5624;
      5496:data<=-16'd5682;
      5497:data<=-16'd5295;
      5498:data<=-16'd3383;
      5499:data<=-16'd2102;
      5500:data<=-16'd1557;
      5501:data<=-16'd1944;
      5502:data<=-16'd2414;
      5503:data<=-16'd1577;
      5504:data<=-16'd1735;
      5505:data<=-16'd1871;
      5506:data<=-16'd1312;
      5507:data<=-16'd1915;
      5508:data<=-16'd1451;
      5509:data<=-16'd1313;
      5510:data<=-16'd1962;
      5511:data<=-16'd663;
      5512:data<=-16'd1340;
      5513:data<=-16'd1642;
      5514:data<=16'd503;
      5515:data<=-16'd488;
      5516:data<=16'd5247;
      5517:data<=16'd19367;
      5518:data<=16'd23135;
      5519:data<=16'd19767;
      5520:data<=16'd19884;
      5521:data<=16'd18483;
      5522:data<=16'd17305;
      5523:data<=16'd17643;
      5524:data<=16'd16007;
      5525:data<=16'd15540;
      5526:data<=16'd15256;
      5527:data<=16'd13955;
      5528:data<=16'd14286;
      5529:data<=16'd13459;
      5530:data<=16'd11705;
      5531:data<=16'd12157;
      5532:data<=16'd13009;
      5533:data<=16'd13066;
      5534:data<=16'd12370;
      5535:data<=16'd11361;
      5536:data<=16'd10874;
      5537:data<=16'd10149;
      5538:data<=16'd9392;
      5539:data<=16'd8857;
      5540:data<=16'd8258;
      5541:data<=16'd7944;
      5542:data<=16'd7432;
      5543:data<=16'd7043;
      5544:data<=16'd6546;
      5545:data<=16'd5624;
      5546:data<=16'd5685;
      5547:data<=16'd5513;
      5548:data<=16'd5409;
      5549:data<=16'd6725;
      5550:data<=16'd6622;
      5551:data<=16'd6150;
      5552:data<=16'd6067;
      5553:data<=16'd4388;
      5554:data<=16'd4481;
      5555:data<=16'd4584;
      5556:data<=16'd3248;
      5557:data<=16'd4457;
      5558:data<=-16'd206;
      5559:data<=-16'd11177;
      5560:data<=-16'd13879;
      5561:data<=-16'd11940;
      5562:data<=-16'd12671;
      5563:data<=-16'd12111;
      5564:data<=-16'd11432;
      5565:data<=-16'd10190;
      5566:data<=-16'd9012;
      5567:data<=-16'd12110;
      5568:data<=-16'd13937;
      5569:data<=-16'd12740;
      5570:data<=-16'd12803;
      5571:data<=-16'd12098;
      5572:data<=-16'd11317;
      5573:data<=-16'd11685;
      5574:data<=-16'd11439;
      5575:data<=-16'd11458;
      5576:data<=-16'd10957;
      5577:data<=-16'd10389;
      5578:data<=-16'd10734;
      5579:data<=-16'd9859;
      5580:data<=-16'd9318;
      5581:data<=-16'd8975;
      5582:data<=-16'd7043;
      5583:data<=-16'd6499;
      5584:data<=-16'd6614;
      5585:data<=-16'd5852;
      5586:data<=-16'd5783;
      5587:data<=-16'd5627;
      5588:data<=-16'd5756;
      5589:data<=-16'd5774;
      5590:data<=-16'd5160;
      5591:data<=-16'd5745;
      5592:data<=-16'd5419;
      5593:data<=-16'd4784;
      5594:data<=-16'd5588;
      5595:data<=-16'd4737;
      5596:data<=-16'd4632;
      5597:data<=-16'd4957;
      5598:data<=-16'd2883;
      5599:data<=-16'd2946;
      5600:data<=16'd986;
      5601:data<=16'd11820;
      5602:data<=16'd15062;
      5603:data<=16'd12442;
      5604:data<=16'd12866;
      5605:data<=16'd11699;
      5606:data<=16'd10501;
      5607:data<=16'd11080;
      5608:data<=16'd9961;
      5609:data<=16'd9508;
      5610:data<=16'd9288;
      5611:data<=16'd8493;
      5612:data<=16'd8736;
      5613:data<=16'd7746;
      5614:data<=16'd6918;
      5615:data<=16'd7579;
      5616:data<=16'd8187;
      5617:data<=16'd10658;
      5618:data<=16'd12719;
      5619:data<=16'd11755;
      5620:data<=16'd10771;
      5621:data<=16'd10128;
      5622:data<=16'd9721;
      5623:data<=16'd9453;
      5624:data<=16'd8282;
      5625:data<=16'd8078;
      5626:data<=16'd8061;
      5627:data<=16'd7089;
      5628:data<=16'd6855;
      5629:data<=16'd6216;
      5630:data<=16'd5204;
      5631:data<=16'd4949;
      5632:data<=16'd4860;
      5633:data<=16'd5098;
      5634:data<=16'd4287;
      5635:data<=16'd3265;
      5636:data<=16'd3436;
      5637:data<=16'd2702;
      5638:data<=16'd2734;
      5639:data<=16'd2563;
      5640:data<=16'd752;
      5641:data<=16'd2041;
      5642:data<=-16'd919;
      5643:data<=-16'd11913;
      5644:data<=-16'd15870;
      5645:data<=-16'd13473;
      5646:data<=-16'd13928;
      5647:data<=-16'd13139;
      5648:data<=-16'd13142;
      5649:data<=-16'd15347;
      5650:data<=-16'd14615;
      5651:data<=-16'd14041;
      5652:data<=-16'd14304;
      5653:data<=-16'd13503;
      5654:data<=-16'd13891;
      5655:data<=-16'd13521;
      5656:data<=-16'd12414;
      5657:data<=-16'd12704;
      5658:data<=-16'd12712;
      5659:data<=-16'd12689;
      5660:data<=-16'd12093;
      5661:data<=-16'd10798;
      5662:data<=-16'd11010;
      5663:data<=-16'd10778;
      5664:data<=-16'd9984;
      5665:data<=-16'd10658;
      5666:data<=-16'd11570;
      5667:data<=-16'd13286;
      5668:data<=-16'd15400;
      5669:data<=-16'd15584;
      5670:data<=-16'd14592;
      5671:data<=-16'd13787;
      5672:data<=-16'd13954;
      5673:data<=-16'd13893;
      5674:data<=-16'd12807;
      5675:data<=-16'd12581;
      5676:data<=-16'd12043;
      5677:data<=-16'd11329;
      5678:data<=-16'd11896;
      5679:data<=-16'd11298;
      5680:data<=-16'd10807;
      5681:data<=-16'd10818;
      5682:data<=-16'd10419;
      5683:data<=-16'd12504;
      5684:data<=-16'd9047;
      5685:data<=16'd2698;
      5686:data<=16'd6913;
      5687:data<=16'd4141;
      5688:data<=16'd4582;
      5689:data<=16'd4460;
      5690:data<=16'd3938;
      5691:data<=16'd4561;
      5692:data<=16'd3632;
      5693:data<=16'd3845;
      5694:data<=16'd4126;
      5695:data<=16'd2896;
      5696:data<=16'd3133;
      5697:data<=16'd3087;
      5698:data<=16'd2238;
      5699:data<=16'd1750;
      5700:data<=16'd776;
      5701:data<=16'd911;
      5702:data<=16'd1248;
      5703:data<=16'd678;
      5704:data<=16'd867;
      5705:data<=16'd737;
      5706:data<=16'd591;
      5707:data<=16'd769;
      5708:data<=16'd190;
      5709:data<=16'd490;
      5710:data<=16'd616;
      5711:data<=-16'd61;
      5712:data<=-16'd5;
      5713:data<=-16'd567;
      5714:data<=-16'd194;
      5715:data<=16'd331;
      5716:data<=-16'd1938;
      5717:data<=-16'd1494;
      5718:data<=16'd1989;
      5719:data<=16'd2717;
      5720:data<=16'd2140;
      5721:data<=16'd1933;
      5722:data<=16'd2297;
      5723:data<=16'd2211;
      5724:data<=16'd967;
      5725:data<=16'd2132;
      5726:data<=-16'd638;
      5727:data<=-16'd11030;
      5728:data<=-16'd15083;
      5729:data<=-16'd12656;
      5730:data<=-16'd13418;
      5731:data<=-16'd13188;
      5732:data<=-16'd12326;
      5733:data<=-16'd13764;
      5734:data<=-16'd13341;
      5735:data<=-16'd12605;
      5736:data<=-16'd12869;
      5737:data<=-16'd12138;
      5738:data<=-16'd11412;
      5739:data<=-16'd10611;
      5740:data<=-16'd10170;
      5741:data<=-16'd10031;
      5742:data<=-16'd9379;
      5743:data<=-16'd9711;
      5744:data<=-16'd9339;
      5745:data<=-16'd8012;
      5746:data<=-16'd8113;
      5747:data<=-16'd7480;
      5748:data<=-16'd7101;
      5749:data<=-16'd8725;
      5750:data<=-16'd8878;
      5751:data<=-16'd8011;
      5752:data<=-16'd7776;
      5753:data<=-16'd7365;
      5754:data<=-16'd7109;
      5755:data<=-16'd6601;
      5756:data<=-16'd6440;
      5757:data<=-16'd6425;
      5758:data<=-16'd5457;
      5759:data<=-16'd5419;
      5760:data<=-16'd5265;
      5761:data<=-16'd4404;
      5762:data<=-16'd4746;
      5763:data<=-16'd4067;
      5764:data<=-16'd3645;
      5765:data<=-16'd4733;
      5766:data<=-16'd4817;
      5767:data<=-16'd7221;
      5768:data<=-16'd7168;
      5769:data<=16'd2108;
      5770:data<=16'd8210;
      5771:data<=16'd6587;
      5772:data<=16'd6578;
      5773:data<=16'd6583;
      5774:data<=16'd5445;
      5775:data<=16'd6061;
      5776:data<=16'd5846;
      5777:data<=16'd5312;
      5778:data<=16'd5368;
      5779:data<=16'd4965;
      5780:data<=16'd5509;
      5781:data<=16'd5642;
      5782:data<=16'd4313;
      5783:data<=16'd3210;
      5784:data<=16'd2493;
      5785:data<=16'd2740;
      5786:data<=16'd3380;
      5787:data<=16'd3186;
      5788:data<=16'd3110;
      5789:data<=16'd2917;
      5790:data<=16'd2664;
      5791:data<=16'd2955;
      5792:data<=16'd2717;
      5793:data<=16'd2312;
      5794:data<=16'd2346;
      5795:data<=16'd2262;
      5796:data<=16'd2203;
      5797:data<=16'd2378;
      5798:data<=16'd2543;
      5799:data<=16'd1715;
      5800:data<=16'd667;
      5801:data<=16'd820;
      5802:data<=16'd584;
      5803:data<=16'd459;
      5804:data<=16'd978;
      5805:data<=16'd437;
      5806:data<=16'd1002;
      5807:data<=16'd1472;
      5808:data<=16'd346;
      5809:data<=16'd1680;
      5810:data<=-16'd814;
      5811:data<=-16'd10477;
      5812:data<=-16'd15024;
      5813:data<=-16'd13772;
      5814:data<=-16'd13459;
      5815:data<=-16'd12707;
      5816:data<=-16'd12518;
      5817:data<=-16'd11213;
      5818:data<=-16'd7087;
      5819:data<=-16'd5560;
      5820:data<=-16'd5629;
      5821:data<=-16'd4987;
      5822:data<=-16'd5368;
      5823:data<=-16'd4780;
      5824:data<=-16'd3883;
      5825:data<=-16'd3911;
      5826:data<=-16'd3500;
      5827:data<=-16'd3632;
      5828:data<=-16'd3087;
      5829:data<=-16'd2159;
      5830:data<=-16'd2578;
      5831:data<=-16'd1932;
      5832:data<=-16'd2187;
      5833:data<=-16'd4168;
      5834:data<=-16'd3673;
      5835:data<=-16'd2917;
      5836:data<=-16'd3228;
      5837:data<=-16'd2329;
      5838:data<=-16'd1689;
      5839:data<=-16'd1551;
      5840:data<=-16'd1704;
      5841:data<=-16'd1942;
      5842:data<=-16'd1233;
      5843:data<=-16'd1119;
      5844:data<=-16'd725;
      5845:data<=16'd88;
      5846:data<=-16'd620;
      5847:data<=-16'd200;
      5848:data<=16'd328;
      5849:data<=-16'd914;
      5850:data<=-16'd1293;
      5851:data<=-16'd2171;
      5852:data<=16'd50;
      5853:data<=16'd8681;
      5854:data<=16'd13511;
      5855:data<=16'd12308;
      5856:data<=16'd12120;
      5857:data<=16'd12091;
      5858:data<=16'd11350;
      5859:data<=16'd10627;
      5860:data<=16'd9938;
      5861:data<=16'd10332;
      5862:data<=16'd10056;
      5863:data<=16'd9687;
      5864:data<=16'd10319;
      5865:data<=16'd9471;
      5866:data<=16'd8185;
      5867:data<=16'd6472;
      5868:data<=16'd3462;
      5869:data<=16'd2358;
      5870:data<=16'd2314;
      5871:data<=16'd1876;
      5872:data<=16'd2264;
      5873:data<=16'd2165;
      5874:data<=16'd2187;
      5875:data<=16'd2519;
      5876:data<=16'd1797;
      5877:data<=16'd1865;
      5878:data<=16'd2096;
      5879:data<=16'd1459;
      5880:data<=16'd1627;
      5881:data<=16'd1939;
      5882:data<=16'd2021;
      5883:data<=16'd1483;
      5884:data<=16'd302;
      5885:data<=16'd499;
      5886:data<=16'd610;
      5887:data<=16'd276;
      5888:data<=16'd823;
      5889:data<=16'd493;
      5890:data<=16'd849;
      5891:data<=16'd1597;
      5892:data<=16'd637;
      5893:data<=16'd1410;
      5894:data<=-16'd394;
      5895:data<=-16'd8640;
      5896:data<=-16'd13235;
      5897:data<=-16'd11938;
      5898:data<=-16'd10956;
      5899:data<=-16'd10314;
      5900:data<=-16'd10053;
      5901:data<=-16'd9683;
      5902:data<=-16'd8531;
      5903:data<=-16'd8258;
      5904:data<=-16'd7730;
      5905:data<=-16'd7178;
      5906:data<=-16'd7359;
      5907:data<=-16'd6579;
      5908:data<=-16'd5903;
      5909:data<=-16'd5328;
      5910:data<=-16'd4642;
      5911:data<=-16'd5322;
      5912:data<=-16'd5036;
      5913:data<=-16'd3996;
      5914:data<=-16'd3983;
      5915:data<=-16'd2940;
      5916:data<=-16'd1944;
      5917:data<=-16'd751;
      5918:data<=16'd2409;
      5919:data<=16'd4049;
      5920:data<=16'd4350;
      5921:data<=16'd5207;
      5922:data<=16'd4927;
      5923:data<=16'd4760;
      5924:data<=16'd4837;
      5925:data<=16'd4367;
      5926:data<=16'd4904;
      5927:data<=16'd5074;
      5928:data<=16'd4805;
      5929:data<=16'd5181;
      5930:data<=16'd4822;
      5931:data<=16'd4822;
      5932:data<=16'd5266;
      5933:data<=16'd5847;
      5934:data<=16'd7456;
      5935:data<=16'd6772;
      5936:data<=16'd6865;
      5937:data<=16'd13832;
      5938:data<=16'd19936;
      5939:data<=16'd19707;
      5940:data<=16'd18747;
      5941:data<=16'd18215;
      5942:data<=16'd17286;
      5943:data<=16'd17149;
      5944:data<=16'd16631;
      5945:data<=16'd15676;
      5946:data<=16'd15365;
      5947:data<=16'd15059;
      5948:data<=16'd14413;
      5949:data<=16'd14530;
      5950:data<=16'd15380;
      5951:data<=16'd15080;
      5952:data<=16'd14220;
      5953:data<=16'd14117;
      5954:data<=16'd13502;
      5955:data<=16'd12701;
      5956:data<=16'd12339;
      5957:data<=16'd11923;
      5958:data<=16'd11885;
      5959:data<=16'd11221;
      5960:data<=16'd10527;
      5961:data<=16'd10686;
      5962:data<=16'd9395;
      5963:data<=16'd8778;
      5964:data<=16'd9697;
      5965:data<=16'd8602;
      5966:data<=16'd8768;
      5967:data<=16'd10017;
      5968:data<=16'd7354;
      5969:data<=16'd5151;
      5970:data<=16'd5037;
      5971:data<=16'd3833;
      5972:data<=16'd3680;
      5973:data<=16'd3929;
      5974:data<=16'd3891;
      5975:data<=16'd4402;
      5976:data<=16'd3213;
      5977:data<=16'd3210;
      5978:data<=16'd3207;
      5979:data<=-16'd3480;
      5980:data<=-16'd10107;
      5981:data<=-16'd10593;
      5982:data<=-16'd9850;
      5983:data<=-16'd8548;
      5984:data<=-16'd7180;
      5985:data<=-16'd7363;
      5986:data<=-16'd6669;
      5987:data<=-16'd5971;
      5988:data<=-16'd6147;
      5989:data<=-16'd5820;
      5990:data<=-16'd5955;
      5991:data<=-16'd5956;
      5992:data<=-16'd5338;
      5993:data<=-16'd5021;
      5994:data<=-16'd4681;
      5995:data<=-16'd4968;
      5996:data<=-16'd4945;
      5997:data<=-16'd3811;
      5998:data<=-16'd3662;
      5999:data<=-16'd3206;
      6000:data<=-16'd1571;
      6001:data<=-16'd1130;
      6002:data<=-16'd1113;
      6003:data<=-16'd694;
      6004:data<=-16'd579;
      6005:data<=-16'd640;
      6006:data<=-16'd914;
      6007:data<=-16'd472;
      6008:data<=16'd97;
      6009:data<=-16'd497;
      6010:data<=-16'd758;
      6011:data<=-16'd901;
      6012:data<=-16'd1099;
      6013:data<=-16'd331;
      6014:data<=-16'd237;
      6015:data<=-16'd308;
      6016:data<=16'd247;
      6017:data<=16'd837;
      6018:data<=16'd3770;
      6019:data<=16'd6119;
      6020:data<=16'd5967;
      6021:data<=16'd11157;
      6022:data<=16'd18879;
      6023:data<=16'd19409;
      6024:data<=16'd17394;
      6025:data<=16'd17388;
      6026:data<=16'd16324;
      6027:data<=16'd15479;
      6028:data<=16'd15496;
      6029:data<=16'd14600;
      6030:data<=16'd14055;
      6031:data<=16'd13755;
      6032:data<=16'd12977;
      6033:data<=16'd13164;
      6034:data<=16'd13577;
      6035:data<=16'd13109;
      6036:data<=16'd13022;
      6037:data<=16'd12816;
      6038:data<=16'd11486;
      6039:data<=16'd10701;
      6040:data<=16'd10907;
      6041:data<=16'd10769;
      6042:data<=16'd10141;
      6043:data<=16'd9318;
      6044:data<=16'd8701;
      6045:data<=16'd8275;
      6046:data<=16'd7583;
      6047:data<=16'd7139;
      6048:data<=16'd6543;
      6049:data<=16'd5920;
      6050:data<=16'd6755;
      6051:data<=16'd7043;
      6052:data<=16'd6059;
      6053:data<=16'd6388;
      6054:data<=16'd6252;
      6055:data<=16'd5156;
      6056:data<=16'd5318;
      6057:data<=16'd4513;
      6058:data<=16'd3765;
      6059:data<=16'd4683;
      6060:data<=16'd3359;
      6061:data<=16'd2749;
      6062:data<=16'd3974;
      6063:data<=-16'd1519;
      6064:data<=-16'd9994;
      6065:data<=-16'd11705;
      6066:data<=-16'd9629;
      6067:data<=-16'd8019;
      6068:data<=-16'd8584;
      6069:data<=-16'd11565;
      6070:data<=-16'd12254;
      6071:data<=-16'd11421;
      6072:data<=-16'd11990;
      6073:data<=-16'd11332;
      6074:data<=-16'd10707;
      6075:data<=-16'd11082;
      6076:data<=-16'd10016;
      6077:data<=-16'd9545;
      6078:data<=-16'd9832;
      6079:data<=-16'd9168;
      6080:data<=-16'd9086;
      6081:data<=-16'd9227;
      6082:data<=-16'd9259;
      6083:data<=-16'd8573;
      6084:data<=-16'd6106;
      6085:data<=-16'd5527;
      6086:data<=-16'd6655;
      6087:data<=-16'd5876;
      6088:data<=-16'd5392;
      6089:data<=-16'd5492;
      6090:data<=-16'd4822;
      6091:data<=-16'd4999;
      6092:data<=-16'd5139;
      6093:data<=-16'd4851;
      6094:data<=-16'd4949;
      6095:data<=-16'd4625;
      6096:data<=-16'd4381;
      6097:data<=-16'd4404;
      6098:data<=-16'd4447;
      6099:data<=-16'd3971;
      6100:data<=-16'd2532;
      6101:data<=-16'd2218;
      6102:data<=-16'd1736;
      6103:data<=-16'd955;
      6104:data<=-16'd2599;
      6105:data<=16'd926;
      6106:data<=16'd10348;
      6107:data<=16'd12558;
      6108:data<=16'd9871;
      6109:data<=16'd10323;
      6110:data<=16'd9929;
      6111:data<=16'd8523;
      6112:data<=16'd8581;
      6113:data<=16'd8420;
      6114:data<=16'd7605;
      6115:data<=16'd6737;
      6116:data<=16'd7260;
      6117:data<=16'd8372;
      6118:data<=16'd8945;
      6119:data<=16'd10925;
      6120:data<=16'd12129;
      6121:data<=16'd11068;
      6122:data<=16'd10555;
      6123:data<=16'd9950;
      6124:data<=16'd9066;
      6125:data<=16'd8402;
      6126:data<=16'd7429;
      6127:data<=16'd7582;
      6128:data<=16'd7257;
      6129:data<=16'd5943;
      6130:data<=16'd5811;
      6131:data<=16'd5072;
      6132:data<=16'd4563;
      6133:data<=16'd5500;
      6134:data<=16'd5542;
      6135:data<=16'd5497;
      6136:data<=16'd5274;
      6137:data<=16'd4936;
      6138:data<=16'd5309;
      6139:data<=16'd4049;
      6140:data<=16'd3560;
      6141:data<=16'd4206;
      6142:data<=16'd2716;
      6143:data<=16'd2675;
      6144:data<=16'd2275;
      6145:data<=16'd570;
      6146:data<=16'd2660;
      6147:data<=-16'd638;
      6148:data<=-16'd10950;
      6149:data<=-16'd13729;
      6150:data<=-16'd11374;
      6151:data<=-16'd10948;
      6152:data<=-16'd10028;
      6153:data<=-16'd10008;
      6154:data<=-16'd10287;
      6155:data<=-16'd9514;
      6156:data<=-16'd9286;
      6157:data<=-16'd8513;
      6158:data<=-16'd8499;
      6159:data<=-16'd9649;
      6160:data<=-16'd9317;
      6161:data<=-16'd8624;
      6162:data<=-16'd8598;
      6163:data<=-16'd8742;
      6164:data<=-16'd8539;
      6165:data<=-16'd8160;
      6166:data<=-16'd8627;
      6167:data<=-16'd8175;
      6168:data<=-16'd8408;
      6169:data<=-16'd11508;
      6170:data<=-16'd12317;
      6171:data<=-16'd11248;
      6172:data<=-16'd11662;
      6173:data<=-16'd11032;
      6174:data<=-16'd10536;
      6175:data<=-16'd10566;
      6176:data<=-16'd9649;
      6177:data<=-16'd9955;
      6178:data<=-16'd10014;
      6179:data<=-16'd9629;
      6180:data<=-16'd10097;
      6181:data<=-16'd9132;
      6182:data<=-16'd8965;
      6183:data<=-16'd9940;
      6184:data<=-16'd9987;
      6185:data<=-16'd11100;
      6186:data<=-16'd10161;
      6187:data<=-16'd8725;
      6188:data<=-16'd11113;
      6189:data<=-16'd7236;
      6190:data<=16'd2500;
      6191:data<=16'd4672;
      6192:data<=16'd3055;
      6193:data<=16'd3979;
      6194:data<=16'd3627;
      6195:data<=16'd2822;
      6196:data<=16'd3060;
      6197:data<=16'd2479;
      6198:data<=16'd1924;
      6199:data<=16'd2273;
      6200:data<=16'd1952;
      6201:data<=16'd537;
      6202:data<=-16'd306;
      6203:data<=-16'd414;
      6204:data<=-16'd387;
      6205:data<=-16'd111;
      6206:data<=-16'd526;
      6207:data<=-16'd1024;
      6208:data<=-16'd872;
      6209:data<=-16'd1192;
      6210:data<=-16'd1163;
      6211:data<=-16'd1143;
      6212:data<=-16'd1544;
      6213:data<=-16'd863;
      6214:data<=-16'd1428;
      6215:data<=-16'd2620;
      6216:data<=-16'd2032;
      6217:data<=-16'd3206;
      6218:data<=-16'd3488;
      6219:data<=-16'd6;
      6220:data<=16'd834;
      6221:data<=16'd26;
      6222:data<=16'd526;
      6223:data<=-16'd491;
      6224:data<=-16'd523;
      6225:data<=-16'd38;
      6226:data<=-16'd1213;
      6227:data<=-16'd423;
      6228:data<=-16'd546;
      6229:data<=-16'd1811;
      6230:data<=16'd114;
      6231:data<=-16'd3193;
      6232:data<=-16'd12336;
      6233:data<=-16'd15083;
      6234:data<=-16'd14324;
      6235:data<=-16'd15593;
      6236:data<=-16'd14898;
      6237:data<=-16'd13806;
      6238:data<=-16'd13711;
      6239:data<=-16'd12784;
      6240:data<=-16'd12806;
      6241:data<=-16'd12660;
      6242:data<=-16'd11491;
      6243:data<=-16'd11664;
      6244:data<=-16'd11530;
      6245:data<=-16'd10483;
      6246:data<=-16'd10281;
      6247:data<=-16'd9720;
      6248:data<=-16'd9010;
      6249:data<=-16'd9283;
      6250:data<=-16'd9761;
      6251:data<=-16'd10329;
      6252:data<=-16'd10425;
      6253:data<=-16'd9831;
      6254:data<=-16'd9741;
      6255:data<=-16'd9635;
      6256:data<=-16'd8733;
      6257:data<=-16'd8103;
      6258:data<=-16'd8055;
      6259:data<=-16'd7589;
      6260:data<=-16'd7122;
      6261:data<=-16'd7448;
      6262:data<=-16'd7436;
      6263:data<=-16'd6957;
      6264:data<=-16'd6420;
      6265:data<=-16'd5327;
      6266:data<=-16'd4939;
      6267:data<=-16'd5083;
      6268:data<=-16'd6240;
      6269:data<=-16'd10249;
      6270:data<=-16'd11359;
      6271:data<=-16'd9350;
      6272:data<=-16'd10733;
      6273:data<=-16'd7087;
      6274:data<=16'd2940;
      6275:data<=16'd5213;
      6276:data<=16'd3636;
      6277:data<=16'd5080;
      6278:data<=16'd3973;
      6279:data<=16'd3334;
      6280:data<=16'd4734;
      6281:data<=16'd4041;
      6282:data<=16'd3899;
      6283:data<=16'd3662;
      6284:data<=16'd1898;
      6285:data<=16'd1548;
      6286:data<=16'd1569;
      6287:data<=16'd1245;
      6288:data<=16'd1125;
      6289:data<=16'd955;
      6290:data<=16'd1600;
      6291:data<=16'd1539;
      6292:data<=16'd934;
      6293:data<=16'd1504;
      6294:data<=16'd1500;
      6295:data<=16'd1433;
      6296:data<=16'd2097;
      6297:data<=16'd1841;
      6298:data<=16'd1381;
      6299:data<=16'd1334;
      6300:data<=16'd1055;
      6301:data<=-16'd3;
      6302:data<=-16'd1181;
      6303:data<=-16'd817;
      6304:data<=-16'd473;
      6305:data<=-16'd690;
      6306:data<=-16'd469;
      6307:data<=-16'd974;
      6308:data<=-16'd597;
      6309:data<=16'd20;
      6310:data<=-16'd613;
      6311:data<=16'd594;
      6312:data<=16'd375;
      6313:data<=-16'd887;
      6314:data<=16'd1782;
      6315:data<=-16'd1227;
      6316:data<=-16'd10875;
      6317:data<=-16'd14458;
      6318:data<=-16'd13591;
      6319:data<=-16'd11623;
      6320:data<=-16'd8387;
      6321:data<=-16'd8235;
      6322:data<=-16'd8310;
      6323:data<=-16'd7030;
      6324:data<=-16'd7172;
      6325:data<=-16'd6445;
      6326:data<=-16'd5821;
      6327:data<=-16'd5906;
      6328:data<=-16'd4930;
      6329:data<=-16'd4802;
      6330:data<=-16'd4564;
      6331:data<=-16'd4070;
      6332:data<=-16'd4249;
      6333:data<=-16'd3339;
      6334:data<=-16'd3899;
      6335:data<=-16'd5312;
      6336:data<=-16'd4557;
      6337:data<=-16'd4535;
      6338:data<=-16'd4411;
      6339:data<=-16'd3503;
      6340:data<=-16'd3918;
      6341:data<=-16'd3465;
      6342:data<=-16'd2978;
      6343:data<=-16'd2720;
      6344:data<=-16'd1118;
      6345:data<=-16'd1306;
      6346:data<=-16'd1841;
      6347:data<=-16'd1204;
      6348:data<=-16'd1366;
      6349:data<=-16'd384;
      6350:data<=-16'd487;
      6351:data<=-16'd2146;
      6352:data<=-16'd1553;
      6353:data<=-16'd2088;
      6354:data<=-16'd2482;
      6355:data<=-16'd1183;
      6356:data<=-16'd2511;
      6357:data<=16'd1192;
      6358:data<=16'd10915;
      6359:data<=16'd13626;
      6360:data<=16'd11967;
      6361:data<=16'd12569;
      6362:data<=16'd12198;
      6363:data<=16'd11512;
      6364:data<=16'd11292;
      6365:data<=16'd10812;
      6366:data<=16'd11022;
      6367:data<=16'd10299;
      6368:data<=16'd8392;
      6369:data<=16'd6191;
      6370:data<=16'd3676;
      6371:data<=16'd2704;
      6372:data<=16'd3230;
      6373:data<=16'd3412;
      6374:data<=16'd3240;
      6375:data<=16'd3281;
      6376:data<=16'd3597;
      6377:data<=16'd3372;
      6378:data<=16'd2902;
      6379:data<=16'd3106;
      6380:data<=16'd3321;
      6381:data<=16'd3647;
      6382:data<=16'd3859;
      6383:data<=16'd3425;
      6384:data<=16'd3052;
      6385:data<=16'd2018;
      6386:data<=16'd1316;
      6387:data<=16'd2030;
      6388:data<=16'd1582;
      6389:data<=16'd1222;
      6390:data<=16'd2052;
      6391:data<=16'd1516;
      6392:data<=16'd1475;
      6393:data<=16'd1745;
      6394:data<=16'd1011;
      6395:data<=16'd2475;
      6396:data<=16'd2889;
      6397:data<=16'd1416;
      6398:data<=16'd3171;
      6399:data<=16'd811;
      6400:data<=-16'd8298;
      6401:data<=-16'd12343;
      6402:data<=-16'd11655;
      6403:data<=-16'd12031;
      6404:data<=-16'd10894;
      6405:data<=-16'd9480;
      6406:data<=-16'd9448;
      6407:data<=-16'd8831;
      6408:data<=-16'd8570;
      6409:data<=-16'd8288;
      6410:data<=-16'd6930;
      6411:data<=-16'd6232;
      6412:data<=-16'd6263;
      6413:data<=-16'd5976;
      6414:data<=-16'd5548;
      6415:data<=-16'd4946;
      6416:data<=-16'd3997;
      6417:data<=-16'd4121;
      6418:data<=-16'd5673;
      6419:data<=-16'd4405;
      6420:data<=-16'd288;
      6421:data<=16'd716;
      6422:data<=-16'd240;
      6423:data<=16'd255;
      6424:data<=16'd411;
      6425:data<=16'd694;
      6426:data<=16'd1391;
      6427:data<=16'd1510;
      6428:data<=16'd2190;
      6429:data<=16'd2335;
      6430:data<=16'd1905;
      6431:data<=16'd2155;
      6432:data<=16'd2067;
      6433:data<=16'd2629;
      6434:data<=16'd3269;
      6435:data<=16'd3039;
      6436:data<=16'd3657;
      6437:data<=16'd3010;
      6438:data<=16'd2549;
      6439:data<=16'd4196;
      6440:data<=16'd3027;
      6441:data<=16'd5013;
      6442:data<=16'd14205;
      6443:data<=16'd17892;
      6444:data<=16'd15940;
      6445:data<=16'd16261;
      6446:data<=16'd15497;
      6447:data<=16'd14498;
      6448:data<=16'd15283;
      6449:data<=16'd14449;
      6450:data<=16'd13526;
      6451:data<=16'd14046;
      6452:data<=16'd14675;
      6453:data<=16'd14953;
      6454:data<=16'd14304;
      6455:data<=16'd13694;
      6456:data<=16'd13567;
      6457:data<=16'd13361;
      6458:data<=16'd13189;
      6459:data<=16'd12636;
      6460:data<=16'd12319;
      6461:data<=16'd11966;
      6462:data<=16'd11242;
      6463:data<=16'd11411;
      6464:data<=16'd10868;
      6465:data<=16'd9831;
      6466:data<=16'd9864;
      6467:data<=16'd9673;
      6468:data<=16'd10730;
      6469:data<=16'd10690;
      6470:data<=16'd6649;
      6471:data<=16'd5251;
      6472:data<=16'd6529;
      6473:data<=16'd6043;
      6474:data<=16'd6287;
      6475:data<=16'd5920;
      6476:data<=16'd4871;
      6477:data<=16'd5409;
      6478:data<=16'd5037;
      6479:data<=16'd5212;
      6480:data<=16'd5163;
      6481:data<=16'd3786;
      6482:data<=16'd5692;
      6483:data<=16'd3712;
      6484:data<=-16'd5059;
      6485:data<=-16'd7727;
      6486:data<=-16'd5879;
      6487:data<=-16'd6425;
      6488:data<=-16'd5732;
      6489:data<=-16'd5195;
      6490:data<=-16'd5635;
      6491:data<=-16'd4713;
      6492:data<=-16'd4548;
      6493:data<=-16'd4616;
      6494:data<=-16'd4003;
      6495:data<=-16'd3838;
      6496:data<=-16'd3471;
      6497:data<=-16'd3198;
      6498:data<=-16'd2957;
      6499:data<=-16'd2837;
      6500:data<=-16'd3290;
      6501:data<=-16'd2435;
      6502:data<=-16'd873;
      6503:data<=-16'd258;
      6504:data<=16'd250;
      6505:data<=16'd1008;
      6506:data<=16'd2397;
      6507:data<=16'd3268;
      6508:data<=16'd2581;
      6509:data<=16'd2272;
      6510:data<=16'd2191;
      6511:data<=16'd2006;
      6512:data<=16'd2358;
      6513:data<=16'd2012;
      6514:data<=16'd1718;
      6515:data<=16'd1601;
      6516:data<=16'd1048;
      6517:data<=16'd1712;
      6518:data<=16'd2504;
      6519:data<=16'd3903;
      6520:data<=16'd6429;
      6521:data<=16'd5738;
      6522:data<=16'd4817;
      6523:data<=16'd6011;
      6524:data<=16'd4309;
      6525:data<=16'd6108;
      6526:data<=16'd14797;
      6527:data<=16'd18534;
      6528:data<=16'd16873;
      6529:data<=16'd16728;
      6530:data<=16'd15914;
      6531:data<=16'd14647;
      6532:data<=16'd14681;
      6533:data<=16'd14013;
      6534:data<=16'd13797;
      6535:data<=16'd14687;
      6536:data<=16'd14249;
      6537:data<=16'd13010;
      6538:data<=16'd12630;
      6539:data<=16'd12395;
      6540:data<=16'd11721;
      6541:data<=16'd11171;
      6542:data<=16'd10892;
      6543:data<=16'd10601;
      6544:data<=16'd10055;
      6545:data<=16'd9180;
      6546:data<=16'd8419;
      6547:data<=16'd7949;
      6548:data<=16'd7627;
      6549:data<=16'd7304;
      6550:data<=16'd6617;
      6551:data<=16'd6531;
      6552:data<=16'd7442;
      6553:data<=16'd7430;
      6554:data<=16'd6896;
      6555:data<=16'd7071;
      6556:data<=16'd6546;
      6557:data<=16'd5858;
      6558:data<=16'd6068;
      6559:data<=16'd5849;
      6560:data<=16'd5184;
      6561:data<=16'd4397;
      6562:data<=16'd3926;
      6563:data<=16'd4501;
      6564:data<=16'd3891;
      6565:data<=16'd2896;
      6566:data<=16'd4190;
      6567:data<=16'd2244;
      6568:data<=-16'd4972;
      6569:data<=-16'd9482;
      6570:data<=-16'd10038;
      6571:data<=-16'd10404;
      6572:data<=-16'd9674;
      6573:data<=-16'd8871;
      6574:data<=-16'd9268;
      6575:data<=-16'd8872;
      6576:data<=-16'd8448;
      6577:data<=-16'd8768;
      6578:data<=-16'd8411;
      6579:data<=-16'd8111;
      6580:data<=-16'd8117;
      6581:data<=-16'd7538;
      6582:data<=-16'd7444;
      6583:data<=-16'd7923;
      6584:data<=-16'd7245;
      6585:data<=-16'd5706;
      6586:data<=-16'd4911;
      6587:data<=-16'd4525;
      6588:data<=-16'd4027;
      6589:data<=-16'd4326;
      6590:data<=-16'd4696;
      6591:data<=-16'd4202;
      6592:data<=-16'd4081;
      6593:data<=-16'd4279;
      6594:data<=-16'd4129;
      6595:data<=-16'd4035;
      6596:data<=-16'd3761;
      6597:data<=-16'd3847;
      6598:data<=-16'd4328;
      6599:data<=-16'd4175;
      6600:data<=-16'd4014;
      6601:data<=-16'd3192;
      6602:data<=-16'd1348;
      6603:data<=-16'd829;
      6604:data<=-16'd1310;
      6605:data<=-16'd1779;
      6606:data<=-16'd2036;
      6607:data<=-16'd1313;
      6608:data<=-16'd1868;
      6609:data<=-16'd1287;
      6610:data<=16'd5594;
      6611:data<=16'd11489;
      6612:data<=16'd10769;
      6613:data<=16'd9611;
      6614:data<=16'd9279;
      6615:data<=16'd8296;
      6616:data<=16'd8247;
      6617:data<=16'd7776;
      6618:data<=16'd7565;
      6619:data<=16'd9045;
      6620:data<=16'd9818;
      6621:data<=16'd9847;
      6622:data<=16'd9568;
      6623:data<=16'd8393;
      6624:data<=16'd7987;
      6625:data<=16'd8032;
      6626:data<=16'd7309;
      6627:data<=16'd6789;
      6628:data<=16'd6449;
      6629:data<=16'd5897;
      6630:data<=16'd5341;
      6631:data<=16'd4942;
      6632:data<=16'd4601;
      6633:data<=16'd3738;
      6634:data<=16'd3691;
      6635:data<=16'd5031;
      6636:data<=16'd5218;
      6637:data<=16'd4353;
      6638:data<=16'd4064;
      6639:data<=16'd3923;
      6640:data<=16'd3821;
      6641:data<=16'd3389;
      6642:data<=16'd2681;
      6643:data<=16'd2505;
      6644:data<=16'd2203;
      6645:data<=16'd1741;
      6646:data<=16'd1245;
      6647:data<=16'd676;
      6648:data<=16'd839;
      6649:data<=16'd638;
      6650:data<=16'd459;
      6651:data<=16'd82;
      6652:data<=-16'd5301;
      6653:data<=-16'd11952;
      6654:data<=-16'd12292;
      6655:data<=-16'd10887;
      6656:data<=-16'd11248;
      6657:data<=-16'd10678;
      6658:data<=-16'd10343;
      6659:data<=-16'd10169;
      6660:data<=-16'd9571;
      6661:data<=-16'd10107;
      6662:data<=-16'd10061;
      6663:data<=-16'd9236;
      6664:data<=-16'd9189;
      6665:data<=-16'd8739;
      6666:data<=-16'd8598;
      6667:data<=-16'd9268;
      6668:data<=-16'd8530;
      6669:data<=-16'd7347;
      6670:data<=-16'd8158;
      6671:data<=-16'd9538;
      6672:data<=-16'd9165;
      6673:data<=-16'd8191;
      6674:data<=-16'd8011;
      6675:data<=-16'd7735;
      6676:data<=-16'd7706;
      6677:data<=-16'd8103;
      6678:data<=-16'd7917;
      6679:data<=-16'd7835;
      6680:data<=-16'd7867;
      6681:data<=-16'd7756;
      6682:data<=-16'd7858;
      6683:data<=-16'd7344;
      6684:data<=-16'd7119;
      6685:data<=-16'd6924;
      6686:data<=-16'd5385;
      6687:data<=-16'd5010;
      6688:data<=-16'd5098;
      6689:data<=-16'd4449;
      6690:data<=-16'd5579;
      6691:data<=-16'd5647;
      6692:data<=-16'd4751;
      6693:data<=-16'd4895;
      6694:data<=16'd958;
      6695:data<=16'd8951;
      6696:data<=16'd8774;
      6697:data<=16'd6934;
      6698:data<=16'd7692;
      6699:data<=16'd6661;
      6700:data<=16'd5620;
      6701:data<=16'd5093;
      6702:data<=16'd4457;
      6703:data<=16'd5025;
      6704:data<=16'd4673;
      6705:data<=16'd3761;
      6706:data<=16'd3664;
      6707:data<=16'd2946;
      6708:data<=16'd2708;
      6709:data<=16'd2883;
      6710:data<=16'd2350;
      6711:data<=16'd2678;
      6712:data<=16'd2981;
      6713:data<=16'd2118;
      6714:data<=16'd1560;
      6715:data<=16'd1268;
      6716:data<=16'd1019;
      6717:data<=16'd1024;
      6718:data<=16'd106;
      6719:data<=-16'd1453;
      6720:data<=-16'd1337;
      6721:data<=16'd240;
      6722:data<=16'd557;
      6723:data<=-16'd299;
      6724:data<=-16'd778;
      6725:data<=-16'd1010;
      6726:data<=-16'd705;
      6727:data<=-16'd604;
      6728:data<=-16'd1143;
      6729:data<=-16'd723;
      6730:data<=-16'd808;
      6731:data<=-16'd1598;
      6732:data<=-16'd1092;
      6733:data<=-16'd1666;
      6734:data<=-16'd1979;
      6735:data<=-16'd1381;
      6736:data<=-16'd7696;
      6737:data<=-16'd16806;
      6738:data<=-16'd17841;
      6739:data<=-16'd15995;
      6740:data<=-16'd16490;
      6741:data<=-16'd15882;
      6742:data<=-16'd14871;
      6743:data<=-16'd14410;
      6744:data<=-16'd13828;
      6745:data<=-16'd13574;
      6746:data<=-16'd12822;
      6747:data<=-16'd12349;
      6748:data<=-16'd12502;
      6749:data<=-16'd11841;
      6750:data<=-16'd11462;
      6751:data<=-16'd11635;
      6752:data<=-16'd12028;
      6753:data<=-16'd13176;
      6754:data<=-16'd13088;
      6755:data<=-16'd12098;
      6756:data<=-16'd12182;
      6757:data<=-16'd11715;
      6758:data<=-16'd10971;
      6759:data<=-16'd10989;
      6760:data<=-16'd10211;
      6761:data<=-16'd9523;
      6762:data<=-16'd9838;
      6763:data<=-16'd9433;
      6764:data<=-16'd8393;
      6765:data<=-16'd8129;
      6766:data<=-16'd8178;
      6767:data<=-16'd7565;
      6768:data<=-16'd7656;
      6769:data<=-16'd9036;
      6770:data<=-16'd10032;
      6771:data<=-16'd11009;
      6772:data<=-16'd11142;
      6773:data<=-16'd9579;
      6774:data<=-16'd9530;
      6775:data<=-16'd9621;
      6776:data<=-16'd8866;
      6777:data<=-16'd9700;
      6778:data<=-16'd5045;
      6779:data<=16'd4625;
      6780:data<=16'd6593;
      6781:data<=16'd4552;
      6782:data<=16'd5802;
      6783:data<=16'd5856;
      6784:data<=16'd5247;
      6785:data<=16'd4631;
      6786:data<=16'd2349;
      6787:data<=16'd1592;
      6788:data<=16'd1800;
      6789:data<=16'd1861;
      6790:data<=16'd2376;
      6791:data<=16'd1700;
      6792:data<=16'd1638;
      6793:data<=16'd2120;
      6794:data<=16'd1541;
      6795:data<=16'd2247;
      6796:data<=16'd2396;
      6797:data<=16'd1692;
      6798:data<=16'd2736;
      6799:data<=16'd2347;
      6800:data<=16'd1536;
      6801:data<=16'd2613;
      6802:data<=16'd1891;
      6803:data<=16'd344;
      6804:data<=16'd121;
      6805:data<=16'd45;
      6806:data<=16'd185;
      6807:data<=16'd58;
      6808:data<=16'd230;
      6809:data<=16'd763;
      6810:data<=16'd362;
      6811:data<=16'd274;
      6812:data<=16'd490;
      6813:data<=16'd890;
      6814:data<=16'd1369;
      6815:data<=16'd455;
      6816:data<=16'd614;
      6817:data<=16'd1254;
      6818:data<=16'd456;
      6819:data<=16'd614;
      6820:data<=-16'd3518;
      6821:data<=-16'd11515;
      6822:data<=-16'd12454;
      6823:data<=-16'd10477;
      6824:data<=-16'd11295;
      6825:data<=-16'd10064;
      6826:data<=-16'd8681;
      6827:data<=-16'd8645;
      6828:data<=-16'd7894;
      6829:data<=-16'd7589;
      6830:data<=-16'd6852;
      6831:data<=-16'd6367;
      6832:data<=-16'd6704;
      6833:data<=-16'd5794;
      6834:data<=-16'd5195;
      6835:data<=-16'd5468;
      6836:data<=-16'd6346;
      6837:data<=-16'd7783;
      6838:data<=-16'd7292;
      6839:data<=-16'd6563;
      6840:data<=-16'd6666;
      6841:data<=-16'd5717;
      6842:data<=-16'd5462;
      6843:data<=-16'd5204;
      6844:data<=-16'd4405;
      6845:data<=-16'd4587;
      6846:data<=-16'd3753;
      6847:data<=-16'd3104;
      6848:data<=-16'd3350;
      6849:data<=-16'd2654;
      6850:data<=-16'd2728;
      6851:data<=-16'd2188;
      6852:data<=-16'd1876;
      6853:data<=-16'd4111;
      6854:data<=-16'd3953;
      6855:data<=-16'd2966;
      6856:data<=-16'd3507;
      6857:data<=-16'd2194;
      6858:data<=-16'd2584;
      6859:data<=-16'd2907;
      6860:data<=-16'd980;
      6861:data<=-16'd2199;
      6862:data<=16'd1688;
      6863:data<=16'd11897;
      6864:data<=16'd13802;
      6865:data<=16'd11468;
      6866:data<=16'd12395;
      6867:data<=16'd11985;
      6868:data<=16'd11449;
      6869:data<=16'd11027;
      6870:data<=16'd8608;
      6871:data<=16'd6613;
      6872:data<=16'd5803;
      6873:data<=16'd6351;
      6874:data<=16'd6816;
      6875:data<=16'd5914;
      6876:data<=16'd5965;
      6877:data<=16'd5988;
      6878:data<=16'd5506;
      6879:data<=16'd6200;
      6880:data<=16'd6526;
      6881:data<=16'd6587;
      6882:data<=16'd6575;
      6883:data<=16'd6043;
      6884:data<=16'd6510;
      6885:data<=16'd6167;
      6886:data<=16'd4491;
      6887:data<=16'd3896;
      6888:data<=16'd3806;
      6889:data<=16'd4205;
      6890:data<=16'd4355;
      6891:data<=16'd3512;
      6892:data<=16'd3773;
      6893:data<=16'd4021;
      6894:data<=16'd3993;
      6895:data<=16'd4614;
      6896:data<=16'd3720;
      6897:data<=16'd3512;
      6898:data<=16'd4443;
      6899:data<=16'd3662;
      6900:data<=16'd4182;
      6901:data<=16'd4434;
      6902:data<=16'd2719;
      6903:data<=16'd3224;
      6904:data<=-16'd503;
      6905:data<=-16'd9749;
      6906:data<=-16'd11979;
      6907:data<=-16'd9574;
      6908:data<=-16'd10076;
      6909:data<=-16'd9485;
      6910:data<=-16'd8258;
      6911:data<=-16'd8197;
      6912:data<=-16'd7092;
      6913:data<=-16'd6510;
      6914:data<=-16'd6419;
      6915:data<=-16'd5827;
      6916:data<=-16'd5909;
      6917:data<=-16'd5002;
      6918:data<=-16'd3809;
      6919:data<=-16'd4843;
      6920:data<=-16'd5457;
      6921:data<=-16'd4202;
      6922:data<=-16'd3055;
      6923:data<=-16'd2393;
      6924:data<=-16'd2056;
      6925:data<=-16'd2099;
      6926:data<=-16'd2176;
      6927:data<=-16'd2076;
      6928:data<=-16'd1583;
      6929:data<=-16'd939;
      6930:data<=-16'd649;
      6931:data<=-16'd528;
      6932:data<=-16'd102;
      6933:data<=16'd167;
      6934:data<=16'd161;
      6935:data<=16'd522;
      6936:data<=-16'd96;
      6937:data<=-16'd1516;
      6938:data<=-16'd1254;
      6939:data<=-16'd826;
      6940:data<=-16'd596;
      6941:data<=16'd561;
      6942:data<=-16'd45;
      6943:data<=-16'd62;
      6944:data<=16'd1133;
      6945:data<=-16'd722;
      6946:data<=16'd3028;
      6947:data<=16'd13732;
      6948:data<=16'd15931;
      6949:data<=16'd12706;
      6950:data<=16'd13869;
      6951:data<=16'd13937;
      6952:data<=16'd12269;
      6953:data<=16'd11274;
      6954:data<=16'd9627;
      6955:data<=16'd9276;
      6956:data<=16'd9294;
      6957:data<=16'd9153;
      6958:data<=16'd9688;
      6959:data<=16'd8589;
      6960:data<=16'd8132;
      6961:data<=16'd8907;
      6962:data<=16'd8166;
      6963:data<=16'd8501;
      6964:data<=16'd9010;
      6965:data<=16'd7943;
      6966:data<=16'd7970;
      6967:data<=16'd7697;
      6968:data<=16'd7230;
      6969:data<=16'd8109;
      6970:data<=16'd7536;
      6971:data<=16'd5968;
      6972:data<=16'd5322;
      6973:data<=16'd5046;
      6974:data<=16'd4858;
      6975:data<=16'd4519;
      6976:data<=16'd4730;
      6977:data<=16'd4955;
      6978:data<=16'd4585;
      6979:data<=16'd4592;
      6980:data<=16'd4049;
      6981:data<=16'd3997;
      6982:data<=16'd4581;
      6983:data<=16'd3914;
      6984:data<=16'd4623;
      6985:data<=16'd4831;
      6986:data<=16'd3976;
      6987:data<=16'd6660;
      6988:data<=16'd3993;
      6989:data<=-16'd5621;
      6990:data<=-16'd7876;
      6991:data<=-16'd6078;
      6992:data<=-16'd7245;
      6993:data<=-16'd6840;
      6994:data<=-16'd6269;
      6995:data<=-16'd5862;
      6996:data<=-16'd4567;
      6997:data<=-16'd4801;
      6998:data<=-16'd4390;
      6999:data<=-16'd3927;
      7000:data<=-16'd4356;
      7001:data<=-16'd3281;
      7002:data<=-16'd2786;
      7003:data<=-16'd1980;
      7004:data<=-16'd234;
      7005:data<=-16'd705;
      7006:data<=-16'd684;
      7007:data<=16'd29;
      7008:data<=-16'd423;
      7009:data<=16'd41;
      7010:data<=-16'd255;
      7011:data<=-16'd936;
      7012:data<=-16'd274;
      7013:data<=-16'd323;
      7014:data<=16'd36;
      7015:data<=16'd290;
      7016:data<=-16'd144;
      7017:data<=16'd772;
      7018:data<=16'd343;
      7019:data<=16'd92;
      7020:data<=16'd2591;
      7021:data<=16'd3806;
      7022:data<=16'd4646;
      7023:data<=16'd5598;
      7024:data<=16'd5036;
      7025:data<=16'd5203;
      7026:data<=16'd4475;
      7027:data<=16'd4196;
      7028:data<=16'd5415;
      7029:data<=16'd3668;
      7030:data<=16'd6564;
      7031:data<=16'd15807;
      7032:data<=16'd18108;
      7033:data<=16'd16202;
      7034:data<=16'd16575;
      7035:data<=16'd15403;
      7036:data<=16'd15318;
      7037:data<=16'd16765;
      7038:data<=16'd16040;
      7039:data<=16'd15226;
      7040:data<=16'd14665;
      7041:data<=16'd13920;
      7042:data<=16'd13662;
      7043:data<=16'd12925;
      7044:data<=16'd12398;
      7045:data<=16'd11806;
      7046:data<=16'd10790;
      7047:data<=16'd10699;
      7048:data<=16'd10715;
      7049:data<=16'd10501;
      7050:data<=16'd10100;
      7051:data<=16'd9175;
      7052:data<=16'd9313;
      7053:data<=16'd10138;
      7054:data<=16'd10326;
      7055:data<=16'd10070;
      7056:data<=16'd9454;
      7057:data<=16'd9323;
      7058:data<=16'd8874;
      7059:data<=16'd7758;
      7060:data<=16'd7897;
      7061:data<=16'd7785;
      7062:data<=16'd7036;
      7063:data<=16'd7106;
      7064:data<=16'd6376;
      7065:data<=16'd5947;
      7066:data<=16'd6158;
      7067:data<=16'd5171;
      7068:data<=16'd5313;
      7069:data<=16'd5565;
      7070:data<=16'd5147;
      7071:data<=16'd6231;
      7072:data<=16'd1973;
      7073:data<=-16'd7692;
      7074:data<=-16'd10871;
      7075:data<=-16'd9386;
      7076:data<=-16'd10114;
      7077:data<=-16'd10064;
      7078:data<=-16'd9271;
      7079:data<=-16'd9498;
      7080:data<=-16'd9127;
      7081:data<=-16'd8760;
      7082:data<=-16'd8796;
      7083:data<=-16'd8317;
      7084:data<=-16'd7793;
      7085:data<=-16'd7641;
      7086:data<=-16'd7110;
      7087:data<=-16'd5627;
      7088:data<=-16'd4739;
      7089:data<=-16'd5080;
      7090:data<=-16'd5015;
      7091:data<=-16'd4755;
      7092:data<=-16'd4678;
      7093:data<=-16'd4628;
      7094:data<=-16'd5198;
      7095:data<=-16'd4998;
      7096:data<=-16'd4179;
      7097:data<=-16'd4458;
      7098:data<=-16'd4613;
      7099:data<=-16'd4579;
      7100:data<=-16'd4629;
      7101:data<=-16'd4344;
      7102:data<=-16'd5016;
      7103:data<=-16'd4378;
      7104:data<=-16'd1782;
      7105:data<=-16'd1278;
      7106:data<=-16'd1486;
      7107:data<=-16'd1306;
      7108:data<=-16'd2088;
      7109:data<=-16'd1788;
      7110:data<=-16'd1811;
      7111:data<=-16'd2241;
      7112:data<=-16'd1418;
      7113:data<=-16'd2517;
      7114:data<=-16'd56;
      7115:data<=16'd8968;
      7116:data<=16'd12349;
      7117:data<=16'd10235;
      7118:data<=16'd10649;
      7119:data<=16'd10411;
      7120:data<=16'd10402;
      7121:data<=16'd12417;
      7122:data<=16'd12624;
      7123:data<=16'd12260;
      7124:data<=16'd11841;
      7125:data<=16'd10592;
      7126:data<=16'd10334;
      7127:data<=16'd9721;
      7128:data<=16'd8854;
      7129:data<=16'd8883;
      7130:data<=16'd8094;
      7131:data<=16'd7242;
      7132:data<=16'd7031;
      7133:data<=16'd6866;
      7134:data<=16'd6625;
      7135:data<=16'd5574;
      7136:data<=16'd5794;
      7137:data<=16'd7383;
      7138:data<=16'd7110;
      7139:data<=16'd6484;
      7140:data<=16'd6373;
      7141:data<=16'd5454;
      7142:data<=16'd5127;
      7143:data<=16'd5093;
      7144:data<=16'd4664;
      7145:data<=16'd4246;
      7146:data<=16'd3565;
      7147:data<=16'd3385;
      7148:data<=16'd2825;
      7149:data<=16'd1927;
      7150:data<=16'd2300;
      7151:data<=16'd1902;
      7152:data<=16'd1275;
      7153:data<=16'd2000;
      7154:data<=16'd2396;
      7155:data<=16'd3128;
      7156:data<=16'd403;
      7157:data<=-16'd8091;
      7158:data<=-16'd12420;
      7159:data<=-16'd11041;
      7160:data<=-16'd11260;
      7161:data<=-16'd11380;
      7162:data<=-16'd10611;
      7163:data<=-16'd10827;
      7164:data<=-16'd10308;
      7165:data<=-16'd10299;
      7166:data<=-16'd10827;
      7167:data<=-16'd9861;
      7168:data<=-16'd9561;
      7169:data<=-16'd9749;
      7170:data<=-16'd8216;
      7171:data<=-16'd7204;
      7172:data<=-16'd8078;
      7173:data<=-16'd8784;
      7174:data<=-16'd8922;
      7175:data<=-16'd9212;
      7176:data<=-16'd8956;
      7177:data<=-16'd8505;
      7178:data<=-16'd8701;
      7179:data<=-16'd8661;
      7180:data<=-16'd8548;
      7181:data<=-16'd8475;
      7182:data<=-16'd7856;
      7183:data<=-16'd7920;
      7184:data<=-16'd8194;
      7185:data<=-16'd7929;
      7186:data<=-16'd7859;
      7187:data<=-16'd6337;
      7188:data<=-16'd4713;
      7189:data<=-16'd5324;
      7190:data<=-16'd5324;
      7191:data<=-16'd5065;
      7192:data<=-16'd5479;
      7193:data<=-16'd4864;
      7194:data<=-16'd5347;
      7195:data<=-16'd5470;
      7196:data<=-16'd4194;
      7197:data<=-16'd5673;
      7198:data<=-16'd3797;
      7199:data<=16'd4863;
      7200:data<=16'd9247;
      7201:data<=16'd7858;
      7202:data<=16'd7339;
      7203:data<=16'd7576;
      7204:data<=16'd8378;
      7205:data<=16'd9200;
      7206:data<=16'd8660;
      7207:data<=16'd8022;
      7208:data<=16'd7177;
      7209:data<=16'd6464;
      7210:data<=16'd6543;
      7211:data<=16'd5965;
      7212:data<=16'd5336;
      7213:data<=16'd4927;
      7214:data<=16'd3956;
      7215:data<=16'd3873;
      7216:data<=16'd4255;
      7217:data<=16'd3892;
      7218:data<=16'd3489;
      7219:data<=16'd2855;
      7220:data<=16'd2943;
      7221:data<=16'd4836;
      7222:data<=16'd6287;
      7223:data<=16'd6111;
      7224:data<=16'd5833;
      7225:data<=16'd5944;
      7226:data<=16'd5432;
      7227:data<=16'd4490;
      7228:data<=16'd4464;
      7229:data<=16'd4582;
      7230:data<=16'd3926;
      7231:data<=16'd3535;
      7232:data<=16'd3168;
      7233:data<=16'd2692;
      7234:data<=16'd2585;
      7235:data<=16'd2041;
      7236:data<=16'd1858;
      7237:data<=16'd1889;
      7238:data<=16'd1105;
      7239:data<=16'd1436;
      7240:data<=-16'd652;
      7241:data<=-16'd8648;
      7242:data<=-16'd13781;
      7243:data<=-16'd12677;
      7244:data<=-16'd12527;
      7245:data<=-16'd13021;
      7246:data<=-16'd11985;
      7247:data<=-16'd11790;
      7248:data<=-16'd11600;
      7249:data<=-16'd11018;
      7250:data<=-16'd11186;
      7251:data<=-16'd11121;
      7252:data<=-16'd10757;
      7253:data<=-16'd10546;
      7254:data<=-16'd10774;
      7255:data<=-16'd11456;
      7256:data<=-16'd11342;
      7257:data<=-16'd11032;
      7258:data<=-16'd11262;
      7259:data<=-16'd10881;
      7260:data<=-16'd10351;
      7261:data<=-16'd10061;
      7262:data<=-16'd9589;
      7263:data<=-16'd9567;
      7264:data<=-16'd9714;
      7265:data<=-16'd9500;
      7266:data<=-16'd9109;
      7267:data<=-16'd8901;
      7268:data<=-16'd9092;
      7269:data<=-16'd8737;
      7270:data<=-16'd8645;
      7271:data<=-16'd10329;
      7272:data<=-16'd11740;
      7273:data<=-16'd11635;
      7274:data<=-16'd11069;
      7275:data<=-16'd10680;
      7276:data<=-16'd10672;
      7277:data<=-16'd9964;
      7278:data<=-16'd9107;
      7279:data<=-16'd9048;
      7280:data<=-16'd8411;
      7281:data<=-16'd8351;
      7282:data<=-16'd6545;
      7283:data<=16'd948;
      7284:data<=16'd6302;
      7285:data<=16'd5454;
      7286:data<=16'd5204;
      7287:data<=16'd4839;
      7288:data<=16'd2836;
      7289:data<=16'd2692;
      7290:data<=16'd2867;
      7291:data<=16'd2601;
      7292:data<=16'd2904;
      7293:data<=16'd2510;
      7294:data<=16'd2388;
      7295:data<=16'd2728;
      7296:data<=16'd2463;
      7297:data<=16'd2170;
      7298:data<=16'd1847;
      7299:data<=16'd2118;
      7300:data<=16'd2481;
      7301:data<=16'd1903;
      7302:data<=16'd2100;
      7303:data<=16'd2052;
      7304:data<=16'd517;
      7305:data<=-16'd61;
      7306:data<=16'd259;
      7307:data<=16'd496;
      7308:data<=16'd663;
      7309:data<=16'd449;
      7310:data<=16'd749;
      7311:data<=16'd846;
      7312:data<=16'd461;
      7313:data<=16'd863;
      7314:data<=16'd764;
      7315:data<=16'd752;
      7316:data<=16'd1245;
      7317:data<=16'd268;
      7318:data<=16'd168;
      7319:data<=16'd1033;
      7320:data<=16'd36;
      7321:data<=-16'd732;
      7322:data<=-16'd444;
      7323:data<=16'd584;
      7324:data<=16'd323;
      7325:data<=-16'd6199;
      7326:data<=-16'd12845;
      7327:data<=-16'd12478;
      7328:data<=-16'd11488;
      7329:data<=-16'd11820;
      7330:data<=-16'd10561;
      7331:data<=-16'd10248;
      7332:data<=-16'd10285;
      7333:data<=-16'd9494;
      7334:data<=-16'd9339;
      7335:data<=-16'd8766;
      7336:data<=-16'd8113;
      7337:data<=-16'd8522;
      7338:data<=-16'd9019;
      7339:data<=-16'd8963;
      7340:data<=-16'd8272;
      7341:data<=-16'd8028;
      7342:data<=-16'd8294;
      7343:data<=-16'd7702;
      7344:data<=-16'd7053;
      7345:data<=-16'd6667;
      7346:data<=-16'd6232;
      7347:data<=-16'd6260;
      7348:data<=-16'd5920;
      7349:data<=-16'd5494;
      7350:data<=-16'd5430;
      7351:data<=-16'd4893;
      7352:data<=-16'd4658;
      7353:data<=-16'd4817;
      7354:data<=-16'd5372;
      7355:data<=-16'd6398;
      7356:data<=-16'd6009;
      7357:data<=-16'd5409;
      7358:data<=-16'd5453;
      7359:data<=-16'd4513;
      7360:data<=-16'd4493;
      7361:data<=-16'd4639;
      7362:data<=-16'd3497;
      7363:data<=-16'd3603;
      7364:data<=-16'd2960;
      7365:data<=-16'd2123;
      7366:data<=-16'd2446;
      7367:data<=16'd3366;
      7368:data<=16'd11518;
      7369:data<=16'd12251;
      7370:data<=16'd10683;
      7371:data<=16'd9400;
      7372:data<=16'd6263;
      7373:data<=16'd5436;
      7374:data<=16'd6078;
      7375:data<=16'd5623;
      7376:data<=16'd5598;
      7377:data<=16'd5448;
      7378:data<=16'd5426;
      7379:data<=16'd5380;
      7380:data<=16'd4422;
      7381:data<=16'd4220;
      7382:data<=16'd4487;
      7383:data<=16'd4868;
      7384:data<=16'd5412;
      7385:data<=16'd4933;
      7386:data<=16'd4922;
      7387:data<=16'd4478;
      7388:data<=16'd2420;
      7389:data<=16'd2234;
      7390:data<=16'd2763;
      7391:data<=16'd2331;
      7392:data<=16'd2852;
      7393:data<=16'd2664;
      7394:data<=16'd2074;
      7395:data<=16'd2409;
      7396:data<=16'd2124;
      7397:data<=16'd2399;
      7398:data<=16'd2767;
      7399:data<=16'd2402;
      7400:data<=16'd2955;
      7401:data<=16'd2852;
      7402:data<=16'd2799;
      7403:data<=16'd3368;
      7404:data<=16'd1812;
      7405:data<=16'd734;
      7406:data<=16'd403;
      7407:data<=-16'd349;
      7408:data<=16'd531;
      7409:data<=-16'd3732;
      7410:data<=-16'd12602;
      7411:data<=-16'd13940;
      7412:data<=-16'd11658;
      7413:data<=-16'd12196;
      7414:data<=-16'd11365;
      7415:data<=-16'd10480;
      7416:data<=-16'd10220;
      7417:data<=-16'd9139;
      7418:data<=-16'd9165;
      7419:data<=-16'd8660;
      7420:data<=-16'd8264;
      7421:data<=-16'd9144;
      7422:data<=-16'd7658;
      7423:data<=-16'd5783;
      7424:data<=-16'd5994;
      7425:data<=-16'd5950;
      7426:data<=-16'd5874;
      7427:data<=-16'd5656;
      7428:data<=-16'd4928;
      7429:data<=-16'd4570;
      7430:data<=-16'd4067;
      7431:data<=-16'd3964;
      7432:data<=-16'd3797;
      7433:data<=-16'd3107;
      7434:data<=-16'd3489;
      7435:data<=-16'd3250;
      7436:data<=-16'd2080;
      7437:data<=-16'd2570;
      7438:data<=-16'd3694;
      7439:data<=-16'd4275;
      7440:data<=-16'd4049;
      7441:data<=-16'd3350;
      7442:data<=-16'd3566;
      7443:data<=-16'd3298;
      7444:data<=-16'd2535;
      7445:data<=-16'd2355;
      7446:data<=-16'd1679;
      7447:data<=-16'd1727;
      7448:data<=-16'd1447;
      7449:data<=-16'd391;
      7450:data<=-16'd1195;
      7451:data<=16'd2763;
      7452:data<=16'd12079;
      7453:data<=16'd14449;
      7454:data<=16'd11664;
      7455:data<=16'd11112;
      7456:data<=16'd10288;
      7457:data<=16'd9811;
      7458:data<=16'd10187;
      7459:data<=16'd9538;
      7460:data<=16'd9661;
      7461:data<=16'd9838;
      7462:data<=16'd9163;
      7463:data<=16'd8799;
      7464:data<=16'd8331;
      7465:data<=16'd8290;
      7466:data<=16'd8305;
      7467:data<=16'd7824;
      7468:data<=16'd7808;
      7469:data<=16'd7779;
      7470:data<=16'd8019;
      7471:data<=16'd7285;
      7472:data<=16'd4511;
      7473:data<=16'd3486;
      7474:data<=16'd3767;
      7475:data<=16'd3087;
      7476:data<=16'd3286;
      7477:data<=16'd3306;
      7478:data<=16'd3028;
      7479:data<=16'd3432;
      7480:data<=16'd2895;
      7481:data<=16'd2869;
      7482:data<=16'd3260;
      7483:data<=16'd3015;
      7484:data<=16'd3758;
      7485:data<=16'd3665;
      7486:data<=16'd3315;
      7487:data<=16'd3553;
      7488:data<=16'd1671;
      7489:data<=16'd1178;
      7490:data<=16'd1789;
      7491:data<=16'd755;
      7492:data<=16'd1785;
      7493:data<=-16'd1745;
      7494:data<=-16'd11247;
      7495:data<=-16'd13053;
      7496:data<=-16'd10721;
      7497:data<=-16'd11996;
      7498:data<=-16'd11254;
      7499:data<=-16'd9894;
      7500:data<=-16'd10025;
      7501:data<=-16'd9354;
      7502:data<=-16'd9313;
      7503:data<=-16'd8596;
      7504:data<=-16'd7542;
      7505:data<=-16'd7736;
      7506:data<=-16'd6842;
      7507:data<=-16'd6068;
      7508:data<=-16'd5880;
      7509:data<=-16'd5128;
      7510:data<=-16'd5330;
      7511:data<=-16'd5169;
      7512:data<=-16'd4622;
      7513:data<=-16'd4613;
      7514:data<=-16'd3856;
      7515:data<=-16'd4041;
      7516:data<=-16'd4282;
      7517:data<=-16'd3072;
      7518:data<=-16'd2722;
      7519:data<=-16'd2185;
      7520:data<=-16'd1861;
      7521:data<=-16'd2076;
      7522:data<=16'd385;
      7523:data<=16'd2537;
      7524:data<=16'd2538;
      7525:data<=16'd2719;
      7526:data<=16'd2268;
      7527:data<=16'd2473;
      7528:data<=16'd2790;
      7529:data<=16'd1968;
      7530:data<=16'd2692;
      7531:data<=16'd2971;
      7532:data<=16'd3052;
      7533:data<=16'd3871;
      7534:data<=16'd2270;
      7535:data<=16'd6065;
      7536:data<=16'd15858;
      7537:data<=16'd18304;
      7538:data<=16'd17106;
      7539:data<=16'd18471;
      7540:data<=16'd17529;
      7541:data<=16'd16671;
      7542:data<=16'd16835;
      7543:data<=16'd15881;
      7544:data<=16'd15920;
      7545:data<=16'd15359;
      7546:data<=16'd14442;
      7547:data<=16'd14600;
      7548:data<=16'd13667;
      7549:data<=16'd12954;
      7550:data<=16'd12750;
      7551:data<=16'd12284;
      7552:data<=16'd12463;
      7553:data<=16'd11646;
      7554:data<=16'd11459;
      7555:data<=16'd12759;
      7556:data<=16'd12502;
      7557:data<=16'd12343;
      7558:data<=16'd12020;
      7559:data<=16'd10548;
      7560:data<=16'd10927;
      7561:data<=16'd10989;
      7562:data<=16'd9861;
      7563:data<=16'd9829;
      7564:data<=16'd9241;
      7565:data<=16'd8986;
      7566:data<=16'd9150;
      7567:data<=16'd8257;
      7568:data<=16'd8429;
      7569:data<=16'd8173;
      7570:data<=16'd7318;
      7571:data<=16'd8211;
      7572:data<=16'd7982;
      7573:data<=16'd6764;
      7574:data<=16'd5682;
      7575:data<=16'd4742;
      7576:data<=16'd6012;
      7577:data<=16'd2358;
      7578:data<=-16'd7512;
      7579:data<=-16'd10141;
      7580:data<=-16'd7477;
      7581:data<=-16'd8417;
      7582:data<=-16'd8746;
      7583:data<=-16'd8078;
      7584:data<=-16'd8281;
      7585:data<=-16'd7412;
      7586:data<=-16'd7547;
      7587:data<=-16'd7726;
      7588:data<=-16'd5833;
      7589:data<=-16'd4698;
      7590:data<=-16'd4381;
      7591:data<=-16'd3970;
      7592:data<=-16'd4073;
      7593:data<=-16'd3877;
      7594:data<=-16'd3668;
      7595:data<=-16'd3765;
      7596:data<=-16'd3648;
      7597:data<=-16'd3542;
      7598:data<=-16'd3350;
      7599:data<=-16'd3336;
      7600:data<=-16'd3298;
      7601:data<=-16'd2901;
      7602:data<=-16'd3243;
      7603:data<=-16'd3636;
      7604:data<=-16'd2657;
      7605:data<=-16'd1181;
      7606:data<=-16'd491;
      7607:data<=-16'd851;
      7608:data<=-16'd1122;
      7609:data<=-16'd1005;
      7610:data<=-16'd1213;
      7611:data<=-16'd1051;
      7612:data<=-16'd949;
      7613:data<=-16'd1048;
      7614:data<=-16'd772;
      7615:data<=-16'd1298;
      7616:data<=-16'd738;
      7617:data<=16'd176;
      7618:data<=-16'd1521;
      7619:data<=16'd2015;
      7620:data<=16'd11160;
      7621:data<=16'd13858;
      7622:data<=16'd13571;
      7623:data<=16'd16198;
      7624:data<=16'd16031;
      7625:data<=16'd14848;
      7626:data<=16'd15148;
      7627:data<=16'd14211;
      7628:data<=16'd13729;
      7629:data<=16'd13145;
      7630:data<=16'd11690;
      7631:data<=16'd11503;
      7632:data<=16'd11133;
      7633:data<=16'd10499;
      7634:data<=16'd10264;
      7635:data<=16'd9415;
      7636:data<=16'd8842;
      7637:data<=16'd8272;
      7638:data<=16'd8555;
      7639:data<=16'd10181;
      7640:data<=16'd9946;
      7641:data<=16'd9083;
      7642:data<=16'd8900;
      7643:data<=16'd7733;
      7644:data<=16'd7482;
      7645:data<=16'd7617;
      7646:data<=16'd6942;
      7647:data<=16'd6834;
      7648:data<=16'd5938;
      7649:data<=16'd5234;
      7650:data<=16'd5626;
      7651:data<=16'd5300;
      7652:data<=16'd5429;
      7653:data<=16'd5021;
      7654:data<=16'd4132;
      7655:data<=16'd5122;
      7656:data<=16'd5392;
      7657:data<=16'd5247;
      7658:data<=16'd4934;
      7659:data<=16'd3330;
      7660:data<=16'd4246;
      7661:data<=16'd1472;
      7662:data<=-16'd8158;
      7663:data<=-16'd11494;
      7664:data<=-16'd9776;
      7665:data<=-16'd10660;
      7666:data<=-16'd10031;
      7667:data<=-16'd9697;
      7668:data<=-16'd10313;
      7669:data<=-16'd9273;
      7670:data<=-16'd9855;
      7671:data<=-16'd9303;
      7672:data<=-16'd7318;
      7673:data<=-16'd8510;
      7674:data<=-16'd9012;
      7675:data<=-16'd8185;
      7676:data<=-16'd8307;
      7677:data<=-16'd7635;
      7678:data<=-16'd7602;
      7679:data<=-16'd7674;
      7680:data<=-16'd6984;
      7681:data<=-16'd7366;
      7682:data<=-16'd7210;
      7683:data<=-16'd7057;
      7684:data<=-16'd7394;
      7685:data<=-16'd6370;
      7686:data<=-16'd6355;
      7687:data<=-16'd6865;
      7688:data<=-16'd5577;
      7689:data<=-16'd4219;
      7690:data<=-16'd3422;
      7691:data<=-16'd3697;
      7692:data<=-16'd4200;
      7693:data<=-16'd3692;
      7694:data<=-16'd3956;
      7695:data<=-16'd3867;
      7696:data<=-16'd3283;
      7697:data<=-16'd3700;
      7698:data<=-16'd3392;
      7699:data<=-16'd3507;
      7700:data<=-16'd3312;
      7701:data<=-16'd2158;
      7702:data<=-16'd3647;
      7703:data<=-16'd860;
      7704:data<=16'd8490;
      7705:data<=16'd12266;
      7706:data<=16'd11506;
      7707:data<=16'd12123;
      7708:data<=16'd11264;
      7709:data<=16'd10812;
      7710:data<=16'd10880;
      7711:data<=16'd9442;
      7712:data<=16'd9300;
      7713:data<=16'd9297;
      7714:data<=16'd8390;
      7715:data<=16'd8011;
      7716:data<=16'd7165;
      7717:data<=16'd6739;
      7718:data<=16'd7019;
      7719:data<=16'd6786;
      7720:data<=16'd6096;
      7721:data<=16'd5227;
      7722:data<=16'd6570;
      7723:data<=16'd8990;
      7724:data<=16'd8731;
      7725:data<=16'd8184;
      7726:data<=16'd8304;
      7727:data<=16'd7586;
      7728:data<=16'd7319;
      7729:data<=16'd6725;
      7730:data<=16'd5893;
      7731:data<=16'd5920;
      7732:data<=16'd5544;
      7733:data<=16'd5187;
      7734:data<=16'd4792;
      7735:data<=16'd4340;
      7736:data<=16'd4508;
      7737:data<=16'd3733;
      7738:data<=16'd3824;
      7739:data<=16'd5263;
      7740:data<=16'd4813;
      7741:data<=16'd4494;
      7742:data<=16'd4161;
      7743:data<=16'd3183;
      7744:data<=16'd4426;
      7745:data<=16'd873;
      7746:data<=-16'd8592;
      7747:data<=-16'd11565;
      7748:data<=-16'd9702;
      7749:data<=-16'd10273;
      7750:data<=-16'd10345;
      7751:data<=-16'd10006;
      7752:data<=-16'd10073;
      7753:data<=-16'd9345;
      7754:data<=-16'd9538;
      7755:data<=-16'd9106;
      7756:data<=-16'd7131;
      7757:data<=-16'd6410;
      7758:data<=-16'd6432;
      7759:data<=-16'd6272;
      7760:data<=-16'd6313;
      7761:data<=-16'd6046;
      7762:data<=-16'd5771;
      7763:data<=-16'd5589;
      7764:data<=-16'd5592;
      7765:data<=-16'd5873;
      7766:data<=-16'd5524;
      7767:data<=-16'd5142;
      7768:data<=-16'd5416;
      7769:data<=-16'd5571;
      7770:data<=-16'd5435;
      7771:data<=-16'd4990;
      7772:data<=-16'd4868;
      7773:data<=-16'd5841;
      7774:data<=-16'd6878;
      7775:data<=-16'd7054;
      7776:data<=-16'd6567;
      7777:data<=-16'd6338;
      7778:data<=-16'd6601;
      7779:data<=-16'd6188;
      7780:data<=-16'd5644;
      7781:data<=-16'd5556;
      7782:data<=-16'd5483;
      7783:data<=-16'd6011;
      7784:data<=-16'd5341;
      7785:data<=-16'd4208;
      7786:data<=-16'd5495;
      7787:data<=-16'd2517;
      7788:data<=16'd5761;
      7789:data<=16'd8076;
      7790:data<=16'd5779;
      7791:data<=16'd5861;
      7792:data<=16'd5679;
      7793:data<=16'd5388;
      7794:data<=16'd5698;
      7795:data<=16'd4872;
      7796:data<=16'd4904;
      7797:data<=16'd4754;
      7798:data<=16'd3533;
      7799:data<=16'd3532;
      7800:data<=16'd3278;
      7801:data<=16'd2845;
      7802:data<=16'd2983;
      7803:data<=16'd2355;
      7804:data<=16'd2426;
      7805:data<=16'd1794;
      7806:data<=-16'd555;
      7807:data<=-16'd870;
      7808:data<=-16'd482;
      7809:data<=-16'd793;
      7810:data<=-16'd155;
      7811:data<=-16'd467;
      7812:data<=-16'd1257;
      7813:data<=-16'd1134;
      7814:data<=-16'd1489;
      7815:data<=-16'd1556;
      7816:data<=-16'd1342;
      7817:data<=-16'd1347;
      7818:data<=-16'd1089;
      7819:data<=-16'd1230;
      7820:data<=-16'd957;
      7821:data<=-16'd1111;
      7822:data<=-16'd2743;
      7823:data<=-16'd3093;
      7824:data<=-16'd2378;
      7825:data<=-16'd1888;
      7826:data<=-16'd1847;
      7827:data<=-16'd2487;
      7828:data<=-16'd1666;
      7829:data<=-16'd4152;
      7830:data<=-16'd12845;
      7831:data<=-16'd16739;
      7832:data<=-16'd14810;
      7833:data<=-16'd14780;
      7834:data<=-16'd14410;
      7835:data<=-16'd13872;
      7836:data<=-16'd14108;
      7837:data<=-16'd12537;
      7838:data<=-16'd12536;
      7839:data<=-16'd13903;
      7840:data<=-16'd13567;
      7841:data<=-16'd13368;
      7842:data<=-16'd12810;
      7843:data<=-16'd12026;
      7844:data<=-16'd11920;
      7845:data<=-16'd11075;
      7846:data<=-16'd10743;
      7847:data<=-16'd10305;
      7848:data<=-16'd9150;
      7849:data<=-16'd9523;
      7850:data<=-16'd9294;
      7851:data<=-16'd8338;
      7852:data<=-16'd8906;
      7853:data<=-16'd8520;
      7854:data<=-16'd7545;
      7855:data<=-16'd8041;
      7856:data<=-16'd8655;
      7857:data<=-16'd8751;
      7858:data<=-16'd8316;
      7859:data<=-16'd7971;
      7860:data<=-16'd7931;
      7861:data<=-16'd7448;
      7862:data<=-16'd7150;
      7863:data<=-16'd6593;
      7864:data<=-16'd5990;
      7865:data<=-16'd5941;
      7866:data<=-16'd5183;
      7867:data<=-16'd5177;
      7868:data<=-16'd5154;
      7869:data<=-16'd3847;
      7870:data<=-16'd4626;
      7871:data<=-16'd2215;
      7872:data<=16'd5914;
      7873:data<=16'd8143;
      7874:data<=16'd5086;
      7875:data<=16'd5162;
      7876:data<=16'd5598;
      7877:data<=16'd5427;
      7878:data<=16'd5435;
      7879:data<=16'd4299;
      7880:data<=16'd4449;
      7881:data<=16'd4984;
      7882:data<=16'd4197;
      7883:data<=16'd4049;
      7884:data<=16'd3821;
      7885:data<=16'd3453;
      7886:data<=16'd3721;
      7887:data<=16'd3586;
      7888:data<=16'd3310;
      7889:data<=16'd2187;
      7890:data<=16'd699;
      7891:data<=16'd1175;
      7892:data<=16'd1745;
      7893:data<=16'd1221;
      7894:data<=16'd1236;
      7895:data<=16'd1262;
      7896:data<=16'd913;
      7897:data<=16'd693;
      7898:data<=16'd519;
      7899:data<=16'd432;
      7900:data<=16'd514;
      7901:data<=16'd936;
      7902:data<=16'd799;
      7903:data<=16'd265;
      7904:data<=16'd914;
      7905:data<=16'd672;
      7906:data<=-16'd1290;
      7907:data<=-16'd1942;
      7908:data<=-16'd1751;
      7909:data<=-16'd1803;
      7910:data<=-16'd1670;
      7911:data<=-16'd1798;
      7912:data<=-16'd1281;
      7913:data<=-16'd3195;
      7914:data<=-16'd10430;
      7915:data<=-16'd15261;
      7916:data<=-16'd14240;
      7917:data<=-16'd13453;
      7918:data<=-16'd13485;
      7919:data<=-16'd13044;
      7920:data<=-16'd12631;
      7921:data<=-16'd11189;
      7922:data<=-16'd11107;
      7923:data<=-16'd12149;
      7924:data<=-16'd10258;
      7925:data<=-16'd8470;
      7926:data<=-16'd8860;
      7927:data<=-16'd8243;
      7928:data<=-16'd7498;
      7929:data<=-16'd7415;
      7930:data<=-16'd7006;
      7931:data<=-16'd7004;
      7932:data<=-16'd6561;
      7933:data<=-16'd5817;
      7934:data<=-16'd5785;
      7935:data<=-16'd5186;
      7936:data<=-16'd4745;
      7937:data<=-16'd4789;
      7938:data<=-16'd3880;
      7939:data<=-16'd3835;
      7940:data<=-16'd4943;
      7941:data<=-16'd4842;
      7942:data<=-16'd4414;
      7943:data<=-16'd4444;
      7944:data<=-16'd3888;
      7945:data<=-16'd3541;
      7946:data<=-16'd3814;
      7947:data<=-16'd3392;
      7948:data<=-16'd2737;
      7949:data<=-16'd2708;
      7950:data<=-16'd2378;
      7951:data<=-16'd2181;
      7952:data<=-16'd1992;
      7953:data<=-16'd588;
      7954:data<=-16'd420;
      7955:data<=16'd135;
      7956:data<=16'd6031;
      7957:data<=16'd11309;
      7958:data<=16'd10986;
      7959:data<=16'd10457;
      7960:data<=16'd10677;
      7961:data<=16'd10161;
      7962:data<=16'd10014;
      7963:data<=16'd9157;
      7964:data<=16'd8719;
      7965:data<=16'd9091;
      7966:data<=16'd8147;
      7967:data<=16'd7776;
      7968:data<=16'd8156;
      7969:data<=16'd7561;
      7970:data<=16'd7454;
      7971:data<=16'd7818;
      7972:data<=16'd7401;
      7973:data<=16'd5398;
      7974:data<=16'd2749;
      7975:data<=16'd2513;
      7976:data<=16'd3096;
      7977:data<=16'd2549;
      7978:data<=16'd2849;
      7979:data<=16'd3011;
      7980:data<=16'd2537;
      7981:data<=16'd2572;
      7982:data<=16'd2188;
      7983:data<=16'd2177;
      7984:data<=16'd2672;
      7985:data<=16'd2631;
      7986:data<=16'd2567;
      7987:data<=16'd2208;
      7988:data<=16'd2300;
      7989:data<=16'd2150;
      7990:data<=16'd420;
      7991:data<=16'd165;
      7992:data<=16'd690;
      7993:data<=16'd214;
      7994:data<=16'd557;
      7995:data<=-16'd243;
      7996:data<=-16'd664;
      7997:data<=-16'd449;
      7998:data<=-16'd6927;
      7999:data<=-16'd14075;
      8000:data<=-16'd13409;
      8001:data<=-16'd12041;
      8002:data<=-16'd12308;
      8003:data<=-16'd11505;
      8004:data<=-16'd10921;
      8005:data<=-16'd9687;
      8006:data<=-16'd9623;
      8007:data<=-16'd11010;
      8008:data<=-16'd10235;
      8009:data<=-16'd9514;
      8010:data<=-16'd9486;
      8011:data<=-16'd8523;
      8012:data<=-16'd8520;
      8013:data<=-16'd8475;
      8014:data<=-16'd7765;
      8015:data<=-16'd7442;
      8016:data<=-16'd6684;
      8017:data<=-16'd6595;
      8018:data<=-16'd6646;
      8019:data<=-16'd5708;
      8020:data<=-16'd5327;
      8021:data<=-16'd4654;
      8022:data<=-16'd4532;
      8023:data<=-16'd5709;
      8024:data<=-16'd4667;
      8025:data<=-16'd3048;
      8026:data<=-16'd3162;
      8027:data<=-16'd2602;
      8028:data<=-16'd2014;
      8029:data<=-16'd2070;
      8030:data<=-16'd1782;
      8031:data<=-16'd1419;
      8032:data<=-16'd820;
      8033:data<=-16'd685;
      8034:data<=-16'd506;
      8035:data<=16'd21;
      8036:data<=-16'd555;
      8037:data<=16'd132;
      8038:data<=16'd1183;
      8039:data<=16'd1033;
      8040:data<=16'd6575;
      8041:data<=16'd14478;
      8042:data<=16'd14839;
      8043:data<=16'd13195;
      8044:data<=16'd14187;
      8045:data<=16'd13805;
      8046:data<=16'd12833;
      8047:data<=16'd12422;
      8048:data<=16'd12284;
      8049:data<=16'd12475;
      8050:data<=16'd11614;
      8051:data<=16'd10934;
      8052:data<=16'd10966;
      8053:data<=16'd10520;
      8054:data<=16'd10564;
      8055:data<=16'd10580;
      8056:data<=16'd10804;
      8057:data<=16'd11949;
      8058:data<=16'd11779;
      8059:data<=16'd11151;
      8060:data<=16'd11126;
      8061:data<=16'd10325;
      8062:data<=16'd10047;
      8063:data<=16'd10064;
      8064:data<=16'd9567;
      8065:data<=16'd9662;
      8066:data<=16'd9333;
      8067:data<=16'd9004;
      8068:data<=16'd9235;
      8069:data<=16'd8737;
      8070:data<=16'd8405;
      8071:data<=16'd7890;
      8072:data<=16'd7876;
      8073:data<=16'd9324;
      8074:data<=16'd8434;
      8075:data<=16'd6734;
      8076:data<=16'd6995;
      8077:data<=16'd6367;
      8078:data<=16'd6305;
      8079:data<=16'd6200;
      8080:data<=16'd4872;
      8081:data<=16'd5518;
      8082:data<=16'd1293;
      8083:data<=-16'd7900;
      8084:data<=-16'd9273;
      8085:data<=-16'd6986;
      8086:data<=-16'd7993;
      8087:data<=-16'd7685;
      8088:data<=-16'd7260;
      8089:data<=-16'd6516;
      8090:data<=-16'd4023;
      8091:data<=-16'd3576;
      8092:data<=-16'd3377;
      8093:data<=-16'd2887;
      8094:data<=-16'd3771;
      8095:data<=-16'd3295;
      8096:data<=-16'd3052;
      8097:data<=-16'd3495;
      8098:data<=-16'd2540;
      8099:data<=-16'd2648;
      8100:data<=-16'd2802;
      8101:data<=-16'd1917;
      8102:data<=-16'd1891;
      8103:data<=-16'd1303;
      8104:data<=-16'd1077;
      8105:data<=-16'd1782;
      8106:data<=-16'd840;
      8107:data<=16'd453;
      8108:data<=16'd948;
      8109:data<=16'd886;
      8110:data<=16'd520;
      8111:data<=16'd1061;
      8112:data<=16'd1099;
      8113:data<=16'd825;
      8114:data<=16'd1395;
      8115:data<=16'd1155;
      8116:data<=16'd1260;
      8117:data<=16'd1670;
      8118:data<=16'd1171;
      8119:data<=16'd1325;
      8120:data<=16'd1080;
      8121:data<=16'd1500;
      8122:data<=16'd2490;
      8123:data<=16'd1876;
      8124:data<=16'd7896;
      8125:data<=16'd18577;
      8126:data<=16'd19851;
      8127:data<=16'd17356;
      8128:data<=16'd18174;
      8129:data<=16'd16853;
      8130:data<=16'd15584;
      8131:data<=16'd15374;
      8132:data<=16'd13988;
      8133:data<=16'd13975;
      8134:data<=16'd13567;
      8135:data<=16'd12416;
      8136:data<=16'd12604;
      8137:data<=16'd11941;
      8138:data<=16'd11365;
      8139:data<=16'd11799;
      8140:data<=16'd11994;
      8141:data<=16'd12463;
      8142:data<=16'd11668;
      8143:data<=16'd10495;
      8144:data<=16'd10777;
      8145:data<=16'd10069;
      8146:data<=16'd9212;
      8147:data<=16'd9354;
      8148:data<=16'd8663;
      8149:data<=16'd7994;
      8150:data<=16'd7830;
      8151:data<=16'd7511;
      8152:data<=16'd7054;
      8153:data<=16'd6728;
      8154:data<=16'd6743;
      8155:data<=16'd5614;
      8156:data<=16'd5168;
      8157:data<=16'd7000;
      8158:data<=16'd6980;
      8159:data<=16'd6431;
      8160:data<=16'd7130;
      8161:data<=16'd5950;
      8162:data<=16'd5354;
      8163:data<=16'd4996;
      8164:data<=16'd3967;
      8165:data<=16'd5647;
      8166:data<=16'd1718;
      8167:data<=-16'd8531;
      8168:data<=-16'd10571;
      8169:data<=-16'd7746;
      8170:data<=-16'd8411;
      8171:data<=-16'd8520;
      8172:data<=-16'd8307;
      8173:data<=-16'd7764;
      8174:data<=-16'd6106;
      8175:data<=-16'd6670;
      8176:data<=-16'd7051;
      8177:data<=-16'd6155;
      8178:data<=-16'd6434;
      8179:data<=-16'd6446;
      8180:data<=-16'd6361;
      8181:data<=-16'd6088;
      8182:data<=-16'd5278;
      8183:data<=-16'd5779;
      8184:data<=-16'd5832;
      8185:data<=-16'd5350;
      8186:data<=-16'd5736;
      8187:data<=-16'd5024;
      8188:data<=-16'd4538;
      8189:data<=-16'd4695;
      8190:data<=-16'd3465;
      8191:data<=-16'd2830;
      8192:data<=-16'd2968;
      8193:data<=-16'd2534;
      8194:data<=-16'd2041;
      8195:data<=-16'd1644;
      8196:data<=-16'd2114;
      8197:data<=-16'd2111;
      8198:data<=-16'd1234;
      8199:data<=-16'd1642;
      8200:data<=-16'd1612;
      8201:data<=-16'd1347;
      8202:data<=-16'd1883;
      8203:data<=-16'd1310;
      8204:data<=-16'd1829;
      8205:data<=-16'd2070;
      8206:data<=-16'd437;
      8207:data<=-16'd951;
      8208:data<=16'd3052;
      8209:data<=16'd12515;
      8210:data<=16'd14108;
      8211:data<=16'd11561;
      8212:data<=16'd12675;
      8213:data<=16'd12169;
      8214:data<=16'd11075;
      8215:data<=16'd10874;
      8216:data<=16'd9538;
      8217:data<=16'd9838;
      8218:data<=16'd10014;
      8219:data<=16'd8270;
      8220:data<=16'd7679;
      8221:data<=16'd7694;
      8222:data<=16'd7376;
      8223:data<=16'd7275;
      8224:data<=16'd8129;
      8225:data<=16'd9973;
      8226:data<=16'd9962;
      8227:data<=16'd8795;
      8228:data<=16'd8563;
      8229:data<=16'd7774;
      8230:data<=16'd7345;
      8231:data<=16'd7658;
      8232:data<=16'd7235;
      8233:data<=16'd6748;
      8234:data<=16'd6099;
      8235:data<=16'd5706;
      8236:data<=16'd5659;
      8237:data<=16'd4983;
      8238:data<=16'd4664;
      8239:data<=16'd3877;
      8240:data<=16'd3374;
      8241:data<=16'd4974;
      8242:data<=16'd5248;
      8243:data<=16'd4526;
      8244:data<=16'd4488;
      8245:data<=16'd3607;
      8246:data<=16'd4108;
      8247:data<=16'd3794;
      8248:data<=16'd1980;
      8249:data<=16'd3559;
      8250:data<=16'd271;
      8251:data<=-16'd9652;
      8252:data<=-16'd12354;
      8253:data<=-16'd10481;
      8254:data<=-16'd11415;
      8255:data<=-16'd11089;
      8256:data<=-16'd9990;
      8257:data<=-16'd9041;
      8258:data<=-16'd7717;
      8259:data<=-16'd7915;
      8260:data<=-16'd7562;
      8261:data<=-16'd6492;
      8262:data<=-16'd6545;
      8263:data<=-16'd6731;
      8264:data<=-16'd7110;
      8265:data<=-16'd6711;
      8266:data<=-16'd5786;
      8267:data<=-16'd6096;
      8268:data<=-16'd5908;
      8269:data<=-16'd5421;
      8270:data<=-16'd5557;
      8271:data<=-16'd5554;
      8272:data<=-16'd5934;
      8273:data<=-16'd5071;
      8274:data<=-16'd3883;
      8275:data<=-16'd5009;
      8276:data<=-16'd5564;
      8277:data<=-16'd5286;
      8278:data<=-16'd5209;
      8279:data<=-16'd4062;
      8280:data<=-16'd4117;
      8281:data<=-16'd4757;
      8282:data<=-16'd4393;
      8283:data<=-16'd4825;
      8284:data<=-16'd4460;
      8285:data<=-16'd4012;
      8286:data<=-16'd4805;
      8287:data<=-16'd4558;
      8288:data<=-16'd5095;
      8289:data<=-16'd4999;
      8290:data<=-16'd3018;
      8291:data<=-16'd3483;
      8292:data<=16'd155;
      8293:data<=16'd9641;
      8294:data<=16'd11988;
      8295:data<=16'd9254;
      8296:data<=16'd9777;
      8297:data<=16'd9941;
      8298:data<=16'd9268;
      8299:data<=16'd8866;
      8300:data<=16'd7471;
      8301:data<=16'd7141;
      8302:data<=16'd7101;
      8303:data<=16'd6090;
      8304:data<=16'd5818;
      8305:data<=16'd5535;
      8306:data<=16'd4760;
      8307:data<=16'd4373;
      8308:data<=16'd4111;
      8309:data<=16'd3701;
      8310:data<=16'd2984;
      8311:data<=16'd2385;
      8312:data<=16'd2144;
      8313:data<=16'd2032;
      8314:data<=16'd2087;
      8315:data<=16'd1756;
      8316:data<=16'd1606;
      8317:data<=16'd1753;
      8318:data<=16'd931;
      8319:data<=16'd268;
      8320:data<=16'd20;
      8321:data<=-16'd155;
      8322:data<=16'd414;
      8323:data<=-16'd798;
      8324:data<=-16'd2319;
      8325:data<=-16'd720;
      8326:data<=-16'd109;
      8327:data<=-16'd822;
      8328:data<=-16'd470;
      8329:data<=-16'd1133;
      8330:data<=-16'd967;
      8331:data<=-16'd701;
      8332:data<=-16'd1830;
      8333:data<=-16'd614;
      8334:data<=-16'd3892;
      8335:data<=-16'd13822;
      8336:data<=-16'd16738;
      8337:data<=-16'd14045;
      8338:data<=-16'd14337;
      8339:data<=-16'd14280;
      8340:data<=-16'd14428;
      8341:data<=-16'd15571;
      8342:data<=-16'd14716;
      8343:data<=-16'd14384;
      8344:data<=-16'd14519;
      8345:data<=-16'd13311;
      8346:data<=-16'd12483;
      8347:data<=-16'd11846;
      8348:data<=-16'd11626;
      8349:data<=-16'd11972;
      8350:data<=-16'd11447;
      8351:data<=-16'd10804;
      8352:data<=-16'd10437;
      8353:data<=-16'd10138;
      8354:data<=-16'd9906;
      8355:data<=-16'd9080;
      8356:data<=-16'd8522;
      8357:data<=-16'd8792;
      8358:data<=-16'd9738;
      8359:data<=-16'd10678;
      8360:data<=-16'd10119;
      8361:data<=-16'd9673;
      8362:data<=-16'd9624;
      8363:data<=-16'd8464;
      8364:data<=-16'd8307;
      8365:data<=-16'd8341;
      8366:data<=-16'd7356;
      8367:data<=-16'd7482;
      8368:data<=-16'd7430;
      8369:data<=-16'd7215;
      8370:data<=-16'd7163;
      8371:data<=-16'd6023;
      8372:data<=-16'd6440;
      8373:data<=-16'd6583;
      8374:data<=-16'd6570;
      8375:data<=-16'd10231;
      8376:data<=-16'd7283;
      8377:data<=16'd3145;
      8378:data<=16'd5538;
      8379:data<=16'd3468;
      8380:data<=16'd4849;
      8381:data<=16'd4898;
      8382:data<=16'd4457;
      8383:data<=16'd4299;
      8384:data<=16'd3163;
      8385:data<=16'd3574;
      8386:data<=16'd3738;
      8387:data<=16'd2889;
      8388:data<=16'd2886;
      8389:data<=16'd2731;
      8390:data<=16'd2181;
      8391:data<=16'd699;
      8392:data<=-16'd587;
      8393:data<=-16'd112;
      8394:data<=-16'd194;
      8395:data<=-16'd373;
      8396:data<=-16'd180;
      8397:data<=-16'd860;
      8398:data<=-16'd437;
      8399:data<=-16'd115;
      8400:data<=-16'd740;
      8401:data<=-16'd253;
      8402:data<=-16'd402;
      8403:data<=-16'd623;
      8404:data<=-16'd208;
      8405:data<=-16'd826;
      8406:data<=-16'd508;
      8407:data<=-16'd845;
      8408:data<=-16'd2911;
      8409:data<=-16'd2914;
      8410:data<=-16'd2731;
      8411:data<=-16'd3063;
      8412:data<=-16'd2362;
      8413:data<=-16'd2337;
      8414:data<=-16'd1489;
      8415:data<=-16'd1613;
      8416:data<=-16'd3347;
      8417:data<=-16'd1721;
      8418:data<=-16'd4041;
      8419:data<=-16'd13277;
      8420:data<=-16'd16498;
      8421:data<=-16'd14219;
      8422:data<=-16'd14163;
      8423:data<=-16'd14110;
      8424:data<=-16'd13641;
      8425:data<=-16'd13236;
      8426:data<=-16'd12138;
      8427:data<=-16'd11749;
      8428:data<=-16'd11089;
      8429:data<=-16'd9809;
      8430:data<=-16'd9095;
      8431:data<=-16'd8530;
      8432:data<=-16'd8291;
      8433:data<=-16'd7947;
      8434:data<=-16'd7339;
      8435:data<=-16'd7294;
      8436:data<=-16'd6974;
      8437:data<=-16'd6300;
      8438:data<=-16'd5557;
      8439:data<=-16'd4722;
      8440:data<=-16'd5395;
      8441:data<=-16'd6927;
      8442:data<=-16'd6915;
      8443:data<=-16'd5984;
      8444:data<=-16'd5893;
      8445:data<=-16'd6349;
      8446:data<=-16'd5802;
      8447:data<=-16'd4808;
      8448:data<=-16'd4576;
      8449:data<=-16'd3947;
      8450:data<=-16'd3309;
      8451:data<=-16'd3606;
      8452:data<=-16'd3401;
      8453:data<=-16'd3043;
      8454:data<=-16'd3112;
      8455:data<=-16'd2817;
      8456:data<=-16'd2682;
      8457:data<=-16'd2575;
      8458:data<=-16'd3369;
      8459:data<=-16'd5016;
      8460:data<=-16'd1442;
      8461:data<=16'd7133;
      8462:data<=16'd11048;
      8463:data<=16'd9652;
      8464:data<=16'd9380;
      8465:data<=16'd9871;
      8466:data<=16'd9520;
      8467:data<=16'd9497;
      8468:data<=16'd9097;
      8469:data<=16'd8345;
      8470:data<=16'd8082;
      8471:data<=16'd7332;
      8472:data<=16'd6956;
      8473:data<=16'd7497;
      8474:data<=16'd6134;
      8475:data<=16'd3388;
      8476:data<=16'd2510;
      8477:data<=16'd2813;
      8478:data<=16'd2643;
      8479:data<=16'd2173;
      8480:data<=16'd1644;
      8481:data<=16'd1566;
      8482:data<=16'd1842;
      8483:data<=16'd1792;
      8484:data<=16'd1709;
      8485:data<=16'd1662;
      8486:data<=16'd1600;
      8487:data<=16'd1789;
      8488:data<=16'd1630;
      8489:data<=16'd1478;
      8490:data<=16'd1870;
      8491:data<=16'd1115;
      8492:data<=-16'd346;
      8493:data<=-16'd488;
      8494:data<=-16'd320;
      8495:data<=-16'd170;
      8496:data<=16'd247;
      8497:data<=-16'd58;
      8498:data<=-16'd150;
      8499:data<=-16'd390;
      8500:data<=-16'd701;
      8501:data<=16'd945;
      8502:data<=-16'd1198;
      8503:data<=-16'd9464;
      8504:data<=-16'd13600;
      8505:data<=-16'd12076;
      8506:data<=-16'd11418;
      8507:data<=-16'd11532;
      8508:data<=-16'd12132;
      8509:data<=-16'd12464;
      8510:data<=-16'd11332;
      8511:data<=-16'd11182;
      8512:data<=-16'd10701;
      8513:data<=-16'd9051;
      8514:data<=-16'd8815;
      8515:data<=-16'd8291;
      8516:data<=-16'd7301;
      8517:data<=-16'd7465;
      8518:data<=-16'd7269;
      8519:data<=-16'd6672;
      8520:data<=-16'd5729;
      8521:data<=-16'd4825;
      8522:data<=-16'd4948;
      8523:data<=-16'd4578;
      8524:data<=-16'd4582;
      8525:data<=-16'd4855;
      8526:data<=-16'd3251;
      8527:data<=-16'd2746;
      8528:data<=-16'd3354;
      8529:data<=-16'd2623;
      8530:data<=-16'd2585;
      8531:data<=-16'd2240;
      8532:data<=-16'd1048;
      8533:data<=-16'd1095;
      8534:data<=-16'd901;
      8535:data<=-16'd760;
      8536:data<=-16'd1128;
      8537:data<=-16'd585;
      8538:data<=-16'd111;
      8539:data<=16'd519;
      8540:data<=16'd567;
      8541:data<=-16'd558;
      8542:data<=-16'd789;
      8543:data<=-16'd1577;
      8544:data<=16'd593;
      8545:data<=16'd9307;
      8546:data<=16'd14105;
      8547:data<=16'd12372;
      8548:data<=16'd12355;
      8549:data<=16'd12401;
      8550:data<=16'd11373;
      8551:data<=16'd11696;
      8552:data<=16'd11292;
      8553:data<=16'd10924;
      8554:data<=16'd10894;
      8555:data<=16'd9781;
      8556:data<=16'd9652;
      8557:data<=16'd9461;
      8558:data<=16'd7733;
      8559:data<=16'd7001;
      8560:data<=16'd7084;
      8561:data<=16'd6739;
      8562:data<=16'd6743;
      8563:data<=16'd6780;
      8564:data<=16'd6184;
      8565:data<=16'd5744;
      8566:data<=16'd6053;
      8567:data<=16'd6108;
      8568:data<=16'd5638;
      8569:data<=16'd5506;
      8570:data<=16'd5330;
      8571:data<=16'd5140;
      8572:data<=16'd5244;
      8573:data<=16'd5072;
      8574:data<=16'd5045;
      8575:data<=16'd4999;
      8576:data<=16'd4739;
      8577:data<=16'd5157;
      8578:data<=16'd5366;
      8579:data<=16'd5093;
      8580:data<=16'd5030;
      8581:data<=16'd4679;
      8582:data<=16'd5046;
      8583:data<=16'd5438;
      8584:data<=16'd4589;
      8585:data<=16'd5077;
      8586:data<=16'd3929;
      8587:data<=-16'd2701;
      8588:data<=-16'd7236;
      8589:data<=-16'd6290;
      8590:data<=-16'd5841;
      8591:data<=-16'd5274;
      8592:data<=-16'd3016;
      8593:data<=-16'd2543;
      8594:data<=-16'd2964;
      8595:data<=-16'd2452;
      8596:data<=-16'd2208;
      8597:data<=-16'd1926;
      8598:data<=-16'd1656;
      8599:data<=-16'd1374;
      8600:data<=-16'd308;
      8601:data<=-16'd6;
      8602:data<=-16'd432;
      8603:data<=-16'd270;
      8604:data<=-16'd305;
      8605:data<=16'd187;
      8606:data<=16'd974;
      8607:data<=16'd646;
      8608:data<=16'd1387;
      8609:data<=16'd3008;
      8610:data<=16'd3209;
      8611:data<=16'd3341;
      8612:data<=16'd3333;
      8613:data<=16'd2482;
      8614:data<=16'd2437;
      8615:data<=16'd2907;
      8616:data<=16'd3095;
      8617:data<=16'd3154;
      8618:data<=16'd3052;
      8619:data<=16'd3206;
      8620:data<=16'd3066;
      8621:data<=16'd2707;
      8622:data<=16'd2836;
      8623:data<=16'd2423;
      8624:data<=16'd2326;
      8625:data<=16'd4012;
      8626:data<=16'd5256;
      8627:data<=16'd4560;
      8628:data<=16'd5495;
      8629:data<=16'd11351;
      8630:data<=16'd16625;
      8631:data<=16'd15638;
      8632:data<=16'd13797;
      8633:data<=16'd14193;
      8634:data<=16'd13544;
      8635:data<=16'd13399;
      8636:data<=16'd13532;
      8637:data<=16'd11953;
      8638:data<=16'd11646;
      8639:data<=16'd11841;
      8640:data<=16'd10545;
      8641:data<=16'd10399;
      8642:data<=16'd11342;
      8643:data<=16'd11747;
      8644:data<=16'd11617;
      8645:data<=16'd10969;
      8646:data<=16'd10457;
      8647:data<=16'd9873;
      8648:data<=16'd9260;
      8649:data<=16'd9291;
      8650:data<=16'd8812;
      8651:data<=16'd7876;
      8652:data<=16'd7479;
      8653:data<=16'd7090;
      8654:data<=16'd6953;
      8655:data<=16'd7307;
      8656:data<=16'd7169;
      8657:data<=16'd6472;
      8658:data<=16'd6810;
      8659:data<=16'd8188;
      8660:data<=16'd8120;
      8661:data<=16'd7228;
      8662:data<=16'd7198;
      8663:data<=16'd6734;
      8664:data<=16'd6522;
      8665:data<=16'd6707;
      8666:data<=16'd5891;
      8667:data<=16'd5683;
      8668:data<=16'd5468;
      8669:data<=16'd4708;
      8670:data<=16'd3952;
      8671:data<=-16'd1010;
      8672:data<=-16'd7074;
      8673:data<=-16'd7037;
      8674:data<=-16'd5404;
      8675:data<=-16'd5093;
      8676:data<=-16'd3695;
      8677:data<=-16'd3356;
      8678:data<=-16'd3783;
      8679:data<=-16'd3510;
      8680:data<=-16'd3485;
      8681:data<=-16'd2964;
      8682:data<=-16'd2552;
      8683:data<=-16'd2529;
      8684:data<=-16'd2127;
      8685:data<=-16'd2303;
      8686:data<=-16'd2428;
      8687:data<=-16'd2473;
      8688:data<=-16'd2684;
      8689:data<=-16'd1917;
      8690:data<=-16'd1879;
      8691:data<=-16'd1745;
      8692:data<=16'd346;
      8693:data<=16'd893;
      8694:data<=16'd15;
      8695:data<=16'd191;
      8696:data<=16'd140;
      8697:data<=-16'd42;
      8698:data<=-16'd255;
      8699:data<=-16'd599;
      8700:data<=-16'd352;
      8701:data<=-16'd514;
      8702:data<=-16'd397;
      8703:data<=-16'd105;
      8704:data<=-16'd898;
      8705:data<=-16'd696;
      8706:data<=-16'd314;
      8707:data<=-16'd740;
      8708:data<=16'd412;
      8709:data<=16'd1497;
      8710:data<=16'd1697;
      8711:data<=16'd1606;
      8712:data<=16'd1127;
      8713:data<=16'd5348;
      8714:data<=16'd11899;
      8715:data<=16'd12222;
      8716:data<=16'd10596;
      8717:data<=16'd10937;
      8718:data<=16'd9858;
      8719:data<=16'd9072;
      8720:data<=16'd8957;
      8721:data<=16'd8263;
      8722:data<=16'd8304;
      8723:data<=16'd7382;
      8724:data<=16'd6379;
      8725:data<=16'd7460;
      8726:data<=16'd7799;
      8727:data<=16'd7265;
      8728:data<=16'd7150;
      8729:data<=16'd6508;
      8730:data<=16'd6166;
      8731:data<=16'd5902;
      8732:data<=16'd5125;
      8733:data<=16'd4719;
      8734:data<=16'd4181;
      8735:data<=16'd3855;
      8736:data<=16'd3815;
      8737:data<=16'd2993;
      8738:data<=16'd2623;
      8739:data<=16'd2802;
      8740:data<=16'd2382;
      8741:data<=16'd2281;
      8742:data<=16'd2816;
      8743:data<=16'd3410;
      8744:data<=16'd3475;
      8745:data<=16'd3001;
      8746:data<=16'd2874;
      8747:data<=16'd2634;
      8748:data<=16'd2356;
      8749:data<=16'd2457;
      8750:data<=16'd2035;
      8751:data<=16'd1859;
      8752:data<=16'd1691;
      8753:data<=16'd1321;
      8754:data<=16'd1692;
      8755:data<=-16'd1930;
      8756:data<=-16'd9135;
      8757:data<=-16'd10941;
      8758:data<=-16'd8890;
      8759:data<=-16'd8390;
      8760:data<=-16'd7820;
      8761:data<=-16'd7577;
      8762:data<=-16'd7680;
      8763:data<=-16'd7282;
      8764:data<=-16'd7532;
      8765:data<=-16'd6954;
      8766:data<=-16'd6264;
      8767:data<=-16'd6736;
      8768:data<=-16'd6120;
      8769:data<=-16'd5641;
      8770:data<=-16'd6049;
      8771:data<=-16'd5937;
      8772:data<=-16'd6024;
      8773:data<=-16'd5477;
      8774:data<=-16'd4896;
      8775:data<=-16'd5007;
      8776:data<=-16'd3630;
      8777:data<=-16'd2616;
      8778:data<=-16'd2802;
      8779:data<=-16'd2355;
      8780:data<=-16'd2667;
      8781:data<=-16'd3075;
      8782:data<=-16'd2987;
      8783:data<=-16'd3157;
      8784:data<=-16'd2508;
      8785:data<=-16'd2796;
      8786:data<=-16'd3432;
      8787:data<=-16'd2544;
      8788:data<=-16'd2890;
      8789:data<=-16'd3254;
      8790:data<=-16'd2757;
      8791:data<=-16'd2719;
      8792:data<=-16'd1093;
      8793:data<=-16'd626;
      8794:data<=-16'd1519;
      8795:data<=-16'd1007;
      8796:data<=-16'd2338;
      8797:data<=16'd503;
      8798:data<=16'd9169;
      8799:data<=16'd10345;
      8800:data<=16'd7410;
      8801:data<=16'd8322;
      8802:data<=16'd7799;
      8803:data<=16'd7307;
      8804:data<=16'd7612;
      8805:data<=16'd6235;
      8806:data<=16'd6367;
      8807:data<=16'd5900;
      8808:data<=16'd5033;
      8809:data<=16'd6907;
      8810:data<=16'd6940;
      8811:data<=16'd5783;
      8812:data<=16'd6169;
      8813:data<=16'd5457;
      8814:data<=16'd4610;
      8815:data<=16'd4002;
      8816:data<=16'd3381;
      8817:data<=16'd3641;
      8818:data<=16'd2805;
      8819:data<=16'd2185;
      8820:data<=16'd2458;
      8821:data<=16'd1629;
      8822:data<=16'd1801;
      8823:data<=16'd2153;
      8824:data<=16'd1236;
      8825:data<=16'd1677;
      8826:data<=16'd2632;
      8827:data<=16'd2986;
      8828:data<=16'd2808;
      8829:data<=16'd1903;
      8830:data<=16'd1906;
      8831:data<=16'd1829;
      8832:data<=16'd1327;
      8833:data<=16'd1145;
      8834:data<=16'd36;
      8835:data<=16'd497;
      8836:data<=16'd1265;
      8837:data<=-16'd99;
      8838:data<=16'd713;
      8839:data<=-16'd1783;
      8840:data<=-16'd10199;
      8841:data<=-16'd12175;
      8842:data<=-16'd9917;
      8843:data<=-16'd11351;
      8844:data<=-16'd11294;
      8845:data<=-16'd10085;
      8846:data<=-16'd10305;
      8847:data<=-16'd9979;
      8848:data<=-16'd10067;
      8849:data<=-16'd9679;
      8850:data<=-16'd9034;
      8851:data<=-16'd9321;
      8852:data<=-16'd8502;
      8853:data<=-16'd8390;
      8854:data<=-16'd9063;
      8855:data<=-16'd8263;
      8856:data<=-16'd8299;
      8857:data<=-16'd8302;
      8858:data<=-16'd7712;
      8859:data<=-16'd8790;
      8860:data<=-16'd8931;
      8861:data<=-16'd8222;
      8862:data<=-16'd8728;
      8863:data<=-16'd8429;
      8864:data<=-16'd7909;
      8865:data<=-16'd8146;
      8866:data<=-16'd8384;
      8867:data<=-16'd8539;
      8868:data<=-16'd7859;
      8869:data<=-16'd7673;
      8870:data<=-16'd8058;
      8871:data<=-16'd7224;
      8872:data<=-16'd7006;
      8873:data<=-16'd7275;
      8874:data<=-16'd6858;
      8875:data<=-16'd7212;
      8876:data<=-16'd7971;
      8877:data<=-16'd8997;
      8878:data<=-16'd8937;
      8879:data<=-16'd7705;
      8880:data<=-16'd8745;
      8881:data<=-16'd6187;
      8882:data<=16'd2238;
      8883:data<=16'd4673;
      8884:data<=16'd2275;
      8885:data<=16'd3143;
      8886:data<=16'd3156;
      8887:data<=16'd2197;
      8888:data<=16'd2863;
      8889:data<=16'd2382;
      8890:data<=16'd1847;
      8891:data<=16'd1824;
      8892:data<=16'd667;
      8893:data<=-16'd458;
      8894:data<=-16'd1174;
      8895:data<=-16'd1342;
      8896:data<=-16'd1158;
      8897:data<=-16'd1450;
      8898:data<=-16'd1374;
      8899:data<=-16'd1283;
      8900:data<=-16'd1387;
      8901:data<=-16'd1395;
      8902:data<=-16'd2296;
      8903:data<=-16'd2510;
      8904:data<=-16'd1776;
      8905:data<=-16'd2438;
      8906:data<=-16'd2854;
      8907:data<=-16'd1879;
      8908:data<=-16'd1801;
      8909:data<=-16'd3151;
      8910:data<=-16'd4099;
      8911:data<=-16'd3577;
      8912:data<=-16'd3307;
      8913:data<=-16'd3566;
      8914:data<=-16'd3101;
      8915:data<=-16'd3330;
      8916:data<=-16'd3629;
      8917:data<=-16'd3359;
      8918:data<=-16'd3958;
      8919:data<=-16'd3466;
      8920:data<=-16'd2913;
      8921:data<=-16'd3275;
      8922:data<=-16'd1809;
      8923:data<=-16'd4517;
      8924:data<=-16'd12319;
      8925:data<=-16'd14854;
      8926:data<=-16'd14017;
      8927:data<=-16'd14748;
      8928:data<=-16'd14204;
      8929:data<=-16'd13814;
      8930:data<=-16'd13667;
      8931:data<=-16'd12610;
      8932:data<=-16'd12524;
      8933:data<=-16'd11781;
      8934:data<=-16'd10803;
      8935:data<=-16'd10813;
      8936:data<=-16'd9873;
      8937:data<=-16'd9320;
      8938:data<=-16'd9157;
      8939:data<=-16'd8654;
      8940:data<=-16'd8830;
      8941:data<=-16'd7652;
      8942:data<=-16'd6960;
      8943:data<=-16'd8508;
      8944:data<=-16'd8402;
      8945:data<=-16'd7783;
      8946:data<=-16'd7877;
      8947:data<=-16'd7283;
      8948:data<=-16'd7591;
      8949:data<=-16'd7297;
      8950:data<=-16'd6211;
      8951:data<=-16'd6394;
      8952:data<=-16'd5990;
      8953:data<=-16'd5802;
      8954:data<=-16'd6008;
      8955:data<=-16'd5150;
      8956:data<=-16'd5322;
      8957:data<=-16'd5060;
      8958:data<=-16'd4085;
      8959:data<=-16'd4854;
      8960:data<=-16'd5456;
      8961:data<=-16'd6203;
      8962:data<=-16'd5930;
      8963:data<=-16'd4150;
      8964:data<=-16'd5554;
      8965:data<=-16'd3198;
      8966:data<=16'd5627;
      8967:data<=16'd8116;
      8968:data<=16'd6294;
      8969:data<=16'd6777;
      8970:data<=16'd5547;
      8971:data<=16'd5335;
      8972:data<=16'd6490;
      8973:data<=16'd5400;
      8974:data<=16'd5439;
      8975:data<=16'd5545;
      8976:data<=16'd3938;
      8977:data<=16'd3015;
      8978:data<=16'd2261;
      8979:data<=16'd2761;
      8980:data<=16'd3821;
      8981:data<=16'd3133;
      8982:data<=16'd3063;
      8983:data<=16'd2948;
      8984:data<=16'd2235;
      8985:data<=16'd2875;
      8986:data<=16'd2319;
      8987:data<=16'd1303;
      8988:data<=16'd2232;
      8989:data<=16'd2440;
      8990:data<=16'd2379;
      8991:data<=16'd3077;
      8992:data<=16'd2331;
      8993:data<=16'd1048;
      8994:data<=16'd899;
      8995:data<=16'd1080;
      8996:data<=16'd878;
      8997:data<=16'd808;
      8998:data<=16'd1087;
      8999:data<=16'd1063;
      9000:data<=16'd1227;
      9001:data<=16'd1286;
      9002:data<=16'd1010;
      9003:data<=16'd1859;
      9004:data<=16'd1814;
      9005:data<=16'd1166;
      9006:data<=16'd2585;
      9007:data<=-16'd138;
      9008:data<=-16'd7547;
      9009:data<=-16'd10063;
      9010:data<=-16'd9368;
      9011:data<=-16'd10323;
      9012:data<=-16'd9970;
      9013:data<=-16'd8948;
      9014:data<=-16'd8746;
      9015:data<=-16'd7841;
      9016:data<=-16'd6804;
      9017:data<=-16'd6273;
      9018:data<=-16'd6156;
      9019:data<=-16'd6096;
      9020:data<=-16'd5636;
      9021:data<=-16'd5203;
      9022:data<=-16'd4619;
      9023:data<=-16'd4334;
      9024:data<=-16'd4356;
      9025:data<=-16'd3852;
      9026:data<=-16'd4219;
      9027:data<=-16'd4790;
      9028:data<=-16'd4129;
      9029:data<=-16'd4091;
      9030:data<=-16'd4120;
      9031:data<=-16'd3471;
      9032:data<=-16'd3169;
      9033:data<=-16'd2555;
      9034:data<=-16'd2634;
      9035:data<=-16'd2914;
      9036:data<=-16'd2024;
      9037:data<=-16'd2140;
      9038:data<=-16'd1756;
      9039:data<=-16'd367;
      9040:data<=-16'd745;
      9041:data<=-16'd459;
      9042:data<=-16'd414;
      9043:data<=-16'd2218;
      9044:data<=-16'd2187;
      9045:data<=-16'd2221;
      9046:data<=-16'd1976;
      9047:data<=-16'd82;
      9048:data<=-16'd1447;
      9049:data<=16'd467;
      9050:data<=16'd8660;
      9051:data<=16'd11042;
      9052:data<=16'd9999;
      9053:data<=16'd11217;
      9054:data<=16'd9844;
      9055:data<=16'd9242;
      9056:data<=16'd10336;
      9057:data<=16'd9289;
      9058:data<=16'd9163;
      9059:data<=16'd8743;
      9060:data<=16'd7206;
      9061:data<=16'd7376;
      9062:data<=16'd6858;
      9063:data<=16'd6404;
      9064:data<=16'd6774;
      9065:data<=16'd5739;
      9066:data<=16'd6040;
      9067:data<=16'd6724;
      9068:data<=16'd5611;
      9069:data<=16'd5530;
      9070:data<=16'd5218;
      9071:data<=16'd4781;
      9072:data<=16'd6352;
      9073:data<=16'd6646;
      9074:data<=16'd5724;
      9075:data<=16'd5826;
      9076:data<=16'd5294;
      9077:data<=16'd4228;
      9078:data<=16'd3894;
      9079:data<=16'd4237;
      9080:data<=16'd4505;
      9081:data<=16'd4049;
      9082:data<=16'd3841;
      9083:data<=16'd4067;
      9084:data<=16'd4206;
      9085:data<=16'd4053;
      9086:data<=16'd3491;
      9087:data<=16'd3711;
      9088:data<=16'd3638;
      9089:data<=16'd3342;
      9090:data<=16'd5002;
      9091:data<=16'd2649;
      9092:data<=-16'd5156;
      9093:data<=-16'd8396;
      9094:data<=-16'd7382;
      9095:data<=-16'd7721;
      9096:data<=-16'd7655;
      9097:data<=-16'd7536;
      9098:data<=-16'd7188;
      9099:data<=-16'd5523;
      9100:data<=-16'd5356;
      9101:data<=-16'd5641;
      9102:data<=-16'd5112;
      9103:data<=-16'd5172;
      9104:data<=-16'd4282;
      9105:data<=-16'd3469;
      9106:data<=-16'd3892;
      9107:data<=-16'd3225;
      9108:data<=-16'd2787;
      9109:data<=-16'd2839;
      9110:data<=-16'd1483;
      9111:data<=-16'd1010;
      9112:data<=-16'd1544;
      9113:data<=-16'd930;
      9114:data<=-16'd387;
      9115:data<=-16'd517;
      9116:data<=-16'd770;
      9117:data<=-16'd816;
      9118:data<=16'd50;
      9119:data<=16'd625;
      9120:data<=16'd244;
      9121:data<=16'd469;
      9122:data<=16'd995;
      9123:data<=16'd816;
      9124:data<=16'd534;
      9125:data<=16'd434;
      9126:data<=16'd1121;
      9127:data<=16'd3072;
      9128:data<=16'd4035;
      9129:data<=16'd3271;
      9130:data<=16'd3698;
      9131:data<=16'd4252;
      9132:data<=16'd2916;
      9133:data<=16'd5215;
      9134:data<=16'd12141;
      9135:data<=16'd15139;
      9136:data<=16'd13726;
      9137:data<=16'd13553;
      9138:data<=16'd13336;
      9139:data<=16'd12481;
      9140:data<=16'd12828;
      9141:data<=16'd12226;
      9142:data<=16'd11200;
      9143:data<=16'd12513;
      9144:data<=16'd13975;
      9145:data<=16'd13562;
      9146:data<=16'd12583;
      9147:data<=16'd12172;
      9148:data<=16'd12258;
      9149:data<=16'd11489;
      9150:data<=16'd10122;
      9151:data<=16'd10251;
      9152:data<=16'd10878;
      9153:data<=16'd10379;
      9154:data<=16'd9630;
      9155:data<=16'd8707;
      9156:data<=16'd8105;
      9157:data<=16'd8583;
      9158:data<=16'd8178;
      9159:data<=16'd7421;
      9160:data<=16'd8689;
      9161:data<=16'd9514;
      9162:data<=16'd8724;
      9163:data<=16'd8683;
      9164:data<=16'd8592;
      9165:data<=16'd8120;
      9166:data<=16'd8049;
      9167:data<=16'd7175;
      9168:data<=16'd6871;
      9169:data<=16'd7291;
      9170:data<=16'd6463;
      9171:data<=16'd6520;
      9172:data<=16'd6648;
      9173:data<=16'd5553;
      9174:data<=16'd6296;
      9175:data<=16'd4193;
      9176:data<=-16'd2331;
      9177:data<=-16'd4061;
      9178:data<=-16'd3004;
      9179:data<=-16'd4361;
      9180:data<=-16'd3644;
      9181:data<=-16'd2572;
      9182:data<=-16'd3791;
      9183:data<=-16'd3782;
      9184:data<=-16'd3266;
      9185:data<=-16'd3377;
      9186:data<=-16'd3674;
      9187:data<=-16'd3953;
      9188:data<=-16'd2716;
      9189:data<=-16'd2258;
      9190:data<=-16'd3137;
      9191:data<=-16'd2748;
      9192:data<=-16'd3018;
      9193:data<=-16'd2616;
      9194:data<=-16'd200;
      9195:data<=-16'd133;
      9196:data<=-16'd472;
      9197:data<=16'd328;
      9198:data<=-16'd1061;
      9199:data<=-16'd1697;
      9200:data<=-16'd649;
      9201:data<=-16'd696;
      9202:data<=-16'd332;
      9203:data<=-16'd118;
      9204:data<=-16'd708;
      9205:data<=-16'd459;
      9206:data<=-16'd382;
      9207:data<=-16'd246;
      9208:data<=16'd161;
      9209:data<=-16'd61;
      9210:data<=16'd1022;
      9211:data<=16'd2831;
      9212:data<=16'd2842;
      9213:data<=16'd1900;
      9214:data<=16'd1489;
      9215:data<=16'd1604;
      9216:data<=16'd1207;
      9217:data<=16'd2682;
      9218:data<=16'd8469;
      9219:data<=16'd12392;
      9220:data<=16'd11952;
      9221:data<=16'd12134;
      9222:data<=16'd11585;
      9223:data<=16'd9858;
      9224:data<=16'd9955;
      9225:data<=16'd9547;
      9226:data<=16'd9412;
      9227:data<=16'd11092;
      9228:data<=16'd10721;
      9229:data<=16'd9136;
      9230:data<=16'd8498;
      9231:data<=16'd7714;
      9232:data<=16'd7670;
      9233:data<=16'd7614;
      9234:data<=16'd6962;
      9235:data<=16'd7342;
      9236:data<=16'd7279;
      9237:data<=16'd6399;
      9238:data<=16'd5850;
      9239:data<=16'd5060;
      9240:data<=16'd5148;
      9241:data<=16'd5457;
      9242:data<=16'd4587;
      9243:data<=16'd5159;
      9244:data<=16'd6420;
      9245:data<=16'd5633;
      9246:data<=16'd4899;
      9247:data<=16'd5312;
      9248:data<=16'd5501;
      9249:data<=16'd5247;
      9250:data<=16'd4510;
      9251:data<=16'd3660;
      9252:data<=16'd3069;
      9253:data<=16'd2566;
      9254:data<=16'd2449;
      9255:data<=16'd2387;
      9256:data<=16'd1770;
      9257:data<=16'd1454;
      9258:data<=16'd1677;
      9259:data<=-16'd247;
      9260:data<=-16'd5089;
      9261:data<=-16'd8085;
      9262:data<=-16'd7498;
      9263:data<=-16'd7313;
      9264:data<=-16'd7858;
      9265:data<=-16'd7489;
      9266:data<=-16'd7591;
      9267:data<=-16'd7694;
      9268:data<=-16'd6470;
      9269:data<=-16'd5495;
      9270:data<=-16'd6079;
      9271:data<=-16'd7206;
      9272:data<=-16'd6925;
      9273:data<=-16'd5356;
      9274:data<=-16'd4672;
      9275:data<=-16'd5204;
      9276:data<=-16'd5668;
      9277:data<=-16'd5319;
      9278:data<=-16'd4546;
      9279:data<=-16'd4695;
      9280:data<=-16'd5147;
      9281:data<=-16'd4300;
      9282:data<=-16'd3330;
      9283:data<=-16'd3325;
      9284:data<=-16'd3544;
      9285:data<=-16'd3827;
      9286:data<=-16'd3892;
      9287:data<=-16'd3524;
      9288:data<=-16'd3792;
      9289:data<=-16'd4391;
      9290:data<=-16'd3892;
      9291:data<=-16'd3553;
      9292:data<=-16'd4059;
      9293:data<=-16'd3046;
      9294:data<=-16'd1565;
      9295:data<=-16'd1938;
      9296:data<=-16'd1633;
      9297:data<=-16'd479;
      9298:data<=-16'd855;
      9299:data<=-16'd1286;
      9300:data<=-16'd1483;
      9301:data<=-16'd341;
      9302:data<=16'd4993;
      9303:data<=16'd9163;
      9304:data<=16'd8294;
      9305:data<=16'd7524;
      9306:data<=16'd7398;
      9307:data<=16'd6657;
      9308:data<=16'd7124;
      9309:data<=16'd6466;
      9310:data<=16'd5330;
      9311:data<=16'd7269;
      9312:data<=16'd8493;
      9313:data<=16'd6608;
      9314:data<=16'd5274;
      9315:data<=16'd5691;
      9316:data<=16'd6304;
      9317:data<=16'd6140;
      9318:data<=16'd5792;
      9319:data<=16'd5375;
      9320:data<=16'd3926;
      9321:data<=16'd3181;
      9322:data<=16'd3783;
      9323:data<=16'd3362;
      9324:data<=16'd2616;
      9325:data<=16'd2848;
      9326:data<=16'd3284;
      9327:data<=16'd3524;
      9328:data<=16'd3240;
      9329:data<=16'd3292;
      9330:data<=16'd3891;
      9331:data<=16'd3598;
      9332:data<=16'd2952;
      9333:data<=16'd2255;
      9334:data<=16'd1597;
      9335:data<=16'd1876;
      9336:data<=16'd1510;
      9337:data<=16'd246;
      9338:data<=-16'd399;
      9339:data<=-16'd517;
      9340:data<=16'd55;
      9341:data<=-16'd59;
      9342:data<=-16'd640;
      9343:data<=-16'd164;
      9344:data<=-16'd3107;
      9345:data<=-16'd8865;
      9346:data<=-16'd10748;
      9347:data<=-16'd10196;
      9348:data<=-16'd9388;
      9349:data<=-16'd8853;
      9350:data<=-16'd10349;
      9351:data<=-16'd9850;
      9352:data<=-16'd7727;
      9353:data<=-16'd8523;
      9354:data<=-16'd8778;
      9355:data<=-16'd8228;
      9356:data<=-16'd9233;
      9357:data<=-16'd8881;
      9358:data<=-16'd7976;
      9359:data<=-16'd7451;
      9360:data<=-16'd6194;
      9361:data<=-16'd6052;
      9362:data<=-16'd5768;
      9363:data<=-16'd4887;
      9364:data<=-16'd5824;
      9365:data<=-16'd6288;
      9366:data<=-16'd5621;
      9367:data<=-16'd5962;
      9368:data<=-16'd5855;
      9369:data<=-16'd5066;
      9370:data<=-16'd5230;
      9371:data<=-16'd5655;
      9372:data<=-16'd5238;
      9373:data<=-16'd4573;
      9374:data<=-16'd4687;
      9375:data<=-16'd5260;
      9376:data<=-16'd5583;
      9377:data<=-16'd5184;
      9378:data<=-16'd4514;
      9379:data<=-16'd4943;
      9380:data<=-16'd5090;
      9381:data<=-16'd4369;
      9382:data<=-16'd4532;
      9383:data<=-16'd3970;
      9384:data<=-16'd3786;
      9385:data<=-16'd5098;
      9386:data<=-16'd1378;
      9387:data<=16'd5198;
      9388:data<=16'd6335;
      9389:data<=16'd5447;
      9390:data<=16'd5280;
      9391:data<=16'd4267;
      9392:data<=16'd4814;
      9393:data<=16'd4801;
      9394:data<=16'd2261;
      9395:data<=16'd1074;
      9396:data<=16'd772;
      9397:data<=16'd258;
      9398:data<=16'd1133;
      9399:data<=16'd1263;
      9400:data<=-16'd58;
      9401:data<=-16'd73;
      9402:data<=16'd804;
      9403:data<=16'd658;
      9404:data<=-16'd132;
      9405:data<=-16'd511;
      9406:data<=-16'd397;
      9407:data<=-16'd303;
      9408:data<=-16'd476;
      9409:data<=-16'd755;
      9410:data<=-16'd1535;
      9411:data<=-16'd3116;
      9412:data<=-16'd3829;
      9413:data<=-16'd3459;
      9414:data<=-16'd4212;
      9415:data<=-16'd4748;
      9416:data<=-16'd3917;
      9417:data<=-16'd4217;
      9418:data<=-16'd4473;
      9419:data<=-16'd3871;
      9420:data<=-16'd4798;
      9421:data<=-16'd4911;
      9422:data<=-16'd3586;
      9423:data<=-16'd3988;
      9424:data<=-16'd4293;
      9425:data<=-16'd3635;
      9426:data<=-16'd3160;
      9427:data<=-16'd3231;
      9428:data<=-16'd8510;
      9429:data<=-16'd16507;
      9430:data<=-16'd17462;
      9431:data<=-16'd14566;
      9432:data<=-16'd14578;
      9433:data<=-16'd15086;
      9434:data<=-16'd15035;
      9435:data<=-16'd14575;
      9436:data<=-16'd13212;
      9437:data<=-16'd12745;
      9438:data<=-16'd12346;
      9439:data<=-16'd11354;
      9440:data<=-16'd11486;
      9441:data<=-16'd11747;
      9442:data<=-16'd11279;
      9443:data<=-16'd10715;
      9444:data<=-16'd10436;
      9445:data<=-16'd11115;
      9446:data<=-16'd11749;
      9447:data<=-16'd11452;
      9448:data<=-16'd10780;
      9449:data<=-16'd9770;
      9450:data<=-16'd9286;
      9451:data<=-16'd9544;
      9452:data<=-16'd9723;
      9453:data<=-16'd9750;
      9454:data<=-16'd8605;
      9455:data<=-16'd6884;
      9456:data<=-16'd6558;
      9457:data<=-16'd6664;
      9458:data<=-16'd6237;
      9459:data<=-16'd5868;
      9460:data<=-16'd6420;
      9461:data<=-16'd7714;
      9462:data<=-16'd8014;
      9463:data<=-16'd7793;
      9464:data<=-16'd7156;
      9465:data<=-16'd5726;
      9466:data<=-16'd5789;
      9467:data<=-16'd5190;
      9468:data<=-16'd3940;
      9469:data<=-16'd5839;
      9470:data<=-16'd3196;
      9471:data<=16'd5139;
      9472:data<=16'd7474;
      9473:data<=16'd6363;
      9474:data<=16'd6633;
      9475:data<=16'd5412;
      9476:data<=16'd5874;
      9477:data<=16'd6173;
      9478:data<=16'd3833;
      9479:data<=16'd3745;
      9480:data<=16'd3263;
      9481:data<=16'd2055;
      9482:data<=16'd3789;
      9483:data<=16'd4053;
      9484:data<=16'd3896;
      9485:data<=16'd5033;
      9486:data<=16'd3294;
      9487:data<=16'd2952;
      9488:data<=16'd5150;
      9489:data<=16'd4526;
      9490:data<=16'd3753;
      9491:data<=16'd3682;
      9492:data<=16'd2411;
      9493:data<=16'd2669;
      9494:data<=16'd2986;
      9495:data<=16'd1111;
      9496:data<=-16'd64;
      9497:data<=16'd208;
      9498:data<=16'd493;
      9499:data<=16'd905;
      9500:data<=16'd937;
      9501:data<=-16'd490;
      9502:data<=-16'd1412;
      9503:data<=16'd155;
      9504:data<=16'd1727;
      9505:data<=16'd1882;
      9506:data<=16'd1754;
      9507:data<=16'd1635;
      9508:data<=16'd1970;
      9509:data<=16'd1381;
      9510:data<=16'd358;
      9511:data<=16'd873;
      9512:data<=-16'd2957;
      9513:data<=-16'd10948;
      9514:data<=-16'd12684;
      9515:data<=-16'd10457;
      9516:data<=-16'd10470;
      9517:data<=-16'd9603;
      9518:data<=-16'd8925;
      9519:data<=-16'd9453;
      9520:data<=-16'd7946;
      9521:data<=-16'd6549;
      9522:data<=-16'd6730;
      9523:data<=-16'd6670;
      9524:data<=-16'd6525;
      9525:data<=-16'd5856;
      9526:data<=-16'd4833;
      9527:data<=-16'd5136;
      9528:data<=-16'd6623;
      9529:data<=-16'd7371;
      9530:data<=-16'd6144;
      9531:data<=-16'd4990;
      9532:data<=-16'd5253;
      9533:data<=-16'd4793;
      9534:data<=-16'd3770;
      9535:data<=-16'd3805;
      9536:data<=-16'd3889;
      9537:data<=-16'd2890;
      9538:data<=-16'd1773;
      9539:data<=-16'd2093;
      9540:data<=-16'd2476;
      9541:data<=-16'd1453;
      9542:data<=-16'd989;
      9543:data<=-16'd922;
      9544:data<=-16'd365;
      9545:data<=-16'd1125;
      9546:data<=-16'd2135;
      9547:data<=-16'd1545;
      9548:data<=-16'd391;
      9549:data<=16'd284;
      9550:data<=16'd464;
      9551:data<=16'd972;
      9552:data<=16'd179;
      9553:data<=-16'd1492;
      9554:data<=16'd2711;
      9555:data<=16'd10275;
      9556:data<=16'd11876;
      9557:data<=16'd10557;
      9558:data<=16'd11473;
      9559:data<=16'd12425;
      9560:data<=16'd12270;
      9561:data<=16'd10484;
      9562:data<=16'd7830;
      9563:data<=16'd7280;
      9564:data<=16'd8624;
      9565:data<=16'd9643;
      9566:data<=16'd9276;
      9567:data<=16'd8580;
      9568:data<=16'd8481;
      9569:data<=16'd7721;
      9570:data<=16'd7507;
      9571:data<=16'd8762;
      9572:data<=16'd8501;
      9573:data<=16'd7107;
      9574:data<=16'd6868;
      9575:data<=16'd7077;
      9576:data<=16'd7068;
      9577:data<=16'd6414;
      9578:data<=16'd5486;
      9579:data<=16'd5145;
      9580:data<=16'd4202;
      9581:data<=16'd3039;
      9582:data<=16'd3509;
      9583:data<=16'd4278;
      9584:data<=16'd3962;
      9585:data<=16'd3771;
      9586:data<=16'd3647;
      9587:data<=16'd2869;
      9588:data<=16'd3272;
      9589:data<=16'd4460;
      9590:data<=16'd3606;
      9591:data<=16'd3033;
      9592:data<=16'd3885;
      9593:data<=16'd2384;
      9594:data<=16'd1198;
      9595:data<=16'd2435;
      9596:data<=-16'd930;
      9597:data<=-16'd7940;
      9598:data<=-16'd9656;
      9599:data<=-16'd7984;
      9600:data<=-16'd8625;
      9601:data<=-16'd9144;
      9602:data<=-16'd7931;
      9603:data<=-16'd7359;
      9604:data<=-16'd7624;
      9605:data<=-16'd7520;
      9606:data<=-16'd6017;
      9607:data<=-16'd4231;
      9608:data<=-16'd4725;
      9609:data<=-16'd5758;
      9610:data<=-16'd5929;
      9611:data<=-16'd6830;
      9612:data<=-16'd6892;
      9613:data<=-16'd6196;
      9614:data<=-16'd6158;
      9615:data<=-16'd5092;
      9616:data<=-16'd5251;
      9617:data<=-16'd6916;
      9618:data<=-16'd5462;
      9619:data<=-16'd3398;
      9620:data<=-16'd3610;
      9621:data<=-16'd3486;
      9622:data<=-16'd2860;
      9623:data<=-16'd2411;
      9624:data<=-16'd2083;
      9625:data<=-16'd1480;
      9626:data<=-16'd405;
      9627:data<=-16'd754;
      9628:data<=-16'd1481;
      9629:data<=-16'd1058;
      9630:data<=-16'd1246;
      9631:data<=-16'd1601;
      9632:data<=-16'd1715;
      9633:data<=-16'd2141;
      9634:data<=-16'd1958;
      9635:data<=-16'd945;
      9636:data<=16'd249;
      9637:data<=-16'd191;
      9638:data<=16'd1172;
      9639:data<=16'd8655;
      9640:data<=16'd13211;
      9641:data<=16'd10815;
      9642:data<=16'd9972;
      9643:data<=16'd10564;
      9644:data<=16'd10463;
      9645:data<=16'd10781;
      9646:data<=16'd9592;
      9647:data<=16'd8692;
      9648:data<=16'd8927;
      9649:data<=16'd9373;
      9650:data<=16'd10615;
      9651:data<=16'd9668;
      9652:data<=16'd7920;
      9653:data<=16'd8214;
      9654:data<=16'd8237;
      9655:data<=16'd8343;
      9656:data<=16'd7902;
      9657:data<=16'd6924;
      9658:data<=16'd6960;
      9659:data<=16'd6184;
      9660:data<=16'd7033;
      9661:data<=16'd8205;
      9662:data<=16'd6734;
      9663:data<=16'd7686;
      9664:data<=16'd7785;
      9665:data<=16'd7000;
      9666:data<=16'd9186;
      9667:data<=16'd6863;
      9668:data<=16'd12768;
      9669:data<=16'd32116;
      9670:data<=16'd30964;
      9671:data<=16'd9759;
      9672:data<=16'd1386;
      9673:data<=16'd3900;
      9674:data<=16'd2525;
      9675:data<=-16'd438;
      9676:data<=16'd920;
      9677:data<=16'd1754;
      9678:data<=16'd129;
      9679:data<=16'd11191;
      9680:data<=16'd29017;
      9681:data<=16'd32608;
      9682:data<=16'd29613;
      9683:data<=16'd23008;
      9684:data<=16'd7714;
      9685:data<=16'd1594;
      9686:data<=16'd7702;
      9687:data<=16'd9820;
      9688:data<=16'd5112;
      9689:data<=-16'd3604;
      9690:data<=-16'd9235;
      9691:data<=-16'd4816;
      9692:data<=16'd2228;
      9693:data<=16'd3389;
      9694:data<=-16'd852;
      9695:data<=-16'd4880;
      9696:data<=-16'd3301;
      9697:data<=-16'd1343;
      9698:data<=-16'd4998;
      9699:data<=-16'd5742;
      9700:data<=-16'd1436;
      9701:data<=-16'd785;
      9702:data<=16'd2126;
      9703:data<=16'd4692;
      9704:data<=-16'd7514;
      9705:data<=-16'd14562;
      9706:data<=-16'd3576;
      9707:data<=-16'd1303;
      9708:data<=-16'd9310;
      9709:data<=-16'd10111;
      9710:data<=-16'd7118;
      9711:data<=-16'd4937;
      9712:data<=-16'd3366;
      9713:data<=-16'd17;
      9714:data<=16'd658;
      9715:data<=-16'd6266;
      9716:data<=-16'd6164;
      9717:data<=-16'd2228;
      9718:data<=-16'd3099;
      9719:data<=16'd4364;
      9720:data<=16'd3287;
      9721:data<=-16'd8238;
      9722:data<=16'd804;
      9723:data<=16'd4449;
      9724:data<=-16'd11814;
      9725:data<=-16'd10172;
      9726:data<=16'd2817;
      9727:data<=16'd7412;
      9728:data<=16'd7144;
      9729:data<=16'd2722;
      9730:data<=16'd7417;
      9731:data<=16'd16029;
      9732:data<=16'd11623;
      9733:data<=16'd8710;
      9734:data<=16'd10793;
      9735:data<=16'd11074;
      9736:data<=16'd13893;
      9737:data<=16'd10022;
      9738:data<=16'd2349;
      9739:data<=16'd3542;
      9740:data<=16'd4141;
      9741:data<=16'd5582;
      9742:data<=16'd16120;
      9743:data<=16'd19685;
      9744:data<=16'd12609;
      9745:data<=16'd13723;
      9746:data<=16'd18803;
      9747:data<=16'd11923;
      9748:data<=16'd3789;
      9749:data<=16'd6470;
      9750:data<=16'd11891;
      9751:data<=16'd13405;
      9752:data<=16'd11731;
      9753:data<=16'd9784;
      9754:data<=16'd7319;
      9755:data<=16'd4886;
      9756:data<=16'd8586;
      9757:data<=16'd7717;
      9758:data<=-16'd2764;
      9759:data<=-16'd1149;
      9760:data<=16'd5215;
      9761:data<=-16'd212;
      9762:data<=16'd1485;
      9763:data<=16'd6775;
      9764:data<=-16'd2258;
      9765:data<=-16'd8410;
      9766:data<=-16'd4073;
      9767:data<=-16'd3888;
      9768:data<=-16'd4091;
      9769:data<=16'd696;
      9770:data<=-16'd6693;
      9771:data<=-16'd25243;
      9772:data<=-16'd27219;
      9773:data<=-16'd18927;
      9774:data<=-16'd21155;
      9775:data<=-16'd24127;
      9776:data<=-16'd25972;
      9777:data<=-16'd24694;
      9778:data<=-16'd12740;
      9779:data<=-16'd11697;
      9780:data<=-16'd20104;
      9781:data<=-16'd16313;
      9782:data<=-16'd14028;
      9783:data<=-16'd16233;
      9784:data<=-16'd12703;
      9785:data<=-16'd11709;
      9786:data<=-16'd14431;
      9787:data<=-16'd16412;
      9788:data<=-16'd12019;
      9789:data<=-16'd8329;
      9790:data<=-16'd20501;
      9791:data<=-16'd24777;
      9792:data<=-16'd12094;
      9793:data<=-16'd11476;
      9794:data<=-16'd15907;
      9795:data<=-16'd16516;
      9796:data<=-16'd22136;
      9797:data<=-16'd21623;
      9798:data<=-16'd18240;
      9799:data<=-16'd18494;
      9800:data<=-16'd17509;
      9801:data<=-16'd19722;
      9802:data<=-16'd15095;
      9803:data<=-16'd9417;
      9804:data<=-16'd18759;
      9805:data<=-16'd17799;
      9806:data<=-16'd8901;
      9807:data<=-16'd15741;
      9808:data<=-16'd15822;
      9809:data<=-16'd9098;
      9810:data<=-16'd13916;
      9811:data<=-16'd12569;
      9812:data<=-16'd6206;
      9813:data<=-16'd9568;
      9814:data<=-16'd10257;
      9815:data<=-16'd1996;
      9816:data<=16'd6294;
      9817:data<=16'd11051;
      9818:data<=16'd14231;
      9819:data<=16'd12927;
      9820:data<=16'd6516;
      9821:data<=16'd9242;
      9822:data<=16'd18656;
      9823:data<=16'd15896;
      9824:data<=16'd12157;
      9825:data<=16'd18066;
      9826:data<=16'd16624;
      9827:data<=16'd10687;
      9828:data<=16'd13690;
      9829:data<=16'd14650;
      9830:data<=16'd9996;
      9831:data<=16'd10712;
      9832:data<=16'd11301;
      9833:data<=16'd7260;
      9834:data<=16'd8345;
      9835:data<=16'd12330;
      9836:data<=16'd12942;
      9837:data<=16'd13191;
      9838:data<=16'd13605;
      9839:data<=16'd15292;
      9840:data<=16'd13517;
      9841:data<=16'd7180;
      9842:data<=16'd11007;
      9843:data<=16'd13679;
      9844:data<=16'd3089;
      9845:data<=16'd3660;
      9846:data<=16'd9044;
      9847:data<=16'd4258;
      9848:data<=16'd10862;
      9849:data<=16'd19893;
      9850:data<=16'd17573;
      9851:data<=16'd18923;
      9852:data<=16'd17754;
      9853:data<=16'd16052;
      9854:data<=16'd20510;
      9855:data<=16'd14909;
      9856:data<=16'd8319;
      9857:data<=16'd9633;
      9858:data<=16'd11793;
      9859:data<=16'd19011;
      9860:data<=16'd12634;
      9861:data<=-16'd7022;
      9862:data<=-16'd7257;
      9863:data<=-16'd2937;
      9864:data<=-16'd7118;
      9865:data<=-16'd2564;
      9866:data<=-16'd1084;
      9867:data<=-16'd5476;
      9868:data<=-16'd1061;
      9869:data<=16'd3253;
      9870:data<=-16'd174;
      9871:data<=-16'd4531;
      9872:data<=-16'd1219;
      9873:data<=16'd4827;
      9874:data<=16'd1615;
      9875:data<=-16'd2366;
      9876:data<=-16'd3327;
      9877:data<=-16'd6169;
      9878:data<=-16'd1359;
      9879:data<=16'd4868;
      9880:data<=16'd2171;
      9881:data<=16'd640;
      9882:data<=16'd2290;
      9883:data<=16'd2852;
      9884:data<=16'd766;
      9885:data<=-16'd667;
      9886:data<=16'd5080;
      9887:data<=16'd4687;
      9888:data<=-16'd4379;
      9889:data<=-16'd1897;
      9890:data<=16'd4619;
      9891:data<=16'd1750;
      9892:data<=-16'd611;
      9893:data<=16'd1665;
      9894:data<=16'd4334;
      9895:data<=16'd3391;
      9896:data<=16'd14;
      9897:data<=-16'd983;
      9898:data<=-16'd2243;
      9899:data<=-16'd432;
      9900:data<=16'd5617;
      9901:data<=16'd2561;
      9902:data<=-16'd6299;
      9903:data<=-16'd7667;
      9904:data<=-16'd4278;
      9905:data<=16'd2455;
      9906:data<=16'd12778;
      9907:data<=16'd15928;
      9908:data<=16'd10730;
      9909:data<=16'd10305;
      9910:data<=16'd13844;
      9911:data<=16'd12548;
      9912:data<=16'd11201;
      9913:data<=16'd11397;
      9914:data<=16'd11832;
      9915:data<=16'd16089;
      9916:data<=16'd14251;
      9917:data<=16'd5671;
      9918:data<=16'd6968;
      9919:data<=16'd12160;
      9920:data<=16'd10367;
      9921:data<=16'd9185;
      9922:data<=16'd10422;
      9923:data<=16'd9661;
      9924:data<=16'd9191;
      9925:data<=16'd12393;
      9926:data<=16'd14266;
      9927:data<=16'd11492;
      9928:data<=16'd10796;
      9929:data<=16'd9527;
      9930:data<=16'd5548;
      9931:data<=16'd5614;
      9932:data<=16'd4748;
      9933:data<=16'd5953;
      9934:data<=16'd12152;
      9935:data<=16'd8111;
      9936:data<=16'd719;
      9937:data<=16'd917;
      9938:data<=16'd1513;
      9939:data<=16'd4223;
      9940:data<=16'd5010;
      9941:data<=16'd3621;
      9942:data<=16'd4939;
      9943:data<=-16'd1092;
      9944:data<=-16'd2575;
      9945:data<=16'd4827;
      9946:data<=16'd1245;
      9947:data<=16'd787;
      9948:data<=16'd3560;
      9949:data<=-16'd9614;
      9950:data<=-16'd18907;
      9951:data<=-16'd18419;
      9952:data<=-16'd18410;
      9953:data<=-16'd14307;
      9954:data<=-16'd11238;
      9955:data<=-16'd7489;
      9956:data<=-16'd4214;
      9957:data<=-16'd7156;
      9958:data<=-16'd5852;
      9959:data<=-16'd6931;
      9960:data<=-16'd10090;
      9961:data<=-16'd5416;
      9962:data<=-16'd8263;
      9963:data<=-16'd8616;
      9964:data<=-16'd974;
      9965:data<=-16'd8150;
      9966:data<=-16'd12305;
      9967:data<=-16'd7468;
      9968:data<=-16'd11412;
      9969:data<=-16'd10141;
      9970:data<=-16'd7815;
      9971:data<=-16'd10871;
      9972:data<=-16'd8792;
      9973:data<=-16'd11374;
      9974:data<=-16'd10537;
      9975:data<=-16'd4755;
      9976:data<=-16'd12480;
      9977:data<=-16'd14066;
      9978:data<=-16'd6193;
      9979:data<=-16'd8608;
      9980:data<=-16'd11077;
      9981:data<=-16'd12117;
      9982:data<=-16'd11324;
      9983:data<=-16'd4272;
      9984:data<=-16'd6860;
      9985:data<=-16'd12806;
      9986:data<=-16'd9665;
      9987:data<=-16'd5245;
      9988:data<=-16'd1293;
      9989:data<=-16'd5635;
      9990:data<=-16'd13138;
      9991:data<=-16'd7429;
      9992:data<=-16'd5313;
      9993:data<=-16'd8443;
      9994:data<=16'd3950;
      9995:data<=16'd14408;
      9996:data<=16'd8909;
      9997:data<=16'd8150;
      9998:data<=16'd12313;
      9999:data<=16'd4757;
      10000:data<=-16'd200;
      10001:data<=16'd9574;
      10002:data<=16'd10731;
      10003:data<=16'd1359;
      10004:data<=16'd1679;
      10005:data<=16'd3574;
      10006:data<=-16'd428;
      10007:data<=-16'd7454;
      10008:data<=-16'd16073;
      10009:data<=-16'd12963;
      10010:data<=-16'd5372;
      10011:data<=-16'd7705;
      10012:data<=-16'd9054;
      10013:data<=-16'd10107;
      10014:data<=-16'd9653;
      10015:data<=-16'd2143;
      10016:data<=-16'd4372;
      10017:data<=-16'd10894;
      10018:data<=-16'd8210;
      10019:data<=-16'd5077;
      10020:data<=-16'd1871;
      10021:data<=-16'd4551;
      10022:data<=-16'd10561;
      10023:data<=-16'd6152;
      10024:data<=-16'd5821;
      10025:data<=-16'd7301;
      10026:data<=-16'd4190;
      10027:data<=-16'd14070;
      10028:data<=-16'd15985;
      10029:data<=-16'd3997;
      10030:data<=-16'd6648;
      10031:data<=-16'd7912;
      10032:data<=-16'd4255;
      10033:data<=-16'd9342;
      10034:data<=-16'd6652;
      10035:data<=-16'd4719;
      10036:data<=-16'd7333;
      10037:data<=-16'd2637;
      10038:data<=-16'd11932;
      10039:data<=-16'd27457;
      10040:data<=-16'd26250;
      10041:data<=-16'd23673;
      10042:data<=-16'd22193;
      10043:data<=-16'd19237;
      10044:data<=-16'd19371;
      10045:data<=-16'd15976;
      10046:data<=-16'd18269;
      10047:data<=-16'd25877;
      10048:data<=-16'd22845;
      10049:data<=-16'd18912;
      10050:data<=-16'd19745;
      10051:data<=-16'd16181;
      10052:data<=-16'd11283;
      10053:data<=-16'd11483;
      10054:data<=-16'd15623;
      10055:data<=-16'd14959;
      10056:data<=-16'd10196;
      10057:data<=-16'd11227;
      10058:data<=-16'd13459;
      10059:data<=-16'd11916;
      10060:data<=-16'd9379;
      10061:data<=-16'd6032;
      10062:data<=-16'd2987;
      10063:data<=-16'd108;
      10064:data<=-16'd992;
      10065:data<=-16'd3927;
      10066:data<=-16'd1216;
      10067:data<=-16'd1800;
      10068:data<=-16'd4558;
      10069:data<=-16'd1312;
      10070:data<=-16'd3024;
      10071:data<=-16'd2617;
      10072:data<=16'd4037;
      10073:data<=16'd1760;
      10074:data<=16'd1894;
      10075:data<=16'd5059;
      10076:data<=-16'd717;
      10077:data<=-16'd939;
      10078:data<=16'd549;
      10079:data<=-16'd1871;
      10080:data<=16'd3536;
      10081:data<=16'd3639;
      10082:data<=-16'd132;
      10083:data<=16'd9072;
      10084:data<=16'd17165;
      10085:data<=16'd17820;
      10086:data<=16'd18201;
      10087:data<=16'd16172;
      10088:data<=16'd15852;
      10089:data<=16'd18428;
      10090:data<=16'd20154;
      10091:data<=16'd21581;
      10092:data<=16'd20192;
      10093:data<=16'd16043;
      10094:data<=16'd14361;
      10095:data<=16'd17185;
      10096:data<=16'd17540;
      10097:data<=16'd13218;
      10098:data<=16'd16657;
      10099:data<=16'd22979;
      10100:data<=16'd18025;
      10101:data<=16'd12692;
      10102:data<=16'd14236;
      10103:data<=16'd16745;
      10104:data<=16'd18225;
      10105:data<=16'd15819;
      10106:data<=16'd15693;
      10107:data<=16'd20058;
      10108:data<=16'd18026;
      10109:data<=16'd11903;
      10110:data<=16'd7065;
      10111:data<=16'd7106;
      10112:data<=16'd14569;
      10113:data<=16'd12524;
      10114:data<=16'd1525;
      10115:data<=16'd2044;
      10116:data<=16'd5897;
      10117:data<=16'd7119;
      10118:data<=16'd11247;
      10119:data<=16'd6017;
      10120:data<=-16'd393;
      10121:data<=16'd7853;
      10122:data<=16'd10191;
      10123:data<=16'd479;
      10124:data<=-16'd1251;
      10125:data<=16'd2664;
      10126:data<=16'd4472;
      10127:data<=16'd3451;
      10128:data<=-16'd7215;
      10129:data<=-16'd17561;
      10130:data<=-16'd14892;
      10131:data<=-16'd11371;
      10132:data<=-16'd12126;
      10133:data<=-16'd11492;
      10134:data<=-16'd11655;
      10135:data<=-16'd7827;
      10136:data<=-16'd2012;
      10137:data<=-16'd6357;
      10138:data<=-16'd11825;
      10139:data<=-16'd8238;
      10140:data<=-16'd2123;
      10141:data<=16'd2358;
      10142:data<=16'd214;
      10143:data<=-16'd4473;
      10144:data<=-16'd919;
      10145:data<=-16'd1575;
      10146:data<=-16'd7451;
      10147:data<=-16'd73;
      10148:data<=16'd3955;
      10149:data<=-16'd5046;
      10150:data<=-16'd3475;
      10151:data<=-16'd35;
      10152:data<=-16'd2487;
      10153:data<=16'd5768;
      10154:data<=16'd6082;
      10155:data<=-16'd4212;
      10156:data<=16'd1759;
      10157:data<=16'd5145;
      10158:data<=-16'd2934;
      10159:data<=-16'd1309;
      10160:data<=16'd1507;
      10161:data<=16'd5297;
      10162:data<=16'd10875;
      10163:data<=16'd2619;
      10164:data<=-16'd558;
      10165:data<=16'd7312;
      10166:data<=16'd6652;
      10167:data<=16'd8813;
      10168:data<=16'd13561;
      10169:data<=16'd11271;
      10170:data<=16'd12419;
      10171:data<=16'd11765;
      10172:data<=16'd13282;
      10173:data<=16'd26874;
      10174:data<=16'd32767;
      10175:data<=16'd28911;
      10176:data<=16'd28013;
      10177:data<=16'd26224;
      10178:data<=16'd26119;
      10179:data<=16'd27008;
      10180:data<=16'd23388;
      10181:data<=16'd21182;
      10182:data<=16'd21520;
      10183:data<=16'd21426;
      10184:data<=16'd21290;
      10185:data<=16'd21464;
      10186:data<=16'd21690;
      10187:data<=16'd20163;
      10188:data<=16'd19136;
      10189:data<=16'd17814;
      10190:data<=16'd14234;
      10191:data<=16'd15227;
      10192:data<=16'd17629;
      10193:data<=16'd16594;
      10194:data<=16'd16310;
      10195:data<=16'd11183;
      10196:data<=16'd5081;
      10197:data<=16'd9679;
      10198:data<=16'd15606;
      10199:data<=16'd14998;
      10200:data<=16'd12090;
      10201:data<=16'd10037;
      10202:data<=16'd10067;
      10203:data<=16'd8698;
      10204:data<=16'd6084;
      10205:data<=16'd4516;
      10206:data<=16'd4770;
      10207:data<=16'd8064;
      10208:data<=16'd5661;
      10209:data<=16'd1231;
      10210:data<=16'd6384;
      10211:data<=16'd7395;
      10212:data<=16'd3664;
      10213:data<=16'd4775;
      10214:data<=16'd787;
      10215:data<=16'd741;
      10216:data<=16'd3338;
      10217:data<=-16'd11920;
      10218:data<=-16'd22157;
      10219:data<=-16'd16730;
      10220:data<=-16'd20430;
      10221:data<=-16'd25566;
      10222:data<=-16'd24439;
      10223:data<=-16'd26233;
      10224:data<=-16'd25012;
      10225:data<=-16'd24427;
      10226:data<=-16'd28154;
      10227:data<=-16'd24691;
      10228:data<=-16'd19628;
      10229:data<=-16'd23514;
      10230:data<=-16'd26435;
      10231:data<=-16'd21957;
      10232:data<=-16'd21739;
      10233:data<=-16'd25669;
      10234:data<=-16'd22234;
      10235:data<=-16'd20101;
      10236:data<=-16'd20926;
      10237:data<=-16'd15312;
      10238:data<=-16'd16803;
      10239:data<=-16'd21605;
      10240:data<=-16'd16895;
      10241:data<=-16'd19828;
      10242:data<=-16'd22116;
      10243:data<=-16'd11888;
      10244:data<=-16'd10786;
      10245:data<=-16'd12195;
      10246:data<=-16'd10696;
      10247:data<=-16'd19842;
      10248:data<=-16'd20213;
      10249:data<=-16'd12158;
      10250:data<=-16'd16315;
      10251:data<=-16'd18195;
      10252:data<=-16'd14577;
      10253:data<=-16'd15335;
      10254:data<=-16'd16495;
      10255:data<=-16'd18691;
      10256:data<=-16'd15831;
      10257:data<=-16'd9994;
      10258:data<=-16'd12725;
      10259:data<=-16'd13486;
      10260:data<=-16'd9417;
      10261:data<=-16'd4602;
      10262:data<=16'd4910;
      10263:data<=16'd7403;
      10264:data<=16'd4510;
      10265:data<=16'd7219;
      10266:data<=16'd5750;
      10267:data<=16'd3623;
      10268:data<=16'd5145;
      10269:data<=16'd1798;
      10270:data<=16'd984;
      10271:data<=16'd3266;
      10272:data<=16'd4322;
      10273:data<=16'd9081;
      10274:data<=16'd9380;
      10275:data<=16'd5771;
      10276:data<=16'd6681;
      10277:data<=16'd4752;
      10278:data<=16'd3797;
      10279:data<=16'd8398;
      10280:data<=16'd7036;
      10281:data<=16'd2573;
      10282:data<=16'd4323;
      10283:data<=16'd7758;
      10284:data<=16'd9021;
      10285:data<=16'd9949;
      10286:data<=16'd8437;
      10287:data<=16'd3838;
      10288:data<=16'd4637;
      10289:data<=16'd8822;
      10290:data<=16'd4734;
      10291:data<=-16'd1092;
      10292:data<=-16'd453;
      10293:data<=16'd306;
      10294:data<=-16'd1503;
      10295:data<=-16'd1729;
      10296:data<=16'd2860;
      10297:data<=16'd4614;
      10298:data<=-16'd1462;
      10299:data<=-16'd3576;
      10300:data<=-16'd3268;
      10301:data<=-16'd6009;
      10302:data<=-16'd4067;
      10303:data<=-16'd3107;
      10304:data<=-16'd2194;
      10305:data<=16'd1037;
      10306:data<=-16'd9920;
      10307:data<=-16'd22019;
      10308:data<=-16'd22112;
      10309:data<=-16'd27338;
      10310:data<=-16'd27693;
      10311:data<=-16'd18158;
      10312:data<=-16'd16976;
      10313:data<=-16'd16603;
      10314:data<=-16'd14859;
      10315:data<=-16'd17526;
      10316:data<=-16'd15778;
      10317:data<=-16'd14439;
      10318:data<=-16'd14886;
      10319:data<=-16'd11082;
      10320:data<=-16'd9690;
      10321:data<=-16'd10246;
      10322:data<=-16'd11550;
      10323:data<=-16'd12236;
      10324:data<=-16'd7031;
      10325:data<=-16'd8120;
      10326:data<=-16'd15872;
      10327:data<=-16'd15935;
      10328:data<=-16'd17691;
      10329:data<=-16'd24459;
      10330:data<=-16'd22656;
      10331:data<=-16'd17723;
      10332:data<=-16'd19751;
      10333:data<=-16'd20688;
      10334:data<=-16'd15402;
      10335:data<=-16'd13133;
      10336:data<=-16'd13402;
      10337:data<=-16'd12182;
      10338:data<=-16'd17644;
      10339:data<=-16'd20621;
      10340:data<=-16'd13461;
      10341:data<=-16'd12715;
      10342:data<=-16'd12971;
      10343:data<=-16'd7990;
      10344:data<=-16'd11398;
      10345:data<=-16'd12026;
      10346:data<=-16'd3885;
      10347:data<=-16'd1445;
      10348:data<=-16'd3683;
      10349:data<=-16'd6209;
      10350:data<=-16'd570;
      10351:data<=16'd12960;
      10352:data<=16'd16343;
      10353:data<=16'd15315;
      10354:data<=16'd15476;
      10355:data<=16'd12516;
      10356:data<=16'd17203;
      10357:data<=16'd16113;
      10358:data<=16'd5899;
      10359:data<=16'd12313;
      10360:data<=16'd17790;
      10361:data<=16'd11850;
      10362:data<=16'd15931;
      10363:data<=16'd16900;
      10364:data<=16'd12481;
      10365:data<=16'd17423;
      10366:data<=16'd17888;
      10367:data<=16'd14273;
      10368:data<=16'd15769;
      10369:data<=16'd15782;
      10370:data<=16'd15192;
      10371:data<=16'd12452;
      10372:data<=16'd8000;
      10373:data<=16'd8113;
      10374:data<=16'd7304;
      10375:data<=16'd8055;
      10376:data<=16'd14807;
      10377:data<=16'd14639;
      10378:data<=16'd7050;
      10379:data<=16'd9564;
      10380:data<=16'd21071;
      10381:data<=16'd20600;
      10382:data<=16'd12590;
      10383:data<=16'd18230;
      10384:data<=16'd24577;
      10385:data<=16'd19221;
      10386:data<=16'd17464;
      10387:data<=16'd18231;
      10388:data<=16'd15737;
      10389:data<=16'd16237;
      10390:data<=16'd17247;
      10391:data<=16'd17220;
      10392:data<=16'd16618;
      10393:data<=16'd15430;
      10394:data<=16'd14164;
      10395:data<=16'd5515;
      10396:data<=-16'd3800;
      10397:data<=-16'd3650;
      10398:data<=-16'd3985;
      10399:data<=-16'd4440;
      10400:data<=-16'd1136;
      10401:data<=-16'd314;
      10402:data<=-16'd86;
      10403:data<=-16'd2118;
      10404:data<=-16'd2406;
      10405:data<=16'd5269;
      10406:data<=16'd5174;
      10407:data<=-16'd30;
      10408:data<=16'd3563;
      10409:data<=16'd2124;
      10410:data<=-16'd3054;
      10411:data<=16'd1554;
      10412:data<=16'd4716;
      10413:data<=16'd926;
      10414:data<=-16'd299;
      10415:data<=16'd2584;
      10416:data<=16'd3526;
      10417:data<=16'd1495;
      10418:data<=16'd3469;
      10419:data<=16'd7356;
      10420:data<=16'd4545;
      10421:data<=-16'd399;
      10422:data<=16'd1111;
      10423:data<=16'd4978;
      10424:data<=16'd805;
      10425:data<=-16'd4355;
      10426:data<=16'd2215;
      10427:data<=16'd7459;
      10428:data<=16'd3798;
      10429:data<=16'd3644;
      10430:data<=16'd5673;
      10431:data<=16'd6413;
      10432:data<=16'd6457;
      10433:data<=16'd3712;
      10434:data<=16'd3206;
      10435:data<=16'd106;
      10436:data<=-16'd4925;
      10437:data<=16'd238;
      10438:data<=16'd334;
      10439:data<=-16'd4613;
      10440:data<=16'd10111;
      10441:data<=16'd25061;
      10442:data<=16'd20221;
      10443:data<=16'd14800;
      10444:data<=16'd12906;
      10445:data<=16'd9867;
      10446:data<=16'd12295;
      10447:data<=16'd14220;
      10448:data<=16'd10710;
      10449:data<=16'd12328;
      10450:data<=16'd15720;
      10451:data<=16'd8627;
      10452:data<=16'd4687;
      10453:data<=16'd11110;
      10454:data<=16'd10084;
      10455:data<=16'd7336;
      10456:data<=16'd9815;
      10457:data<=16'd6416;
      10458:data<=16'd9903;
      10459:data<=16'd18271;
      10460:data<=16'd12313;
      10461:data<=16'd9843;
      10462:data<=16'd14428;
      10463:data<=16'd9797;
      10464:data<=16'd7612;
      10465:data<=16'd10132;
      10466:data<=16'd10116;
      10467:data<=16'd11514;
      10468:data<=16'd11521;
      10469:data<=16'd11377;
      10470:data<=16'd9529;
      10471:data<=16'd2937;
      10472:data<=16'd2221;
      10473:data<=16'd3460;
      10474:data<=16'd1902;
      10475:data<=16'd5022;
      10476:data<=16'd5685;
      10477:data<=16'd3941;
      10478:data<=16'd4538;
      10479:data<=16'd1623;
      10480:data<=16'd2560;
      10481:data<=16'd6411;
      10482:data<=16'd4425;
      10483:data<=16'd1968;
      10484:data<=-16'd7501;
      10485:data<=-16'd18982;
      10486:data<=-16'd14333;
      10487:data<=-16'd10857;
      10488:data<=-16'd15891;
      10489:data<=-16'd10742;
      10490:data<=-16'd5071;
      10491:data<=-16'd8611;
      10492:data<=-16'd10530;
      10493:data<=-16'd10517;
      10494:data<=-16'd9203;
      10495:data<=-16'd5556;
      10496:data<=-16'd5844;
      10497:data<=-16'd8113;
      10498:data<=-16'd7511;
      10499:data<=-16'd6813;
      10500:data<=-16'd7755;
      10501:data<=-16'd10364;
      10502:data<=-16'd12508;
      10503:data<=-16'd11593;
      10504:data<=-16'd10948;
      10505:data<=-16'd9979;
      10506:data<=-16'd8241;
      10507:data<=-16'd13696;
      10508:data<=-16'd18055;
      10509:data<=-16'd10587;
      10510:data<=-16'd7984;
      10511:data<=-16'd13432;
      10512:data<=-16'd10405;
      10513:data<=-16'd4726;
      10514:data<=-16'd4757;
      10515:data<=-16'd8590;
      10516:data<=-16'd14871;
      10517:data<=-16'd13318;
      10518:data<=-16'd8047;
      10519:data<=-16'd12298;
      10520:data<=-16'd13881;
      10521:data<=-16'd8017;
      10522:data<=-16'd6636;
      10523:data<=-16'd8443;
      10524:data<=-16'd9680;
      10525:data<=-16'd7664;
      10526:data<=-16'd5882;
      10527:data<=-16'd13204;
      10528:data<=-16'd14069;
      10529:data<=16'd879;
      10530:data<=16'd10933;
      10531:data<=16'd12261;
      10532:data<=16'd12408;
      10533:data<=16'd7406;
      10534:data<=16'd2493;
      10535:data<=16'd3292;
      10536:data<=16'd4020;
      10537:data<=16'd1325;
      10538:data<=-16'd625;
      10539:data<=16'd2695;
      10540:data<=16'd1679;
      10541:data<=-16'd9039;
      10542:data<=-16'd11373;
      10543:data<=-16'd4038;
      10544:data<=-16'd5142;
      10545:data<=-16'd9435;
      10546:data<=-16'd6946;
      10547:data<=-16'd4278;
      10548:data<=-16'd3566;
      10549:data<=-16'd3157;
      10550:data<=-16'd6428;
      10551:data<=-16'd11568;
      10552:data<=-16'd10111;
      10553:data<=-16'd2275;
      10554:data<=16'd1997;
      10555:data<=16'd2362;
      10556:data<=16'd3789;
      10557:data<=16'd3413;
      10558:data<=16'd1894;
      10559:data<=16'd837;
      10560:data<=-16'd1829;
      10561:data<=-16'd1624;
      10562:data<=16'd1155;
      10563:data<=16'd1016;
      10564:data<=16'd699;
      10565:data<=16'd50;
      10566:data<=-16'd2447;
      10567:data<=-16'd3086;
      10568:data<=-16'd2613;
      10569:data<=-16'd1947;
      10570:data<=-16'd1682;
      10571:data<=-16'd1739;
      10572:data<=16'd1027;
      10573:data<=-16'd3295;
      10574:data<=-16'd17914;
      10575:data<=-16'd22239;
      10576:data<=-16'd16055;
      10577:data<=-16'd16509;
      10578:data<=-16'd19537;
      10579:data<=-16'd19247;
      10580:data<=-16'd18914;
      10581:data<=-16'd17752;
      10582:data<=-16'd15945;
      10583:data<=-16'd14305;
      10584:data<=-16'd13538;
      10585:data<=-16'd15033;
      10586:data<=-16'd16437;
      10587:data<=-16'd16349;
      10588:data<=-16'd14882;
      10589:data<=-16'd12687;
      10590:data<=-16'd12261;
      10591:data<=-16'd12433;
      10592:data<=-16'd11044;
      10593:data<=-16'd7600;
      10594:data<=-16'd3324;
      10595:data<=-16'd3410;
      10596:data<=-16'd6382;
      10597:data<=-16'd5903;
      10598:data<=-16'd3183;
      10599:data<=-16'd1942;
      10600:data<=-16'd5001;
      10601:data<=-16'd8443;
      10602:data<=-16'd5204;
      10603:data<=-16'd2504;
      10604:data<=-16'd4282;
      10605:data<=-16'd2743;
      10606:data<=-16'd1051;
      10607:data<=-16'd2861;
      10608:data<=-16'd4040;
      10609:data<=-16'd4281;
      10610:data<=-16'd3089;
      10611:data<=-16'd1950;
      10612:data<=-16'd2290;
      10613:data<=-16'd1616;
      10614:data<=-16'd1821;
      10615:data<=-16'd1727;
      10616:data<=-16'd161;
      10617:data<=-16'd45;
      10618:data<=16'd6299;
      10619:data<=16'd18055;
      10620:data<=16'd20721;
      10621:data<=16'd17062;
      10622:data<=16'd15732;
      10623:data<=16'd15952;
      10624:data<=16'd17459;
      10625:data<=16'd17926;
      10626:data<=16'd16540;
      10627:data<=16'd15338;
      10628:data<=16'd13700;
      10629:data<=16'd13383;
      10630:data<=16'd14225;
      10631:data<=16'd13678;
      10632:data<=16'd13565;
      10633:data<=16'd14308;
      10634:data<=16'd14502;
      10635:data<=16'd14161;
      10636:data<=16'd13955;
      10637:data<=16'd14316;
      10638:data<=16'd13499;
      10639:data<=16'd12223;
      10640:data<=16'd11906;
      10641:data<=16'd11590;
      10642:data<=16'd12574;
      10643:data<=16'd12696;
      10644:data<=16'd10520;
      10645:data<=16'd9012;
      10646:data<=16'd4376;
      10647:data<=-16'd1340;
      10648:data<=-16'd462;
      10649:data<=16'd1917;
      10650:data<=16'd2074;
      10651:data<=16'd2411;
      10652:data<=16'd3339;
      10653:data<=16'd4746;
      10654:data<=16'd2848;
      10655:data<=16'd1465;
      10656:data<=16'd4347;
      10657:data<=16'd3058;
      10658:data<=16'd1844;
      10659:data<=16'd3727;
      10660:data<=16'd1124;
      10661:data<=16'd2009;
      10662:data<=16'd1662;
      10663:data<=-16'd10355;
      10664:data<=-16'd15396;
      10665:data<=-16'd11482;
      10666:data<=-16'd12402;
      10667:data<=-16'd11764;
      10668:data<=-16'd10060;
      10669:data<=-16'd10525;
      10670:data<=-16'd8223;
      10671:data<=-16'd7139;
      10672:data<=-16'd7417;
      10673:data<=-16'd7092;
      10674:data<=-16'd7667;
      10675:data<=-16'd5489;
      10676:data<=-16'd3685;
      10677:data<=-16'd4073;
      10678:data<=-16'd2557;
      10679:data<=-16'd3388;
      10680:data<=-16'd4899;
      10681:data<=-16'd3698;
      10682:data<=-16'd5227;
      10683:data<=-16'd5474;
      10684:data<=-16'd1641;
      10685:data<=-16'd613;
      10686:data<=-16'd1340;
      10687:data<=-16'd1331;
      10688:data<=-16'd2159;
      10689:data<=-16'd2581;
      10690:data<=-16'd2275;
      10691:data<=-16'd1395;
      10692:data<=16'd622;
      10693:data<=16'd1468;
      10694:data<=16'd121;
      10695:data<=16'd250;
      10696:data<=16'd1378;
      10697:data<=-16'd347;
      10698:data<=16'd773;
      10699:data<=16'd6598;
      10700:data<=16'd8734;
      10701:data<=16'd10792;
      10702:data<=16'd13711;
      10703:data<=16'd9438;
      10704:data<=16'd7473;
      10705:data<=16'd9530;
      10706:data<=16'd5510;
      10707:data<=16'd9100;
      10708:data<=16'd22620;
      10709:data<=16'd26785;
      10710:data<=16'd25642;
      10711:data<=16'd25846;
      10712:data<=16'd21607;
      10713:data<=16'd18942;
      10714:data<=16'd20447;
      10715:data<=16'd20275;
      10716:data<=16'd19714;
      10717:data<=16'd18907;
      10718:data<=16'd16775;
      10719:data<=16'd15705;
      10720:data<=16'd15866;
      10721:data<=16'd16571;
      10722:data<=16'd16868;
      10723:data<=16'd15499;
      10724:data<=16'd13368;
      10725:data<=16'd12534;
      10726:data<=16'd13582;
      10727:data<=16'd13160;
      10728:data<=16'd11069;
      10729:data<=16'd11940;
      10730:data<=16'd12716;
      10731:data<=16'd9641;
      10732:data<=16'd7633;
      10733:data<=16'd8564;
      10734:data<=16'd10002;
      10735:data<=16'd9982;
      10736:data<=16'd8135;
      10737:data<=16'd8452;
      10738:data<=16'd9967;
      10739:data<=16'd8047;
      10740:data<=16'd5817;
      10741:data<=16'd5395;
      10742:data<=16'd5494;
      10743:data<=16'd6393;
      10744:data<=16'd5463;
      10745:data<=16'd3353;
      10746:data<=16'd3744;
      10747:data<=16'd4026;
      10748:data<=16'd2737;
      10749:data<=16'd3002;
      10750:data<=16'd3824;
      10751:data<=-16'd1842;
      10752:data<=-16'd16075;
      10753:data<=-16'd27261;
      10754:data<=-16'd27875;
      10755:data<=-16'd25680;
      10756:data<=-16'd25153;
      10757:data<=-16'd23681;
      10758:data<=-16'd22021;
      10759:data<=-16'd22889;
      10760:data<=-16'd24968;
      10761:data<=-16'd23309;
      10762:data<=-16'd20407;
      10763:data<=-16'd21619;
      10764:data<=-16'd22242;
      10765:data<=-16'd20383;
      10766:data<=-16'd19241;
      10767:data<=-16'd17787;
      10768:data<=-16'd17890;
      10769:data<=-16'd19177;
      10770:data<=-16'd17843;
      10771:data<=-16'd16539;
      10772:data<=-16'd16175;
      10773:data<=-16'd15415;
      10774:data<=-16'd15161;
      10775:data<=-16'd15176;
      10776:data<=-16'd16258;
      10777:data<=-16'd16004;
      10778:data<=-16'd13593;
      10779:data<=-16'd14085;
      10780:data<=-16'd14703;
      10781:data<=-16'd13376;
      10782:data<=-16'd13728;
      10783:data<=-16'd13050;
      10784:data<=-16'd12073;
      10785:data<=-16'd13194;
      10786:data<=-16'd13397;
      10787:data<=-16'd12915;
      10788:data<=-16'd11367;
      10789:data<=-16'd10085;
      10790:data<=-16'd10971;
      10791:data<=-16'd10204;
      10792:data<=-16'd10577;
      10793:data<=-16'd13059;
      10794:data<=-16'd13964;
      10795:data<=-16'd15393;
      10796:data<=-16'd9262;
      10797:data<=16'd4167;
      10798:data<=16'd7639;
      10799:data<=16'd5902;
      10800:data<=16'd6343;
      10801:data<=16'd4040;
      10802:data<=16'd5077;
      10803:data<=16'd6000;
      10804:data<=16'd2359;
      10805:data<=16'd6053;
      10806:data<=16'd12496;
      10807:data<=16'd12531;
      10808:data<=16'd11734;
      10809:data<=16'd10154;
      10810:data<=16'd7571;
      10811:data<=16'd7283;
      10812:data<=16'd7653;
      10813:data<=16'd7254;
      10814:data<=16'd6067;
      10815:data<=16'd5627;
      10816:data<=16'd5448;
      10817:data<=16'd4002;
      10818:data<=16'd4096;
      10819:data<=16'd4131;
      10820:data<=16'd2954;
      10821:data<=16'd3797;
      10822:data<=16'd3798;
      10823:data<=16'd2810;
      10824:data<=16'd2679;
      10825:data<=16'd1262;
      10826:data<=16'd1528;
      10827:data<=16'd2449;
      10828:data<=16'd449;
      10829:data<=16'd334;
      10830:data<=16'd1820;
      10831:data<=16'd864;
      10832:data<=-16'd948;
      10833:data<=-16'd1331;
      10834:data<=-16'd613;
      10835:data<=-16'd2437;
      10836:data<=-16'd3906;
      10837:data<=-16'd1058;
      10838:data<=-16'd986;
      10839:data<=-16'd1902;
      10840:data<=16'd133;
      10841:data<=-16'd5263;
      10842:data<=-16'd15732;
      10843:data<=-16'd19870;
      10844:data<=-16'd19273;
      10845:data<=-16'd17400;
      10846:data<=-16'd16641;
      10847:data<=-16'd17429;
      10848:data<=-16'd16325;
      10849:data<=-16'd14293;
      10850:data<=-16'd13060;
      10851:data<=-16'd13876;
      10852:data<=-16'd15496;
      10853:data<=-16'd12871;
      10854:data<=-16'd11101;
      10855:data<=-16'd14383;
      10856:data<=-16'd14129;
      10857:data<=-16'd10455;
      10858:data<=-16'd11556;
      10859:data<=-16'd16554;
      10860:data<=-16'd19811;
      10861:data<=-16'd19353;
      10862:data<=-16'd17776;
      10863:data<=-16'd17139;
      10864:data<=-16'd16719;
      10865:data<=-16'd15095;
      10866:data<=-16'd12387;
      10867:data<=-16'd12648;
      10868:data<=-16'd15045;
      10869:data<=-16'd14210;
      10870:data<=-16'd12518;
      10871:data<=-16'd12301;
      10872:data<=-16'd12472;
      10873:data<=-16'd12649;
      10874:data<=-16'd9805;
      10875:data<=-16'd7517;
      10876:data<=-16'd9401;
      10877:data<=-16'd8592;
      10878:data<=-16'd5515;
      10879:data<=-16'd4679;
      10880:data<=-16'd4952;
      10881:data<=-16'd6307;
      10882:data<=-16'd5354;
      10883:data<=-16'd3791;
      10884:data<=-16'd5752;
      10885:data<=-16'd651;
      10886:data<=16'd11985;
      10887:data<=16'd17638;
      10888:data<=16'd16756;
      10889:data<=16'd16242;
      10890:data<=16'd16389;
      10891:data<=16'd16325;
      10892:data<=16'd15691;
      10893:data<=16'd16449;
      10894:data<=16'd17531;
      10895:data<=16'd16493;
      10896:data<=16'd15364;
      10897:data<=16'd14839;
      10898:data<=16'd15192;
      10899:data<=16'd14759;
      10900:data<=16'd12390;
      10901:data<=16'd13740;
      10902:data<=16'd15760;
      10903:data<=16'd13320;
      10904:data<=16'd13538;
      10905:data<=16'd15097;
      10906:data<=16'd13103;
      10907:data<=16'd12539;
      10908:data<=16'd12974;
      10909:data<=16'd12370;
      10910:data<=16'd12907;
      10911:data<=16'd15799;
      10912:data<=16'd20961;
      10913:data<=16'd22058;
      10914:data<=16'd18774;
      10915:data<=16'd18697;
      10916:data<=16'd19252;
      10917:data<=16'd19405;
      10918:data<=16'd20579;
      10919:data<=16'd18442;
      10920:data<=16'd17682;
      10921:data<=16'd19150;
      10922:data<=16'd16727;
      10923:data<=16'd15367;
      10924:data<=16'd14683;
      10925:data<=16'd12944;
      10926:data<=16'd15822;
      10927:data<=16'd16600;
      10928:data<=16'd14577;
      10929:data<=16'd16777;
      10930:data<=16'd11597;
      10931:data<=-16'd1513;
      10932:data<=-16'd5495;
      10933:data<=-16'd2335;
      10934:data<=-16'd1306;
      10935:data<=-16'd1021;
      10936:data<=-16'd315;
      10937:data<=-16'd509;
      10938:data<=-16'd1757;
      10939:data<=-16'd1903;
      10940:data<=-16'd481;
      10941:data<=-16'd607;
      10942:data<=-16'd1706;
      10943:data<=-16'd1148;
      10944:data<=16'd226;
      10945:data<=16'd872;
      10946:data<=16'd895;
      10947:data<=16'd1066;
      10948:data<=16'd1069;
      10949:data<=16'd1186;
      10950:data<=16'd2118;
      10951:data<=16'd2673;
      10952:data<=16'd3284;
      10953:data<=16'd4021;
      10954:data<=16'd3516;
      10955:data<=16'd3485;
      10956:data<=16'd3527;
      10957:data<=16'd2729;
      10958:data<=16'd3098;
      10959:data<=16'd3212;
      10960:data<=16'd3539;
      10961:data<=16'd4908;
      10962:data<=16'd3876;
      10963:data<=16'd2878;
      10964:data<=16'd1938;
      10965:data<=-16'd2881;
      10966:data<=-16'd5735;
      10967:data<=-16'd4632;
      10968:data<=-16'd3304;
      10969:data<=-16'd1118;
      10970:data<=-16'd1046;
      10971:data<=-16'd2420;
      10972:data<=-16'd2570;
      10973:data<=-16'd4455;
      10974:data<=-16'd987;
      10975:data<=16'd10249;
      10976:data<=16'd15969;
      10977:data<=16'd16070;
      10978:data<=16'd17135;
      10979:data<=16'd15773;
      10980:data<=16'd13201;
      10981:data<=16'd13681;
      10982:data<=16'd14575;
      10983:data<=16'd12683;
      10984:data<=16'd11314;
      10985:data<=16'd13206;
      10986:data<=16'd13159;
      10987:data<=16'd11433;
      10988:data<=16'd12328;
      10989:data<=16'd11136;
      10990:data<=16'd8915;
      10991:data<=16'd10216;
      10992:data<=16'd9996;
      10993:data<=16'd8737;
      10994:data<=16'd9938;
      10995:data<=16'd10508;
      10996:data<=16'd9835;
      10997:data<=16'd8851;
      10998:data<=16'd8787;
      10999:data<=16'd8787;
      11000:data<=16'd5958;
      11001:data<=16'd5814;
      11002:data<=16'd8916;
      11003:data<=16'd7497;
      11004:data<=16'd5465;
      11005:data<=16'd6590;
      11006:data<=16'd6575;
      11007:data<=16'd5623;
      11008:data<=16'd4379;
      11009:data<=16'd3284;
      11010:data<=16'd2914;
      11011:data<=16'd2176;
      11012:data<=16'd2319;
      11013:data<=16'd1448;
      11014:data<=16'd690;
      11015:data<=16'd3324;
      11016:data<=16'd2105;
      11017:data<=16'd1754;
      11018:data<=16'd9691;
      11019:data<=16'd6845;
      11020:data<=-16'd8235;
      11021:data<=-16'd12751;
      11022:data<=-16'd10084;
      11023:data<=-16'd10654;
      11024:data<=-16'd10170;
      11025:data<=-16'd9727;
      11026:data<=-16'd10960;
      11027:data<=-16'd11723;
      11028:data<=-16'd11958;
      11029:data<=-16'd11550;
      11030:data<=-16'd11997;
      11031:data<=-16'd12193;
      11032:data<=-16'd10255;
      11033:data<=-16'd9740;
      11034:data<=-16'd10674;
      11035:data<=-16'd10402;
      11036:data<=-16'd10410;
      11037:data<=-16'd11462;
      11038:data<=-16'd12102;
      11039:data<=-16'd11304;
      11040:data<=-16'd10724;
      11041:data<=-16'd11488;
      11042:data<=-16'd11292;
      11043:data<=-16'd11013;
      11044:data<=-16'd11652;
      11045:data<=-16'd11324;
      11046:data<=-16'd11276;
      11047:data<=-16'd10751;
      11048:data<=-16'd9236;
      11049:data<=-16'd10122;
      11050:data<=-16'd11107;
      11051:data<=-16'd10702;
      11052:data<=-16'd11309;
      11053:data<=-16'd10978;
      11054:data<=-16'd10229;
      11055:data<=-16'd10117;
      11056:data<=-16'd8921;
      11057:data<=-16'd8687;
      11058:data<=-16'd8628;
      11059:data<=-16'd7497;
      11060:data<=-16'd8075;
      11061:data<=-16'd8984;
      11062:data<=-16'd10232;
      11063:data<=-16'd10164;
      11064:data<=-16'd1895;
      11065:data<=16'd8011;
      11066:data<=16'd9673;
      11067:data<=16'd7912;
      11068:data<=16'd6683;
      11069:data<=16'd4983;
      11070:data<=16'd2743;
      11071:data<=-16'd1365;
      11072:data<=-16'd4508;
      11073:data<=-16'd4197;
      11074:data<=-16'd4168;
      11075:data<=-16'd4529;
      11076:data<=-16'd3965;
      11077:data<=-16'd5228;
      11078:data<=-16'd6896;
      11079:data<=-16'd6243;
      11080:data<=-16'd5694;
      11081:data<=-16'd6170;
      11082:data<=-16'd6608;
      11083:data<=-16'd6748;
      11084:data<=-16'd5325;
      11085:data<=-16'd4598;
      11086:data<=-16'd6532;
      11087:data<=-16'd6868;
      11088:data<=-16'd5739;
      11089:data<=-16'd6038;
      11090:data<=-16'd5915;
      11091:data<=-16'd6328;
      11092:data<=-16'd7257;
      11093:data<=-16'd6649;
      11094:data<=-16'd7121;
      11095:data<=-16'd7166;
      11096:data<=-16'd6002;
      11097:data<=-16'd7542;
      11098:data<=-16'd7530;
      11099:data<=-16'd5429;
      11100:data<=-16'd6378;
      11101:data<=-16'd6472;
      11102:data<=-16'd6129;
      11103:data<=-16'd7565;
      11104:data<=-16'd6328;
      11105:data<=-16'd6443;
      11106:data<=-16'd8035;
      11107:data<=-16'd5629;
      11108:data<=-16'd8986;
      11109:data<=-16'd19766;
      11110:data<=-16'd24518;
      11111:data<=-16'd23987;
      11112:data<=-16'd23914;
      11113:data<=-16'd22927;
      11114:data<=-16'd22049;
      11115:data<=-16'd21516;
      11116:data<=-16'd20800;
      11117:data<=-16'd20204;
      11118:data<=-16'd18478;
      11119:data<=-16'd17911;
      11120:data<=-16'd18812;
      11121:data<=-16'd17453;
      11122:data<=-16'd16210;
      11123:data<=-16'd15570;
      11124:data<=-16'd11113;
      11125:data<=-16'd6091;
      11126:data<=-16'd4670;
      11127:data<=-16'd5127;
      11128:data<=-16'd6431;
      11129:data<=-16'd6610;
      11130:data<=-16'd4868;
      11131:data<=-16'd4520;
      11132:data<=-16'd4931;
      11133:data<=-16'd3905;
      11134:data<=-16'd3518;
      11135:data<=-16'd4423;
      11136:data<=-16'd5116;
      11137:data<=-16'd5001;
      11138:data<=-16'd3917;
      11139:data<=-16'd3168;
      11140:data<=-16'd3742;
      11141:data<=-16'd4258;
      11142:data<=-16'd3835;
      11143:data<=-16'd2869;
      11144:data<=-16'd1941;
      11145:data<=-16'd1979;
      11146:data<=-16'd2115;
      11147:data<=-16'd726;
      11148:data<=-16'd132;
      11149:data<=-16'd866;
      11150:data<=16'd494;
      11151:data<=16'd378;
      11152:data<=-16'd1723;
      11153:data<=16'd5257;
      11154:data<=16'd17631;
      11155:data<=16'd20662;
      11156:data<=16'd18287;
      11157:data<=16'd18236;
      11158:data<=16'd17687;
      11159:data<=16'd16824;
      11160:data<=16'd17192;
      11161:data<=16'd18114;
      11162:data<=16'd18639;
      11163:data<=16'd17312;
      11164:data<=16'd16542;
      11165:data<=16'd16769;
      11166:data<=16'd15352;
      11167:data<=16'd14941;
      11168:data<=16'd15832;
      11169:data<=16'd15488;
      11170:data<=16'd15544;
      11171:data<=16'd15746;
      11172:data<=16'd15755;
      11173:data<=16'd16187;
      11174:data<=16'd14784;
      11175:data<=16'd13473;
      11176:data<=16'd13826;
      11177:data<=16'd10991;
      11178:data<=16'd5844;
      11179:data<=16'd4420;
      11180:data<=16'd5803;
      11181:data<=16'd5756;
      11182:data<=16'd4852;
      11183:data<=16'd4931;
      11184:data<=16'd4949;
      11185:data<=16'd5036;
      11186:data<=16'd6317;
      11187:data<=16'd7404;
      11188:data<=16'd6901;
      11189:data<=16'd5567;
      11190:data<=16'd5656;
      11191:data<=16'd6282;
      11192:data<=16'd4711;
      11193:data<=16'd4570;
      11194:data<=16'd6663;
      11195:data<=16'd6755;
      11196:data<=16'd7398;
      11197:data<=16'd5137;
      11198:data<=-16'd5172;
      11199:data<=-16'd11259;
      11200:data<=-16'd9476;
      11201:data<=-16'd10249;
      11202:data<=-16'd10470;
      11203:data<=-16'd7177;
      11204:data<=-16'd6414;
      11205:data<=-16'd6658;
      11206:data<=-16'd5606;
      11207:data<=-16'd5404;
      11208:data<=-16'd5444;
      11209:data<=-16'd4545;
      11210:data<=-16'd3351;
      11211:data<=-16'd2901;
      11212:data<=-16'd2382;
      11213:data<=-16'd1081;
      11214:data<=-16'd928;
      11215:data<=-16'd1259;
      11216:data<=-16'd444;
      11217:data<=-16'd411;
      11218:data<=-16'd1013;
      11219:data<=-16'd86;
      11220:data<=16'd1419;
      11221:data<=16'd1754;
      11222:data<=16'd1295;
      11223:data<=16'd1068;
      11224:data<=16'd1078;
      11225:data<=16'd763;
      11226:data<=16'd246;
      11227:data<=16'd1428;
      11228:data<=16'd3579;
      11229:data<=16'd3075;
      11230:data<=16'd4860;
      11231:data<=16'd11894;
      11232:data<=16'd13640;
      11233:data<=16'd10957;
      11234:data<=16'd12161;
      11235:data<=16'd11994;
      11236:data<=16'd11153;
      11237:data<=16'd12487;
      11238:data<=16'd10895;
      11239:data<=16'd11624;
      11240:data<=16'd13127;
      11241:data<=16'd9069;
      11242:data<=16'd13345;
      11243:data<=16'd25185;
      11244:data<=16'd27499;
      11245:data<=16'd25334;
      11246:data<=16'd25169;
      11247:data<=16'd23575;
      11248:data<=16'd22868;
      11249:data<=16'd22826;
      11250:data<=16'd21931;
      11251:data<=16'd20836;
      11252:data<=16'd19226;
      11253:data<=16'd19153;
      11254:data<=16'd19375;
      11255:data<=16'd18334;
      11256:data<=16'd18269;
      11257:data<=16'd17851;
      11258:data<=16'd17327;
      11259:data<=16'd17082;
      11260:data<=16'd14686;
      11261:data<=16'd13826;
      11262:data<=16'd15326;
      11263:data<=16'd14707;
      11264:data<=16'd13336;
      11265:data<=16'd12518;
      11266:data<=16'd11941;
      11267:data<=16'd12113;
      11268:data<=16'd11538;
      11269:data<=16'd11174;
      11270:data<=16'd11743;
      11271:data<=16'd11300;
      11272:data<=16'd10552;
      11273:data<=16'd10067;
      11274:data<=16'd9204;
      11275:data<=16'd8349;
      11276:data<=16'd8099;
      11277:data<=16'd8041;
      11278:data<=16'd6672;
      11279:data<=16'd5636;
      11280:data<=16'd5532;
      11281:data<=16'd4519;
      11282:data<=16'd4954;
      11283:data<=16'd2749;
      11284:data<=-16'd4845;
      11285:data<=-16'd6455;
      11286:data<=-16'd6391;
      11287:data<=-16'd16983;
      11288:data<=-16'd26172;
      11289:data<=-16'd25602;
      11290:data<=-16'd23532;
      11291:data<=-16'd22623;
      11292:data<=-16'd21925;
      11293:data<=-16'd20914;
      11294:data<=-16'd20879;
      11295:data<=-16'd22154;
      11296:data<=-16'd20688;
      11297:data<=-16'd20110;
      11298:data<=-16'd21547;
      11299:data<=-16'd18848;
      11300:data<=-16'd17396;
      11301:data<=-16'd19014;
      11302:data<=-16'd18023;
      11303:data<=-16'd18242;
      11304:data<=-16'd19183;
      11305:data<=-16'd18031;
      11306:data<=-16'd17594;
      11307:data<=-16'd16198;
      11308:data<=-16'd15588;
      11309:data<=-16'd16603;
      11310:data<=-16'd14718;
      11311:data<=-16'd14038;
      11312:data<=-16'd15547;
      11313:data<=-16'd15085;
      11314:data<=-16'd14760;
      11315:data<=-16'd13900;
      11316:data<=-16'd12922;
      11317:data<=-16'd13383;
      11318:data<=-16'd12164;
      11319:data<=-16'd12043;
      11320:data<=-16'd13520;
      11321:data<=-16'd12885;
      11322:data<=-16'd12845;
      11323:data<=-16'd12463;
      11324:data<=-16'd10915;
      11325:data<=-16'd10473;
      11326:data<=-16'd9157;
      11327:data<=-16'd9471;
      11328:data<=-16'd10496;
      11329:data<=-16'd8904;
      11330:data<=-16'd9888;
      11331:data<=-16'd6385;
      11332:data<=16'd5982;
      11333:data<=16'd10900;
      11334:data<=16'd8466;
      11335:data<=16'd8916;
      11336:data<=16'd8895;
      11337:data<=16'd9903;
      11338:data<=16'd12740;
      11339:data<=16'd12367;
      11340:data<=16'd11236;
      11341:data<=16'd10533;
      11342:data<=16'd9753;
      11343:data<=16'd10369;
      11344:data<=16'd9579;
      11345:data<=16'd7239;
      11346:data<=16'd6108;
      11347:data<=16'd5789;
      11348:data<=16'd5607;
      11349:data<=16'd5015;
      11350:data<=16'd4617;
      11351:data<=16'd4705;
      11352:data<=16'd3955;
      11353:data<=16'd3084;
      11354:data<=16'd2285;
      11355:data<=16'd1544;
      11356:data<=16'd1754;
      11357:data<=16'd1645;
      11358:data<=16'd1720;
      11359:data<=16'd2529;
      11360:data<=16'd2255;
      11361:data<=16'd1536;
      11362:data<=16'd535;
      11363:data<=-16'd428;
      11364:data<=-16'd258;
      11365:data<=-16'd1075;
      11366:data<=-16'd1833;
      11367:data<=-16'd1021;
      11368:data<=-16'd1095;
      11369:data<=-16'd1553;
      11370:data<=-16'd2921;
      11371:data<=-16'd4552;
      11372:data<=-16'd3312;
      11373:data<=-16'd3579;
      11374:data<=-16'd4387;
      11375:data<=-16'd2322;
      11376:data<=-16'd7905;
      11377:data<=-16'd19120;
      11378:data<=-16'd21391;
      11379:data<=-16'd19417;
      11380:data<=-16'd20337;
      11381:data<=-16'd19814;
      11382:data<=-16'd18090;
      11383:data<=-16'd17479;
      11384:data<=-16'd17309;
      11385:data<=-16'd16674;
      11386:data<=-16'd15590;
      11387:data<=-16'd15766;
      11388:data<=-16'd16001;
      11389:data<=-16'd15894;
      11390:data<=-16'd18524;
      11391:data<=-16'd21270;
      11392:data<=-16'd20883;
      11393:data<=-16'd19672;
      11394:data<=-16'd18648;
      11395:data<=-16'd17929;
      11396:data<=-16'd17855;
      11397:data<=-16'd17318;
      11398:data<=-16'd16145;
      11399:data<=-16'd15141;
      11400:data<=-16'd15101;
      11401:data<=-16'd14777;
      11402:data<=-16'd12903;
      11403:data<=-16'd12534;
      11404:data<=-16'd13831;
      11405:data<=-16'd13271;
      11406:data<=-16'd11997;
      11407:data<=-16'd11386;
      11408:data<=-16'd10718;
      11409:data<=-16'd10751;
      11410:data<=-16'd10592;
      11411:data<=-16'd8972;
      11412:data<=-16'd7542;
      11413:data<=-16'd7313;
      11414:data<=-16'd6693;
      11415:data<=-16'd5777;
      11416:data<=-16'd6102;
      11417:data<=-16'd4777;
      11418:data<=-16'd2772;
      11419:data<=-16'd4869;
      11420:data<=-16'd1579;
      11421:data<=16'd11723;
      11422:data<=16'd18812;
      11423:data<=16'd16798;
      11424:data<=16'd16213;
      11425:data<=16'd16372;
      11426:data<=16'd16042;
      11427:data<=16'd15517;
      11428:data<=16'd14327;
      11429:data<=16'd15396;
      11430:data<=16'd15854;
      11431:data<=16'd14634;
      11432:data<=16'd15020;
      11433:data<=16'd14034;
      11434:data<=16'd13470;
      11435:data<=16'd14909;
      11436:data<=16'd13744;
      11437:data<=16'd13725;
      11438:data<=16'd15180;
      11439:data<=16'd13940;
      11440:data<=16'd14029;
      11441:data<=16'd13788;
      11442:data<=16'd12217;
      11443:data<=16'd15009;
      11444:data<=16'd18255;
      11445:data<=16'd19127;
      11446:data<=16'd19807;
      11447:data<=16'd18528;
      11448:data<=16'd17878;
      11449:data<=16'd18856;
      11450:data<=16'd17992;
      11451:data<=16'd16577;
      11452:data<=16'd15300;
      11453:data<=16'd14612;
      11454:data<=16'd15600;
      11455:data<=16'd16029;
      11456:data<=16'd15309;
      11457:data<=16'd14126;
      11458:data<=16'd13650;
      11459:data<=16'd13715;
      11460:data<=16'd12057;
      11461:data<=16'd11867;
      11462:data<=16'd12878;
      11463:data<=16'd12323;
      11464:data<=16'd14004;
      11465:data<=16'd9732;
      11466:data<=-16'd3870;
      11467:data<=-16'd7887;
      11468:data<=-16'd3758;
      11469:data<=-16'd5500;
      11470:data<=-16'd5724;
      11471:data<=-16'd2696;
      11472:data<=-16'd2590;
      11473:data<=-16'd1897;
      11474:data<=-16'd1036;
      11475:data<=-16'd1550;
      11476:data<=-16'd1700;
      11477:data<=-16'd2666;
      11478:data<=-16'd2520;
      11479:data<=-16'd368;
      11480:data<=16'd549;
      11481:data<=16'd520;
      11482:data<=16'd508;
      11483:data<=16'd509;
      11484:data<=16'd1125;
      11485:data<=16'd1293;
      11486:data<=16'd951;
      11487:data<=16'd1885;
      11488:data<=16'd3312;
      11489:data<=16'd2837;
      11490:data<=16'd1577;
      11491:data<=16'd1835;
      11492:data<=16'd2182;
      11493:data<=16'd1263;
      11494:data<=16'd696;
      11495:data<=16'd1623;
      11496:data<=16'd1650;
      11497:data<=-16'd1762;
      11498:data<=-16'd4399;
      11499:data<=-16'd3544;
      11500:data<=-16'd3501;
      11501:data<=-16'd3577;
      11502:data<=-16'd2302;
      11503:data<=-16'd1935;
      11504:data<=-16'd1072;
      11505:data<=-16'd813;
      11506:data<=-16'd531;
      11507:data<=16'd1970;
      11508:data<=16'd450;
      11509:data<=16'd459;
      11510:data<=16'd10655;
      11511:data<=16'd17722;
      11512:data<=16'd17253;
      11513:data<=16'd17949;
      11514:data<=16'd16792;
      11515:data<=16'd14398;
      11516:data<=16'd14895;
      11517:data<=16'd15085;
      11518:data<=16'd14240;
      11519:data<=16'd13059;
      11520:data<=16'd12898;
      11521:data<=16'd13764;
      11522:data<=16'd12790;
      11523:data<=16'd12395;
      11524:data<=16'd12217;
      11525:data<=16'd10219;
      11526:data<=16'd10611;
      11527:data<=16'd11303;
      11528:data<=16'd9881;
      11529:data<=16'd10091;
      11530:data<=16'd10545;
      11531:data<=16'd10090;
      11532:data<=16'd9497;
      11533:data<=16'd8669;
      11534:data<=16'd8822;
      11535:data<=16'd8106;
      11536:data<=16'd7333;
      11537:data<=16'd8123;
      11538:data<=16'd7594;
      11539:data<=16'd7718;
      11540:data<=16'd8008;
      11541:data<=16'd6029;
      11542:data<=16'd6002;
      11543:data<=16'd6217;
      11544:data<=16'd5195;
      11545:data<=16'd5535;
      11546:data<=16'd4520;
      11547:data<=16'd3753;
      11548:data<=16'd3386;
      11549:data<=16'd3142;
      11550:data<=16'd8216;
      11551:data<=16'd9597;
      11552:data<=16'd5823;
      11553:data<=16'd8388;
      11554:data<=16'd4038;
      11555:data<=-16'd10536;
      11556:data<=-16'd15098;
      11557:data<=-16'd13342;
      11558:data<=-16'd13832;
      11559:data<=-16'd12750;
      11560:data<=-16'd12869;
      11561:data<=-16'd13479;
      11562:data<=-16'd13396;
      11563:data<=-16'd14624;
      11564:data<=-16'd13806;
      11565:data<=-16'd12833;
      11566:data<=-16'd13494;
      11567:data<=-16'd12592;
      11568:data<=-16'd12043;
      11569:data<=-16'd11897;
      11570:data<=-16'd11321;
      11571:data<=-16'd12452;
      11572:data<=-16'd13376;
      11573:data<=-16'd13167;
      11574:data<=-16'd12783;
      11575:data<=-16'd12070;
      11576:data<=-16'd12172;
      11577:data<=-16'd11978;
      11578:data<=-16'd10930;
      11579:data<=-16'd11326;
      11580:data<=-16'd12469;
      11581:data<=-16'd12851;
      11582:data<=-16'd12968;
      11583:data<=-16'd13207;
      11584:data<=-16'd12648;
      11585:data<=-16'd11147;
      11586:data<=-16'd10948;
      11587:data<=-16'd11506;
      11588:data<=-16'd11500;
      11589:data<=-16'd12237;
      11590:data<=-16'd12104;
      11591:data<=-16'd11012;
      11592:data<=-16'd10784;
      11593:data<=-16'd9623;
      11594:data<=-16'd9364;
      11595:data<=-16'd10828;
      11596:data<=-16'd10278;
      11597:data<=-16'd10354;
      11598:data<=-16'd10346;
      11599:data<=-16'd3128;
      11600:data<=16'd6523;
      11601:data<=16'd8684;
      11602:data<=16'd4649;
      11603:data<=16'd842;
      11604:data<=-16'd1181;
      11605:data<=-16'd2631;
      11606:data<=-16'd2927;
      11607:data<=-16'd2534;
      11608:data<=-16'd2443;
      11609:data<=-16'd2049;
      11610:data<=-16'd2414;
      11611:data<=-16'd3066;
      11612:data<=-16'd2851;
      11613:data<=-16'd3921;
      11614:data<=-16'd5113;
      11615:data<=-16'd4954;
      11616:data<=-16'd5321;
      11617:data<=-16'd4996;
      11618:data<=-16'd4363;
      11619:data<=-16'd4884;
      11620:data<=-16'd4664;
      11621:data<=-16'd5154;
      11622:data<=-16'd6754;
      11623:data<=-16'd6849;
      11624:data<=-16'd6461;
      11625:data<=-16'd5732;
      11626:data<=-16'd5086;
      11627:data<=-16'd5338;
      11628:data<=-16'd4237;
      11629:data<=-16'd4347;
      11630:data<=-16'd6411;
      11631:data<=-16'd5903;
      11632:data<=-16'd5456;
      11633:data<=-16'd5829;
      11634:data<=-16'd4487;
      11635:data<=-16'd4511;
      11636:data<=-16'd4372;
      11637:data<=-16'd3780;
      11638:data<=-16'd5645;
      11639:data<=-16'd5479;
      11640:data<=-16'd5529;
      11641:data<=-16'd7086;
      11642:data<=-16'd4015;
      11643:data<=-16'd7403;
      11644:data<=-16'd19886;
      11645:data<=-16'd23017;
      11646:data<=-16'd20504;
      11647:data<=-16'd22301;
      11648:data<=-16'd21793;
      11649:data<=-16'd20518;
      11650:data<=-16'd20927;
      11651:data<=-16'd19608;
      11652:data<=-16'd18152;
      11653:data<=-16'd16759;
      11654:data<=-16'd16565;
      11655:data<=-16'd16140;
      11656:data<=-16'd11151;
      11657:data<=-16'd7881;
      11658:data<=-16'd8070;
      11659:data<=-16'd6889;
      11660:data<=-16'd7166;
      11661:data<=-16'd7209;
      11662:data<=-16'd6085;
      11663:data<=-16'd7629;
      11664:data<=-16'd7758;
      11665:data<=-16'd6719;
      11666:data<=-16'd7197;
      11667:data<=-16'd6351;
      11668:data<=-16'd6229;
      11669:data<=-16'd5858;
      11670:data<=-16'd3859;
      11671:data<=-16'd4939;
      11672:data<=-16'd6490;
      11673:data<=-16'd6234;
      11674:data<=-16'd5830;
      11675:data<=-16'd4243;
      11676:data<=-16'd3902;
      11677:data<=-16'd4106;
      11678:data<=-16'd3486;
      11679:data<=-16'd4168;
      11680:data<=-16'd2843;
      11681:data<=-16'd1591;
      11682:data<=-16'd2513;
      11683:data<=-16'd910;
      11684:data<=-16'd804;
      11685:data<=-16'd1169;
      11686:data<=16'd388;
      11687:data<=-16'd1607;
      11688:data<=16'd4472;
      11689:data<=16'd19112;
      11690:data<=16'd21416;
      11691:data<=16'd17663;
      11692:data<=16'd18898;
      11693:data<=16'd18659;
      11694:data<=16'd18545;
      11695:data<=16'd18415;
      11696:data<=16'd17364;
      11697:data<=16'd18927;
      11698:data<=16'd18204;
      11699:data<=16'd16410;
      11700:data<=16'd17326;
      11701:data<=16'd16768;
      11702:data<=16'd16227;
      11703:data<=16'd16019;
      11704:data<=16'd15253;
      11705:data<=16'd16680;
      11706:data<=16'd16686;
      11707:data<=16'd15393;
      11708:data<=16'd14809;
      11709:data<=16'd10895;
      11710:data<=16'd7300;
      11711:data<=16'd7103;
      11712:data<=16'd6951;
      11713:data<=16'd8038;
      11714:data<=16'd9273;
      11715:data<=16'd8657;
      11716:data<=16'd8860;
      11717:data<=16'd9870;
      11718:data<=16'd9911;
      11719:data<=16'd8692;
      11720:data<=16'd8049;
      11721:data<=16'd9222;
      11722:data<=16'd9820;
      11723:data<=16'd9709;
      11724:data<=16'd9699;
      11725:data<=16'd9188;
      11726:data<=16'd9056;
      11727:data<=16'd8601;
      11728:data<=16'd8072;
      11729:data<=16'd8219;
      11730:data<=16'd8566;
      11731:data<=16'd10493;
      11732:data<=16'd7741;
      11733:data<=-16'd3280;
      11734:data<=-16'd9448;
      11735:data<=-16'd7603;
      11736:data<=-16'd6937;
      11737:data<=-16'd6875;
      11738:data<=-16'd5961;
      11739:data<=-16'd5354;
      11740:data<=-16'd4143;
      11741:data<=-16'd3345;
      11742:data<=-16'd2475;
      11743:data<=-16'd1601;
      11744:data<=-16'd1724;
      11745:data<=-16'd930;
      11746:data<=16'd376;
      11747:data<=16'd1357;
      11748:data<=16'd2008;
      11749:data<=16'd1369;
      11750:data<=16'd1351;
      11751:data<=16'd1986;
      11752:data<=16'd1759;
      11753:data<=16'd2065;
      11754:data<=16'd2478;
      11755:data<=16'd3274;
      11756:data<=16'd5012;
      11757:data<=16'd5316;
      11758:data<=16'd4648;
      11759:data<=16'd4153;
      11760:data<=16'd3773;
      11761:data<=16'd4187;
      11762:data<=16'd5744;
      11763:data<=16'd9793;
      11764:data<=16'd13073;
      11765:data<=16'd12081;
      11766:data<=16'd11558;
      11767:data<=16'd11335;
      11768:data<=16'd9662;
      11769:data<=16'd10088;
      11770:data<=16'd9673;
      11771:data<=16'd8990;
      11772:data<=16'd11003;
      11773:data<=16'd10144;
      11774:data<=16'd9514;
      11775:data<=16'd10904;
      11776:data<=16'd8533;
      11777:data<=16'd12490;
      11778:data<=16'd23877;
      11779:data<=16'd26207;
      11780:data<=16'd23913;
      11781:data<=16'd25780;
      11782:data<=16'd25240;
      11783:data<=16'd23323;
      11784:data<=16'd23309;
      11785:data<=16'd21919;
      11786:data<=16'd19973;
      11787:data<=16'd18551;
      11788:data<=16'd17561;
      11789:data<=16'd18063;
      11790:data<=16'd17958;
      11791:data<=16'd16416;
      11792:data<=16'd15411;
      11793:data<=16'd14901;
      11794:data<=16'd14801;
      11795:data<=16'd14759;
      11796:data<=16'd13784;
      11797:data<=16'd13221;
      11798:data<=16'd13321;
      11799:data<=16'd12748;
      11800:data<=16'd12148;
      11801:data<=16'd11226;
      11802:data<=16'd10014;
      11803:data<=16'd10137;
      11804:data<=16'd9941;
      11805:data<=16'd9477;
      11806:data<=16'd10865;
      11807:data<=16'd10699;
      11808:data<=16'd8877;
      11809:data<=16'd9219;
      11810:data<=16'd8837;
      11811:data<=16'd7124;
      11812:data<=16'd7001;
      11813:data<=16'd6742;
      11814:data<=16'd6470;
      11815:data<=16'd4711;
      11816:data<=-16'd798;
      11817:data<=-16'd3063;
      11818:data<=-16'd1682;
      11819:data<=-16'd2908;
      11820:data<=-16'd2543;
      11821:data<=-16'd3488;
      11822:data<=-16'd13737;
      11823:data<=-16'd22571;
      11824:data<=-16'd22360;
      11825:data<=-16'd21328;
      11826:data<=-16'd21472;
      11827:data<=-16'd20613;
      11828:data<=-16'd20007;
      11829:data<=-16'd19414;
      11830:data<=-16'd19581;
      11831:data<=-16'd20256;
      11832:data<=-16'd19517;
      11833:data<=-16'd18803;
      11834:data<=-16'd18636;
      11835:data<=-16'd18160;
      11836:data<=-16'd17892;
      11837:data<=-16'd17092;
      11838:data<=-16'd16553;
      11839:data<=-16'd17802;
      11840:data<=-16'd18442;
      11841:data<=-16'd17117;
      11842:data<=-16'd15876;
      11843:data<=-16'd15597;
      11844:data<=-16'd15277;
      11845:data<=-16'd14405;
      11846:data<=-16'd13999;
      11847:data<=-16'd14331;
      11848:data<=-16'd14509;
      11849:data<=-16'd14882;
      11850:data<=-16'd15477;
      11851:data<=-16'd15026;
      11852:data<=-16'd13781;
      11853:data<=-16'd13502;
      11854:data<=-16'd14095;
      11855:data<=-16'd13902;
      11856:data<=-16'd13541;
      11857:data<=-16'd13702;
      11858:data<=-16'd13320;
      11859:data<=-16'd13135;
      11860:data<=-16'd12731;
      11861:data<=-16'd11444;
      11862:data<=-16'd11408;
      11863:data<=-16'd11321;
      11864:data<=-16'd11486;
      11865:data<=-16'd13333;
      11866:data<=-16'd8731;
      11867:data<=16'd2443;
      11868:data<=16'd8898;
      11869:data<=16'd11248;
      11870:data<=16'd12797;
      11871:data<=16'd11538;
      11872:data<=16'd10493;
      11873:data<=16'd9941;
      11874:data<=16'd8169;
      11875:data<=16'd7180;
      11876:data<=16'd6492;
      11877:data<=16'd6179;
      11878:data<=16'd6191;
      11879:data<=16'd4968;
      11880:data<=16'd4015;
      11881:data<=16'd2972;
      11882:data<=16'd1776;
      11883:data<=16'd1959;
      11884:data<=16'd1585;
      11885:data<=16'd1612;
      11886:data<=16'd2370;
      11887:data<=16'd1233;
      11888:data<=16'd610;
      11889:data<=16'd26;
      11890:data<=-16'd2035;
      11891:data<=-16'd2088;
      11892:data<=-16'd1509;
      11893:data<=-16'd1545;
      11894:data<=-16'd779;
      11895:data<=-16'd793;
      11896:data<=-16'd776;
      11897:data<=-16'd1340;
      11898:data<=-16'd3036;
      11899:data<=-16'd2804;
      11900:data<=-16'd2864;
      11901:data<=-16'd3354;
      11902:data<=-16'd2690;
      11903:data<=-16'd3806;
      11904:data<=-16'd3548;
      11905:data<=-16'd2720;
      11906:data<=-16'd5456;
      11907:data<=-16'd5564;
      11908:data<=-16'd4711;
      11909:data<=-16'd5742;
      11910:data<=-16'd4084;
      11911:data<=-16'd9044;
      11912:data<=-16'd20372;
      11913:data<=-16'd22222;
      11914:data<=-16'd20058;
      11915:data<=-16'd21761;
      11916:data<=-16'd21053;
      11917:data<=-16'd19490;
      11918:data<=-16'd19506;
      11919:data<=-16'd18265;
      11920:data<=-16'd16795;
      11921:data<=-16'd17461;
      11922:data<=-16'd20892;
      11923:data<=-16'd23385;
      11924:data<=-16'd22272;
      11925:data<=-16'd21041;
      11926:data<=-16'd20556;
      11927:data<=-16'd19825;
      11928:data<=-16'd19221;
      11929:data<=-16'd17644;
      11930:data<=-16'd16657;
      11931:data<=-16'd17478;
      11932:data<=-16'd17362;
      11933:data<=-16'd16117;
      11934:data<=-16'd15262;
      11935:data<=-16'd14422;
      11936:data<=-16'd13421;
      11937:data<=-16'd12913;
      11938:data<=-16'd12825;
      11939:data<=-16'd12928;
      11940:data<=-16'd13797;
      11941:data<=-16'd13937;
      11942:data<=-16'd12484;
      11943:data<=-16'd11693;
      11944:data<=-16'd10830;
      11945:data<=-16'd9817;
      11946:data<=-16'd10040;
      11947:data<=-16'd8769;
      11948:data<=-16'd7515;
      11949:data<=-16'd7862;
      11950:data<=-16'd6457;
      11951:data<=-16'd5832;
      11952:data<=-16'd5404;
      11953:data<=-16'd3621;
      11954:data<=-16'd5665;
      11955:data<=-16'd2461;
      11956:data<=16'd10881;
      11957:data<=16'd17086;
      11958:data<=16'd15377;
      11959:data<=16'd16042;
      11960:data<=16'd15505;
      11961:data<=16'd14627;
      11962:data<=16'd15065;
      11963:data<=16'd13917;
      11964:data<=16'd14436;
      11965:data<=16'd15324;
      11966:data<=16'd14142;
      11967:data<=16'd14298;
      11968:data<=16'd14236;
      11969:data<=16'd12815;
      11970:data<=16'd12425;
      11971:data<=16'd12935;
      11972:data<=16'd13635;
      11973:data<=16'd13550;
      11974:data<=16'd14580;
      11975:data<=16'd17760;
      11976:data<=16'd18733;
      11977:data<=16'd18045;
      11978:data<=16'd17623;
      11979:data<=16'd16358;
      11980:data<=16'd16923;
      11981:data<=16'd18472;
      11982:data<=16'd18181;
      11983:data<=16'd17970;
      11984:data<=16'd17265;
      11985:data<=16'd16175;
      11986:data<=16'd16057;
      11987:data<=16'd15394;
      11988:data<=16'd15309;
      11989:data<=16'd15823;
      11990:data<=16'd15808;
      11991:data<=16'd16034;
      11992:data<=16'd14640;
      11993:data<=16'd13306;
      11994:data<=16'd13690;
      11995:data<=16'd12800;
      11996:data<=16'd12839;
      11997:data<=16'd13044;
      11998:data<=16'd12037;
      11999:data<=16'd13853;
      12000:data<=16'd9653;
      12001:data<=-16'd2834;
      12002:data<=-16'd7130;
      12003:data<=-16'd4901;
      12004:data<=-16'd5444;
      12005:data<=-16'd4250;
      12006:data<=-16'd2672;
      12007:data<=-16'd2874;
      12008:data<=-16'd1804;
      12009:data<=-16'd1347;
      12010:data<=-16'd1350;
      12011:data<=-16'd839;
      12012:data<=-16'd1136;
      12013:data<=-16'd1118;
      12014:data<=-16'd365;
      12015:data<=16'd1295;
      12016:data<=16'd2312;
      12017:data<=16'd1092;
      12018:data<=16'd1665;
      12019:data<=16'd3920;
      12020:data<=16'd4381;
      12021:data<=16'd4399;
      12022:data<=16'd4469;
      12023:data<=16'd5103;
      12024:data<=16'd5864;
      12025:data<=16'd4854;
      12026:data<=16'd4569;
      12027:data<=16'd3698;
      12028:data<=-16'd226;
      12029:data<=-16'd2629;
      12030:data<=-16'd2519;
      12031:data<=-16'd1582;
      12032:data<=-16'd543;
      12033:data<=-16'd1021;
      12034:data<=-16'd541;
      12035:data<=16'd505;
      12036:data<=-16'd453;
      12037:data<=-16'd570;
      12038:data<=-16'd177;
      12039:data<=16'd29;
      12040:data<=16'd1324;
      12041:data<=16'd1792;
      12042:data<=16'd2302;
      12043:data<=16'd2235;
      12044:data<=16'd2880;
      12045:data<=16'd10351;
      12046:data<=16'd16732;
      12047:data<=16'd15678;
      12048:data<=16'd16061;
      12049:data<=16'd17095;
      12050:data<=16'd15625;
      12051:data<=16'd15368;
      12052:data<=16'd14181;
      12053:data<=16'd12828;
      12054:data<=16'd12747;
      12055:data<=16'd11230;
      12056:data<=16'd11626;
      12057:data<=16'd13537;
      12058:data<=16'd12898;
      12059:data<=16'd12102;
      12060:data<=16'd11499;
      12061:data<=16'd10577;
      12062:data<=16'd10361;
      12063:data<=16'd9456;
      12064:data<=16'd8866;
      12065:data<=16'd9400;
      12066:data<=16'd9817;
      12067:data<=16'd9987;
      12068:data<=16'd8915;
      12069:data<=16'd7580;
      12070:data<=16'd7374;
      12071:data<=16'd6912;
      12072:data<=16'd6912;
      12073:data<=16'd7896;
      12074:data<=16'd8345;
      12075:data<=16'd7993;
      12076:data<=16'd7224;
      12077:data<=16'd6866;
      12078:data<=16'd6751;
      12079:data<=16'd6314;
      12080:data<=16'd6038;
      12081:data<=16'd6670;
      12082:data<=16'd9609;
      12083:data<=16'd11285;
      12084:data<=16'd9000;
      12085:data<=16'd8933;
      12086:data<=16'd9636;
      12087:data<=16'd7527;
      12088:data<=16'd7771;
      12089:data<=16'd3688;
      12090:data<=-16'd7615;
      12091:data<=-16'd11627;
      12092:data<=-16'd10261;
      12093:data<=-16'd11814;
      12094:data<=-16'd11112;
      12095:data<=-16'd9988;
      12096:data<=-16'd10583;
      12097:data<=-16'd9417;
      12098:data<=-16'd9949;
      12099:data<=-16'd11405;
      12100:data<=-16'd10595;
      12101:data<=-16'd10662;
      12102:data<=-16'd10671;
      12103:data<=-16'd9565;
      12104:data<=-16'd9740;
      12105:data<=-16'd10119;
      12106:data<=-16'd10511;
      12107:data<=-16'd11594;
      12108:data<=-16'd11767;
      12109:data<=-16'd10900;
      12110:data<=-16'd10097;
      12111:data<=-16'd10005;
      12112:data<=-16'd10050;
      12113:data<=-16'd9583;
      12114:data<=-16'd9870;
      12115:data<=-16'd10851;
      12116:data<=-16'd11432;
      12117:data<=-16'd11894;
      12118:data<=-16'd11731;
      12119:data<=-16'd10892;
      12120:data<=-16'd10222;
      12121:data<=-16'd9530;
      12122:data<=-16'd9379;
      12123:data<=-16'd10246;
      12124:data<=-16'd11082;
      12125:data<=-16'd11239;
      12126:data<=-16'd10533;
      12127:data<=-16'd9210;
      12128:data<=-16'd8557;
      12129:data<=-16'd9051;
      12130:data<=-16'd9379;
      12131:data<=-16'd9417;
      12132:data<=-16'd10648;
      12133:data<=-16'd10634;
      12134:data<=-16'd6120;
      12135:data<=-16'd1431;
      12136:data<=-16'd1013;
      12137:data<=-16'd1683;
      12138:data<=-16'd1145;
      12139:data<=-16'd1676;
      12140:data<=-16'd3463;
      12141:data<=-16'd4228;
      12142:data<=-16'd4070;
      12143:data<=-16'd4238;
      12144:data<=-16'd4164;
      12145:data<=-16'd3918;
      12146:data<=-16'd3765;
      12147:data<=-16'd3330;
      12148:data<=-16'd4482;
      12149:data<=-16'd6495;
      12150:data<=-16'd6137;
      12151:data<=-16'd5418;
      12152:data<=-16'd5618;
      12153:data<=-16'd5065;
      12154:data<=-16'd4949;
      12155:data<=-16'd5092;
      12156:data<=-16'd5328;
      12157:data<=-16'd6611;
      12158:data<=-16'd6593;
      12159:data<=-16'd6231;
      12160:data<=-16'd6904;
      12161:data<=-16'd5671;
      12162:data<=-16'd4287;
      12163:data<=-16'd4040;
      12164:data<=-16'd3294;
      12165:data<=-16'd4168;
      12166:data<=-16'd5365;
      12167:data<=-16'd5473;
      12168:data<=-16'd6441;
      12169:data<=-16'd6093;
      12170:data<=-16'd5118;
      12171:data<=-16'd5150;
      12172:data<=-16'd4222;
      12173:data<=-16'd4637;
      12174:data<=-16'd5632;
      12175:data<=-16'd5501;
      12176:data<=-16'd6425;
      12177:data<=-16'd5134;
      12178:data<=-16'd6655;
      12179:data<=-16'd16651;
      12180:data<=-16'd21270;
      12181:data<=-16'd18497;
      12182:data<=-16'd19312;
      12183:data<=-16'd19503;
      12184:data<=-16'd17606;
      12185:data<=-16'd17761;
      12186:data<=-16'd16818;
      12187:data<=-16'd13775;
      12188:data<=-16'd9242;
      12189:data<=-16'd6378;
      12190:data<=-16'd7891;
      12191:data<=-16'd8323;
      12192:data<=-16'd7235;
      12193:data<=-16'd6924;
      12194:data<=-16'd5783;
      12195:data<=-16'd6261;
      12196:data<=-16'd6802;
      12197:data<=-16'd5281;
      12198:data<=-16'd5285;
      12199:data<=-16'd5204;
      12200:data<=-16'd4975;
      12201:data<=-16'd5626;
      12202:data<=-16'd4087;
      12203:data<=-16'd3610;
      12204:data<=-16'd4394;
      12205:data<=-16'd3018;
      12206:data<=-16'd3447;
      12207:data<=-16'd5212;
      12208:data<=-16'd5454;
      12209:data<=-16'd5336;
      12210:data<=-16'd4470;
      12211:data<=-16'd4097;
      12212:data<=-16'd3585;
      12213:data<=-16'd2428;
      12214:data<=-16'd2834;
      12215:data<=-16'd1855;
      12216:data<=-16'd875;
      12217:data<=-16'd2012;
      12218:data<=-16'd1300;
      12219:data<=-16'd1754;
      12220:data<=-16'd1760;
      12221:data<=16'd904;
      12222:data<=-16'd707;
      12223:data<=16'd3366;
      12224:data<=16'd16321;
      12225:data<=16'd19285;
      12226:data<=16'd16463;
      12227:data<=16'd17444;
      12228:data<=16'd15547;
      12229:data<=16'd14877;
      12230:data<=16'd15955;
      12231:data<=16'd13891;
      12232:data<=16'd14930;
      12233:data<=16'd16712;
      12234:data<=16'd14947;
      12235:data<=16'd14910;
      12236:data<=16'd15079;
      12237:data<=16'd13565;
      12238:data<=16'd13468;
      12239:data<=16'd13403;
      12240:data<=16'd11338;
      12241:data<=16'd8886;
      12242:data<=16'd8279;
      12243:data<=16'd8005;
      12244:data<=16'd6546;
      12245:data<=16'd6555;
      12246:data<=16'd6939;
      12247:data<=16'd5927;
      12248:data<=16'd6576;
      12249:data<=16'd8078;
      12250:data<=16'd8416;
      12251:data<=16'd9148;
      12252:data<=16'd9542;
      12253:data<=16'd8587;
      12254:data<=16'd7929;
      12255:data<=16'd7653;
      12256:data<=16'd6778;
      12257:data<=16'd7063;
      12258:data<=16'd8617;
      12259:data<=16'd8605;
      12260:data<=16'd8549;
      12261:data<=16'd8812;
      12262:data<=16'd7345;
      12263:data<=16'd7749;
      12264:data<=16'd8508;
      12265:data<=16'd7327;
      12266:data<=16'd9712;
      12267:data<=16'd8727;
      12268:data<=-16'd1139;
      12269:data<=-16'd6579;
      12270:data<=-16'd5333;
      12271:data<=-16'd4854;
      12272:data<=-16'd4381;
      12273:data<=-16'd4253;
      12274:data<=-16'd3617;
      12275:data<=-16'd1991;
      12276:data<=-16'd2375;
      12277:data<=-16'd2381;
      12278:data<=-16'd1475;
      12279:data<=-16'd1407;
      12280:data<=-16'd1169;
      12281:data<=-16'd1644;
      12282:data<=-16'd617;
      12283:data<=16'd1918;
      12284:data<=16'd1729;
      12285:data<=16'd1404;
      12286:data<=16'd1682;
      12287:data<=16'd1544;
      12288:data<=16'd2717;
      12289:data<=16'd2217;
      12290:data<=16'd2273;
      12291:data<=16'd4667;
      12292:data<=16'd3707;
      12293:data<=16'd4572;
      12294:data<=16'd9265;
      12295:data<=16'd9494;
      12296:data<=16'd8432;
      12297:data<=16'd8752;
      12298:data<=16'd7970;
      12299:data<=16'd8846;
      12300:data<=16'd9802;
      12301:data<=16'd9658;
      12302:data<=16'd9879;
      12303:data<=16'd8940;
      12304:data<=16'd8796;
      12305:data<=16'd8566;
      12306:data<=16'd7225;
      12307:data<=16'd8771;
      12308:data<=16'd9796;
      12309:data<=16'd9298;
      12310:data<=16'd9615;
      12311:data<=16'd7702;
      12312:data<=16'd11353;
      12313:data<=16'd21672;
      12314:data<=16'd23457;
      12315:data<=16'd20886;
      12316:data<=16'd22351;
      12317:data<=16'd21165;
      12318:data<=16'd19943;
      12319:data<=16'd20619;
      12320:data<=16'd18381;
      12321:data<=16'd17344;
      12322:data<=16'd17135;
      12323:data<=16'd14833;
      12324:data<=16'd14862;
      12325:data<=16'd15547;
      12326:data<=16'd14698;
      12327:data<=16'd14877;
      12328:data<=16'd14158;
      12329:data<=16'd12586;
      12330:data<=16'd12222;
      12331:data<=16'd11402;
      12332:data<=16'd10555;
      12333:data<=16'd10690;
      12334:data<=16'd10680;
      12335:data<=16'd10261;
      12336:data<=16'd9815;
      12337:data<=16'd9972;
      12338:data<=16'd9664;
      12339:data<=16'd8076;
      12340:data<=16'd7978;
      12341:data<=16'd9450;
      12342:data<=16'd9404;
      12343:data<=16'd8117;
      12344:data<=16'd7598;
      12345:data<=16'd7652;
      12346:data<=16'd6072;
      12347:data<=16'd2572;
      12348:data<=-16'd284;
      12349:data<=-16'd1453;
      12350:data<=-16'd1589;
      12351:data<=-16'd1917;
      12352:data<=-16'd2681;
      12353:data<=-16'd2640;
      12354:data<=-16'd2908;
      12355:data<=-16'd2913;
      12356:data<=-16'd3095;
      12357:data<=-16'd10452;
      12358:data<=-16'd20139;
      12359:data<=-16'd20817;
      12360:data<=-16'd19049;
      12361:data<=-16'd20063;
      12362:data<=-16'd18763;
      12363:data<=-16'd17831;
      12364:data<=-16'd18343;
      12365:data<=-16'd17801;
      12366:data<=-16'd18501;
      12367:data<=-16'd18765;
      12368:data<=-16'd17491;
      12369:data<=-16'd17030;
      12370:data<=-16'd16196;
      12371:data<=-16'd15850;
      12372:data<=-16'd16020;
      12373:data<=-16'd14662;
      12374:data<=-16'd14880;
      12375:data<=-16'd16330;
      12376:data<=-16'd15673;
      12377:data<=-16'd14985;
      12378:data<=-16'd14418;
      12379:data<=-16'd13021;
      12380:data<=-16'd12965;
      12381:data<=-16'd13649;
      12382:data<=-16'd14032;
      12383:data<=-16'd14748;
      12384:data<=-16'd14815;
      12385:data<=-16'd14734;
      12386:data<=-16'd15183;
      12387:data<=-16'd14258;
      12388:data<=-16'd12927;
      12389:data<=-16'd12698;
      12390:data<=-16'd12245;
      12391:data<=-16'd12972;
      12392:data<=-16'd14328;
      12393:data<=-16'd13191;
      12394:data<=-16'd12592;
      12395:data<=-16'd12754;
      12396:data<=-16'd11256;
      12397:data<=-16'd11250;
      12398:data<=-16'd10662;
      12399:data<=-16'd9418;
      12400:data<=-16'd10561;
      12401:data<=-16'd3941;
      12402:data<=16'd8105;
      12403:data<=16'd10151;
      12404:data<=16'd8516;
      12405:data<=16'd9317;
      12406:data<=16'd7941;
      12407:data<=16'd7946;
      12408:data<=16'd7310;
      12409:data<=16'd4575;
      12410:data<=16'd5143;
      12411:data<=16'd5015;
      12412:data<=16'd3545;
      12413:data<=16'd3850;
      12414:data<=16'd3515;
      12415:data<=16'd3805;
      12416:data<=16'd2754;
      12417:data<=16'd99;
      12418:data<=16'd816;
      12419:data<=16'd453;
      12420:data<=-16'd1151;
      12421:data<=-16'd234;
      12422:data<=-16'd852;
      12423:data<=-16'd1092;
      12424:data<=-16'd1017;
      12425:data<=-16'd3374;
      12426:data<=-16'd2760;
      12427:data<=-16'd1641;
      12428:data<=-16'd2628;
      12429:data<=-16'd1771;
      12430:data<=-16'd2097;
      12431:data<=-16'd2511;
      12432:data<=-16'd1491;
      12433:data<=-16'd2957;
      12434:data<=-16'd3805;
      12435:data<=-16'd3988;
      12436:data<=-16'd4611;
      12437:data<=-16'd3077;
      12438:data<=-16'd3582;
      12439:data<=-16'd4713;
      12440:data<=-16'd3836;
      12441:data<=-16'd5374;
      12442:data<=-16'd5864;
      12443:data<=-16'd5583;
      12444:data<=-16'd6777;
      12445:data<=-16'd4737;
      12446:data<=-16'd8170;
      12447:data<=-16'd18616;
      12448:data<=-16'd20750;
      12449:data<=-16'd18842;
      12450:data<=-16'd20876;
      12451:data<=-16'd20196;
      12452:data<=-16'd18512;
      12453:data<=-16'd20416;
      12454:data<=-16'd22852;
      12455:data<=-16'd23062;
      12456:data<=-16'd21018;
      12457:data<=-16'd19773;
      12458:data<=-16'd20137;
      12459:data<=-16'd19851;
      12460:data<=-16'd19550;
      12461:data<=-16'd19458;
      12462:data<=-16'd18707;
      12463:data<=-16'd17699;
      12464:data<=-16'd16604;
      12465:data<=-16'd15599;
      12466:data<=-16'd14727;
      12467:data<=-16'd14612;
      12468:data<=-16'd15124;
      12469:data<=-16'd14530;
      12470:data<=-16'd13573;
      12471:data<=-16'd13136;
      12472:data<=-16'd12260;
      12473:data<=-16'd11442;
      12474:data<=-16'd11591;
      12475:data<=-16'd12745;
      12476:data<=-16'd12930;
      12477:data<=-16'd11156;
      12478:data<=-16'd10243;
      12479:data<=-16'd9844;
      12480:data<=-16'd8793;
      12481:data<=-16'd8701;
      12482:data<=-16'd7999;
      12483:data<=-16'd6695;
      12484:data<=-16'd5985;
      12485:data<=-16'd4658;
      12486:data<=-16'd4940;
      12487:data<=-16'd5354;
      12488:data<=-16'd3664;
      12489:data<=-16'd4246;
      12490:data<=-16'd1626;
      12491:data<=16'd8762;
      12492:data<=16'd14997;
      12493:data<=16'd14277;
      12494:data<=16'd14252;
      12495:data<=16'd14542;
      12496:data<=16'd14325;
      12497:data<=16'd14305;
      12498:data<=16'd13449;
      12499:data<=16'd13224;
      12500:data<=16'd14415;
      12501:data<=16'd15067;
      12502:data<=16'd14401;
      12503:data<=16'd14170;
      12504:data<=16'd14233;
      12505:data<=16'd13174;
      12506:data<=16'd14477;
      12507:data<=16'd18292;
      12508:data<=16'd19676;
      12509:data<=16'd19948;
      12510:data<=16'd19904;
      12511:data<=16'd18346;
      12512:data<=16'd18081;
      12513:data<=16'd17650;
      12514:data<=16'd16199;
      12515:data<=16'd16480;
      12516:data<=16'd16480;
      12517:data<=16'd16557;
      12518:data<=16'd17722;
      12519:data<=16'd17476;
      12520:data<=16'd17391;
      12521:data<=16'd17229;
      12522:data<=16'd15876;
      12523:data<=16'd15241;
      12524:data<=16'd14169;
      12525:data<=16'd14507;
      12526:data<=16'd16210;
      12527:data<=16'd14869;
      12528:data<=16'd14346;
      12529:data<=16'd14361;
      12530:data<=16'd12151;
      12531:data<=16'd12992;
      12532:data<=16'd12944;
      12533:data<=16'd11917;
      12534:data<=16'd15790;
      12535:data<=16'd11383;
      12536:data<=-16'd1239;
      12537:data<=-16'd3868;
      12538:data<=-16'd1841;
      12539:data<=-16'd2905;
      12540:data<=-16'd1994;
      12541:data<=-16'd1119;
      12542:data<=-16'd414;
      12543:data<=16'd1130;
      12544:data<=16'd588;
      12545:data<=16'd164;
      12546:data<=16'd469;
      12547:data<=16'd599;
      12548:data<=16'd1086;
      12549:data<=16'd450;
      12550:data<=16'd1115;
      12551:data<=16'd3378;
      12552:data<=16'd3416;
      12553:data<=16'd2913;
      12554:data<=16'd2981;
      12555:data<=16'd3218;
      12556:data<=16'd3747;
      12557:data<=16'd3136;
      12558:data<=16'd3776;
      12559:data<=16'd3927;
      12560:data<=16'd6;
      12561:data<=-16'd1453;
      12562:data<=-16'd372;
      12563:data<=-16'd1859;
      12564:data<=-16'd2391;
      12565:data<=-16'd2261;
      12566:data<=-16'd2036;
      12567:data<=16'd502;
      12568:data<=16'd967;
      12569:data<=16'd89;
      12570:data<=16'd714;
      12571:data<=-16'd50;
      12572:data<=-16'd18;
      12573:data<=16'd1060;
      12574:data<=16'd478;
      12575:data<=16'd1259;
      12576:data<=16'd2990;
      12577:data<=16'd3284;
      12578:data<=16'd2585;
      12579:data<=16'd3547;
      12580:data<=16'd11198;
      12581:data<=16'd18679;
      12582:data<=16'd17273;
      12583:data<=16'd15838;
      12584:data<=16'd18002;
      12585:data<=16'd17697;
      12586:data<=16'd16845;
      12587:data<=16'd16031;
      12588:data<=16'd14578;
      12589:data<=16'd14948;
      12590:data<=16'd14678;
      12591:data<=16'd13302;
      12592:data<=16'd13412;
      12593:data<=16'd13565;
      12594:data<=16'd13490;
      12595:data<=16'd13673;
      12596:data<=16'd12897;
      12597:data<=16'd11605;
      12598:data<=16'd10686;
      12599:data<=16'd10248;
      12600:data<=16'd10249;
      12601:data<=16'd10390;
      12602:data<=16'd10154;
      12603:data<=16'd9665;
      12604:data<=16'd9730;
      12605:data<=16'd9473;
      12606:data<=16'd8511;
      12607:data<=16'd7896;
      12608:data<=16'd7664;
      12609:data<=16'd9072;
      12610:data<=16'd10398;
      12611:data<=16'd8522;
      12612:data<=16'd8426;
      12613:data<=16'd11870;
      12614:data<=16'd13465;
      12615:data<=16'd13030;
      12616:data<=16'd11781;
      12617:data<=16'd10709;
      12618:data<=16'd10621;
      12619:data<=16'd9441;
      12620:data<=16'd9380;
      12621:data<=16'd9803;
      12622:data<=16'd7985;
      12623:data<=16'd8458;
      12624:data<=16'd5109;
      12625:data<=-16'd6880;
      12626:data<=-16'd12466;
      12627:data<=-16'd10281;
      12628:data<=-16'd10830;
      12629:data<=-16'd10763;
      12630:data<=-16'd9881;
      12631:data<=-16'd10813;
      12632:data<=-16'd10137;
      12633:data<=-16'd10043;
      12634:data<=-16'd11512;
      12635:data<=-16'd11479;
      12636:data<=-16'd11136;
      12637:data<=-16'd10863;
      12638:data<=-16'd10270;
      12639:data<=-16'd10281;
      12640:data<=-16'd10251;
      12641:data<=-16'd10066;
      12642:data<=-16'd10542;
      12643:data<=-16'd11403;
      12644:data<=-16'd11351;
      12645:data<=-16'd10792;
      12646:data<=-16'd10912;
      12647:data<=-16'd10067;
      12648:data<=-16'd8856;
      12649:data<=-16'd9303;
      12650:data<=-16'd9858;
      12651:data<=-16'd10731;
      12652:data<=-16'd11649;
      12653:data<=-16'd11050;
      12654:data<=-16'd11025;
      12655:data<=-16'd10945;
      12656:data<=-16'd9956;
      12657:data<=-16'd9861;
      12658:data<=-16'd9306;
      12659:data<=-16'd9929;
      12660:data<=-16'd12093;
      12661:data<=-16'd11509;
      12662:data<=-16'd10890;
      12663:data<=-16'd11141;
      12664:data<=-16'd9855;
      12665:data<=-16'd10689;
      12666:data<=-16'd12854;
      12667:data<=-16'd15537;
      12668:data<=-16'd18342;
      12669:data<=-16'd11913;
      12670:data<=-16'd995;
      12671:data<=16'd638;
      12672:data<=-16'd1216;
      12673:data<=-16'd411;
      12674:data<=-16'd834;
      12675:data<=-16'd1759;
      12676:data<=-16'd2441;
      12677:data<=-16'd3054;
      12678:data<=-16'd2989;
      12679:data<=-16'd3450;
      12680:data<=-16'd3551;
      12681:data<=-16'd3112;
      12682:data<=-16'd2807;
      12683:data<=-16'd2156;
      12684:data<=-16'd3083;
      12685:data<=-16'd4772;
      12686:data<=-16'd4943;
      12687:data<=-16'd5147;
      12688:data<=-16'd5100;
      12689:data<=-16'd4672;
      12690:data<=-16'd4996;
      12691:data<=-16'd4911;
      12692:data<=-16'd5327;
      12693:data<=-16'd6537;
      12694:data<=-16'd6702;
      12695:data<=-16'd6443;
      12696:data<=-16'd5686;
      12697:data<=-16'd4754;
      12698:data<=-16'd4725;
      12699:data<=-16'd4382;
      12700:data<=-16'd4948;
      12701:data<=-16'd6827;
      12702:data<=-16'd6975;
      12703:data<=-16'd6288;
      12704:data<=-16'd6244;
      12705:data<=-16'd5644;
      12706:data<=-16'd4963;
      12707:data<=-16'd4869;
      12708:data<=-16'd4746;
      12709:data<=-16'd4766;
      12710:data<=-16'd6217;
      12711:data<=-16'd7060;
      12712:data<=-16'd4739;
      12713:data<=-16'd6760;
      12714:data<=-16'd16716;
      12715:data<=-16'd22052;
      12716:data<=-16'd19186;
      12717:data<=-16'd18550;
      12718:data<=-16'd20249;
      12719:data<=-16'd17528;
      12720:data<=-16'd12448;
      12721:data<=-16'd10410;
      12722:data<=-16'd10473;
      12723:data<=-16'd9700;
      12724:data<=-16'd8972;
      12725:data<=-16'd8758;
      12726:data<=-16'd8842;
      12727:data<=-16'd9553;
      12728:data<=-16'd9356;
      12729:data<=-16'd8878;
      12730:data<=-16'd8986;
      12731:data<=-16'd8041;
      12732:data<=-16'd7180;
      12733:data<=-16'd6579;
      12734:data<=-16'd6003;
      12735:data<=-16'd7185;
      12736:data<=-16'd7512;
      12737:data<=-16'd6790;
      12738:data<=-16'd7247;
      12739:data<=-16'd6410;
      12740:data<=-16'd5686;
      12741:data<=-16'd5923;
      12742:data<=-16'd4940;
      12743:data<=-16'd5864;
      12744:data<=-16'd6789;
      12745:data<=-16'd5143;
      12746:data<=-16'd5245;
      12747:data<=-16'd5154;
      12748:data<=-16'd4112;
      12749:data<=-16'd4896;
      12750:data<=-16'd4481;
      12751:data<=-16'd4172;
      12752:data<=-16'd4461;
      12753:data<=-16'd2572;
      12754:data<=-16'd2299;
      12755:data<=-16'd2129;
      12756:data<=-16'd1180;
      12757:data<=-16'd3371;
      12758:data<=16'd1347;
      12759:data<=16'd14296;
      12760:data<=16'd18592;
      12761:data<=16'd15503;
      12762:data<=16'd15434;
      12763:data<=16'd15434;
      12764:data<=16'd14472;
      12765:data<=16'd14537;
      12766:data<=16'd13486;
      12767:data<=16'd12975;
      12768:data<=16'd14672;
      12769:data<=16'd14603;
      12770:data<=16'd13262;
      12771:data<=16'd13781;
      12772:data<=16'd11835;
      12773:data<=16'd7148;
      12774:data<=16'd6082;
      12775:data<=16'd6739;
      12776:data<=16'd6708;
      12777:data<=16'd8087;
      12778:data<=16'd8204;
      12779:data<=16'd7181;
      12780:data<=16'd7309;
      12781:data<=16'd6540;
      12782:data<=16'd6102;
      12783:data<=16'd6733;
      12784:data<=16'd7118;
      12785:data<=16'd8608;
      12786:data<=16'd9051;
      12787:data<=16'd7990;
      12788:data<=16'd8264;
      12789:data<=16'd7661;
      12790:data<=16'd6564;
      12791:data<=16'd7304;
      12792:data<=16'd8003;
      12793:data<=16'd8425;
      12794:data<=16'd8437;
      12795:data<=16'd8437;
      12796:data<=16'd9232;
      12797:data<=16'd8407;
      12798:data<=16'd7638;
      12799:data<=16'd7585;
      12800:data<=16'd6519;
      12801:data<=16'd8969;
      12802:data<=16'd9277;
      12803:data<=-16'd331;
      12804:data<=-16'd7151;
      12805:data<=-16'd5732;
      12806:data<=-16'd5460;
      12807:data<=-16'd6034;
      12808:data<=-16'd5318;
      12809:data<=-16'd4352;
      12810:data<=-16'd2482;
      12811:data<=-16'd1841;
      12812:data<=-16'd2291;
      12813:data<=-16'd2237;
      12814:data<=-16'd2071;
      12815:data<=-16'd1236;
      12816:data<=-16'd1286;
      12817:data<=-16'd1689;
      12818:data<=-16'd202;
      12819:data<=16'd966;
      12820:data<=16'd1598;
      12821:data<=16'd1768;
      12822:data<=16'd990;
      12823:data<=16'd1651;
      12824:data<=16'd1762;
      12825:data<=16'd2491;
      12826:data<=16'd7641;
      12827:data<=16'd10513;
      12828:data<=16'd9373;
      12829:data<=16'd9024;
      12830:data<=16'd7764;
      12831:data<=16'd7201;
      12832:data<=16'd8002;
      12833:data<=16'd7112;
      12834:data<=16'd7750;
      12835:data<=16'd9268;
      12836:data<=16'd8802;
      12837:data<=16'd8663;
      12838:data<=16'd8084;
      12839:data<=16'd7388;
      12840:data<=16'd7826;
      12841:data<=16'd7497;
      12842:data<=16'd7239;
      12843:data<=16'd7383;
      12844:data<=16'd8293;
      12845:data<=16'd8901;
      12846:data<=16'd6307;
      12847:data<=16'd9386;
      12848:data<=16'd20093;
      12849:data<=16'd22999;
      12850:data<=16'd19669;
      12851:data<=16'd20149;
      12852:data<=16'd20118;
      12853:data<=16'd19118;
      12854:data<=16'd19199;
      12855:data<=16'd17757;
      12856:data<=16'd16724;
      12857:data<=16'd16026;
      12858:data<=16'd14195;
      12859:data<=16'd14131;
      12860:data<=16'd15173;
      12861:data<=16'd14882;
      12862:data<=16'd14449;
      12863:data<=16'd14504;
      12864:data<=16'd13632;
      12865:data<=16'd12222;
      12866:data<=16'd11661;
      12867:data<=16'd10727;
      12868:data<=16'd10354;
      12869:data<=16'd11825;
      12870:data<=16'd11277;
      12871:data<=16'd9591;
      12872:data<=16'd9565;
      12873:data<=16'd8611;
      12874:data<=16'd8167;
      12875:data<=16'd8408;
      12876:data<=16'd7435;
      12877:data<=16'd8567;
      12878:data<=16'd7877;
      12879:data<=16'd2692;
      12880:data<=16'd666;
      12881:data<=16'd643;
      12882:data<=-16'd397;
      12883:data<=-16'd52;
      12884:data<=-16'd796;
      12885:data<=-16'd1598;
      12886:data<=-16'd1237;
      12887:data<=-16'd2264;
      12888:data<=-16'd2100;
      12889:data<=-16'd2046;
      12890:data<=-16'd2887;
      12891:data<=-16'd2308;
      12892:data<=-16'd8166;
      12893:data<=-16'd18298;
      12894:data<=-16'd20040;
      12895:data<=-16'd18255;
      12896:data<=-16'd18906;
      12897:data<=-16'd18199;
      12898:data<=-16'd17399;
      12899:data<=-16'd16950;
      12900:data<=-16'd15940;
      12901:data<=-16'd16428;
      12902:data<=-16'd17297;
      12903:data<=-16'd17212;
      12904:data<=-16'd16979;
      12905:data<=-16'd16768;
      12906:data<=-16'd16393;
      12907:data<=-16'd15816;
      12908:data<=-16'd15487;
      12909:data<=-16'd15089;
      12910:data<=-16'd15094;
      12911:data<=-16'd15887;
      12912:data<=-16'd15412;
      12913:data<=-16'd14818;
      12914:data<=-16'd15089;
      12915:data<=-16'd14113;
      12916:data<=-16'd13441;
      12917:data<=-16'd13221;
      12918:data<=-16'd13018;
      12919:data<=-16'd14789;
      12920:data<=-16'd15323;
      12921:data<=-16'd14377;
      12922:data<=-16'd14716;
      12923:data<=-16'd13759;
      12924:data<=-16'd12771;
      12925:data<=-16'd12568;
      12926:data<=-16'd11682;
      12927:data<=-16'd12783;
      12928:data<=-16'd13077;
      12929:data<=-16'd12084;
      12930:data<=-16'd12941;
      12931:data<=-16'd10504;
      12932:data<=-16'd6496;
      12933:data<=-16'd4825;
      12934:data<=-16'd3556;
      12935:data<=-16'd6196;
      12936:data<=-16'd5037;
      12937:data<=16'd5583;
      12938:data<=16'd9724;
      12939:data<=16'd7359;
      12940:data<=16'd8373;
      12941:data<=16'd7971;
      12942:data<=16'd7403;
      12943:data<=16'd7362;
      12944:data<=16'd4353;
      12945:data<=16'd3717;
      12946:data<=16'd4472;
      12947:data<=16'd3491;
      12948:data<=16'd3482;
      12949:data<=16'd3134;
      12950:data<=16'd3131;
      12951:data<=16'd3156;
      12952:data<=16'd925;
      12953:data<=16'd188;
      12954:data<=16'd422;
      12955:data<=-16'd329;
      12956:data<=-16'd97;
      12957:data<=-16'd406;
      12958:data<=-16'd365;
      12959:data<=16'd519;
      12960:data<=-16'd940;
      12961:data<=-16'd2669;
      12962:data<=-16'd3143;
      12963:data<=-16'd2776;
      12964:data<=-16'd1105;
      12965:data<=-16'd766;
      12966:data<=-16'd1045;
      12967:data<=-16'd346;
      12968:data<=-16'd1334;
      12969:data<=-16'd2981;
      12970:data<=-16'd3181;
      12971:data<=-16'd2531;
      12972:data<=-16'd1974;
      12973:data<=-16'd2416;
      12974:data<=-16'd2347;
      12975:data<=-16'd2155;
      12976:data<=-16'd3106;
      12977:data<=-16'd3295;
      12978:data<=-16'd4337;
      12979:data<=-16'd4937;
      12980:data<=-16'd2494;
      12981:data<=-16'd6670;
      12982:data<=-16'd17623;
      12983:data<=-16'd20101;
      12984:data<=-16'd16815;
      12985:data<=-16'd19892;
      12986:data<=-16'd24371;
      12987:data<=-16'd24069;
      12988:data<=-16'd22660;
      12989:data<=-16'd21420;
      12990:data<=-16'd19923;
      12991:data<=-16'd19349;
      12992:data<=-16'd18389;
      12993:data<=-16'd17559;
      12994:data<=-16'd18403;
      12995:data<=-16'd18368;
      12996:data<=-16'd17749;
      12997:data<=-16'd17641;
      12998:data<=-16'd15995;
      12999:data<=-16'd15054;
      13000:data<=-16'd14910;
      13001:data<=-16'd12822;
      13002:data<=-16'd12584;
      13003:data<=-16'd13731;
      13004:data<=-16'd12533;
      13005:data<=-16'd11838;
      13006:data<=-16'd11436;
      13007:data<=-16'd10313;
      13008:data<=-16'd10143;
      13009:data<=-16'd9279;
      13010:data<=-16'd9313;
      13011:data<=-16'd10957;
      13012:data<=-16'd10241;
      13013:data<=-16'd8959;
      13014:data<=-16'd8573;
      13015:data<=-16'd7726;
      13016:data<=-16'd7694;
      13017:data<=-16'd7233;
      13018:data<=-16'd6396;
      13019:data<=-16'd6363;
      13020:data<=-16'd5362;
      13021:data<=-16'd4951;
      13022:data<=-16'd4514;
      13023:data<=-16'd3139;
      13024:data<=-16'd4419;
      13025:data<=-16'd2006;
      13026:data<=16'd7853;
      13027:data<=16'd13750;
      13028:data<=16'd13849;
      13029:data<=16'd14458;
      13030:data<=16'd14304;
      13031:data<=16'd13600;
      13032:data<=16'd13787;
      13033:data<=16'd13315;
      13034:data<=16'd12801;
      13035:data<=16'd13564;
      13036:data<=16'd14542;
      13037:data<=16'd14554;
      13038:data<=16'd16387;
      13039:data<=16'd20421;
      13040:data<=16'd20800;
      13041:data<=16'd18903;
      13042:data<=16'd19103;
      13043:data<=16'd18707;
      13044:data<=16'd18615;
      13045:data<=16'd19716;
      13046:data<=16'd19124;
      13047:data<=16'd18751;
      13048:data<=16'd18456;
      13049:data<=16'd17185;
      13050:data<=16'd17021;
      13051:data<=16'd16425;
      13052:data<=16'd16495;
      13053:data<=16'd18225;
      13054:data<=16'd18078;
      13055:data<=16'd17819;
      13056:data<=16'd17798;
      13057:data<=16'd16569;
      13058:data<=16'd16486;
      13059:data<=16'd15402;
      13060:data<=16'd14753;
      13061:data<=16'd17011;
      13062:data<=16'd16581;
      13063:data<=16'd15606;
      13064:data<=16'd15963;
      13065:data<=16'd14035;
      13066:data<=16'd14346;
      13067:data<=16'd14105;
      13068:data<=16'd11609;
      13069:data<=16'd14800;
      13070:data<=16'd12709;
      13071:data<=16'd1095;
      13072:data<=-16'd2027;
      13073:data<=16'd452;
      13074:data<=-16'd986;
      13075:data<=-16'd655;
      13076:data<=16'd211;
      13077:data<=16'd350;
      13078:data<=16'd2093;
      13079:data<=16'd2146;
      13080:data<=16'd1809;
      13081:data<=16'd2516;
      13082:data<=16'd2012;
      13083:data<=16'd1820;
      13084:data<=16'd2135;
      13085:data<=16'd2475;
      13086:data<=16'd3800;
      13087:data<=16'd4646;
      13088:data<=16'd4235;
      13089:data<=16'd3811;
      13090:data<=16'd4366;
      13091:data<=16'd3218;
      13092:data<=-16'd1735;
      13093:data<=-16'd3876;
      13094:data<=-16'd1101;
      13095:data<=-16'd180;
      13096:data<=-16'd511;
      13097:data<=16'd115;
      13098:data<=-16'd741;
      13099:data<=-16'd1512;
      13100:data<=-16'd1198;
      13101:data<=-16'd1316;
      13102:data<=-16'd657;
      13103:data<=16'd904;
      13104:data<=16'd1245;
      13105:data<=16'd643;
      13106:data<=16'd1058;
      13107:data<=16'd1394;
      13108:data<=16'd790;
      13109:data<=16'd1538;
      13110:data<=16'd2326;
      13111:data<=16'd2469;
      13112:data<=16'd3915;
      13113:data<=16'd3401;
      13114:data<=16'd3648;
      13115:data<=16'd10989;
      13116:data<=16'd17572;
      13117:data<=16'd17423;
      13118:data<=16'd16119;
      13119:data<=16'd16128;
      13120:data<=16'd16759;
      13121:data<=16'd16627;
      13122:data<=16'd15437;
      13123:data<=16'd15306;
      13124:data<=16'd14882;
      13125:data<=16'd13503;
      13126:data<=16'd12433;
      13127:data<=16'd11711;
      13128:data<=16'd12671;
      13129:data<=16'd13018;
      13130:data<=16'd11532;
      13131:data<=16'd11702;
      13132:data<=16'd11723;
      13133:data<=16'd10960;
      13134:data<=16'd10745;
      13135:data<=16'd9163;
      13136:data<=16'd9221;
      13137:data<=16'd10454;
      13138:data<=16'd9360;
      13139:data<=16'd9266;
      13140:data<=16'd8783;
      13141:data<=16'd7579;
      13142:data<=16'd8511;
      13143:data<=16'd7618;
      13144:data<=16'd8875;
      13145:data<=16'd14593;
      13146:data<=16'd15383;
      13147:data<=16'd13417;
      13148:data<=16'd13074;
      13149:data<=16'd11875;
      13150:data<=16'd11611;
      13151:data<=16'd10869;
      13152:data<=16'd9809;
      13153:data<=16'd9966;
      13154:data<=16'd8126;
      13155:data<=16'd7670;
      13156:data<=16'd7708;
      13157:data<=16'd5733;
      13158:data<=16'd7568;
      13159:data<=16'd4278;
      13160:data<=-16'd7608;
      13161:data<=-16'd11688;
      13162:data<=-16'd10709;
      13163:data<=-16'd12765;
      13164:data<=-16'd12187;
      13165:data<=-16'd11317;
      13166:data<=-16'd11913;
      13167:data<=-16'd11392;
      13168:data<=-16'd11805;
      13169:data<=-16'd12022;
      13170:data<=-16'd12110;
      13171:data<=-16'd12889;
      13172:data<=-16'd12434;
      13173:data<=-16'd12214;
      13174:data<=-16'd12070;
      13175:data<=-16'd11376;
      13176:data<=-16'd11232;
      13177:data<=-16'd11057;
      13178:data<=-16'd12339;
      13179:data<=-16'd13270;
      13180:data<=-16'd11963;
      13181:data<=-16'd12167;
      13182:data<=-16'd12017;
      13183:data<=-16'd10877;
      13184:data<=-16'd11700;
      13185:data<=-16'd11547;
      13186:data<=-16'd11817;
      13187:data<=-16'd13673;
      13188:data<=-16'd13705;
      13189:data<=-16'd13831;
      13190:data<=-16'd13197;
      13191:data<=-16'd12185;
      13192:data<=-16'd13367;
      13193:data<=-16'd11793;
      13194:data<=-16'd10863;
      13195:data<=-16'd13291;
      13196:data<=-16'd11908;
      13197:data<=-16'd12775;
      13198:data<=-16'd17514;
      13199:data<=-16'd17347;
      13200:data<=-16'd16932;
      13201:data<=-16'd16577;
      13202:data<=-16'd14912;
      13203:data<=-16'd17350;
      13204:data<=-16'd13506;
      13205:data<=-16'd2279;
      13206:data<=16'd306;
      13207:data<=-16'd1612;
      13208:data<=-16'd864;
      13209:data<=-16'd1538;
      13210:data<=-16'd1427;
      13211:data<=-16'd1312;
      13212:data<=-16'd3474;
      13213:data<=-16'd4097;
      13214:data<=-16'd3789;
      13215:data<=-16'd3650;
      13216:data<=-16'd3071;
      13217:data<=-16'd3265;
      13218:data<=-16'd3086;
      13219:data<=-16'd3163;
      13220:data<=-16'd4743;
      13221:data<=-16'd5033;
      13222:data<=-16'd4094;
      13223:data<=-16'd3905;
      13224:data<=-16'd4187;
      13225:data<=-16'd4608;
      13226:data<=-16'd4325;
      13227:data<=-16'd3717;
      13228:data<=-16'd4488;
      13229:data<=-16'd5683;
      13230:data<=-16'd5855;
      13231:data<=-16'd5301;
      13232:data<=-16'd4249;
      13233:data<=-16'd3463;
      13234:data<=-16'd3695;
      13235:data<=-16'd3894;
      13236:data<=-16'd4337;
      13237:data<=-16'd6023;
      13238:data<=-16'd6347;
      13239:data<=-16'd5325;
      13240:data<=-16'd5768;
      13241:data<=-16'd5218;
      13242:data<=-16'd4058;
      13243:data<=-16'd5031;
      13244:data<=-16'd4886;
      13245:data<=-16'd5498;
      13246:data<=-16'd7329;
      13247:data<=-16'd4545;
      13248:data<=-16'd6451;
      13249:data<=-16'd17450;
      13250:data<=-16'd20698;
      13251:data<=-16'd15065;
      13252:data<=-16'd12302;
      13253:data<=-16'd12013;
      13254:data<=-16'd12851;
      13255:data<=-16'd13521;
      13256:data<=-16'd12125;
      13257:data<=-16'd11746;
      13258:data<=-16'd11271;
      13259:data<=-16'd9740;
      13260:data<=-16'd9674;
      13261:data<=-16'd9683;
      13262:data<=-16'd10207;
      13263:data<=-16'd11453;
      13264:data<=-16'd10684;
      13265:data<=-16'd9580;
      13266:data<=-16'd9646;
      13267:data<=-16'd9683;
      13268:data<=-16'd8775;
      13269:data<=-16'd7339;
      13270:data<=-16'd8204;
      13271:data<=-16'd9374;
      13272:data<=-16'd8131;
      13273:data<=-16'd7937;
      13274:data<=-16'd8260;
      13275:data<=-16'd7758;
      13276:data<=-16'd7840;
      13277:data<=-16'd6811;
      13278:data<=-16'd6733;
      13279:data<=-16'd8385;
      13280:data<=-16'd7993;
      13281:data<=-16'd7457;
      13282:data<=-16'd6866;
      13283:data<=-16'd5322;
      13284:data<=-16'd5594;
      13285:data<=-16'd5112;
      13286:data<=-16'd3994;
      13287:data<=-16'd4262;
      13288:data<=-16'd3055;
      13289:data<=-16'd2682;
      13290:data<=-16'd2742;
      13291:data<=-16'd1721;
      13292:data<=-16'd3539;
      13293:data<=16'd402;
      13294:data<=16'd11987;
      13295:data<=16'd15556;
      13296:data<=16'd14076;
      13297:data<=16'd15773;
      13298:data<=16'd14651;
      13299:data<=16'd13406;
      13300:data<=16'd14854;
      13301:data<=16'd13740;
      13302:data<=16'd12443;
      13303:data<=16'd12671;
      13304:data<=16'd10781;
      13305:data<=16'd8181;
      13306:data<=16'd8002;
      13307:data<=16'd8619;
      13308:data<=16'd7818;
      13309:data<=16'd7558;
      13310:data<=16'd8069;
      13311:data<=16'd7790;
      13312:data<=16'd8704;
      13313:data<=16'd9533;
      13314:data<=16'd8777;
      13315:data<=16'd9289;
      13316:data<=16'd9385;
      13317:data<=16'd8408;
      13318:data<=16'd8528;
      13319:data<=16'd8160;
      13320:data<=16'd8934;
      13321:data<=16'd10921;
      13322:data<=16'd10425;
      13323:data<=16'd9882;
      13324:data<=16'd10134;
      13325:data<=16'd9517;
      13326:data<=16'd9226;
      13327:data<=16'd8472;
      13328:data<=16'd8654;
      13329:data<=16'd10342;
      13330:data<=16'd10006;
      13331:data<=16'd9062;
      13332:data<=16'd8957;
      13333:data<=16'd8910;
      13334:data<=16'd8819;
      13335:data<=16'd7454;
      13336:data<=16'd7921;
      13337:data<=16'd7932;
      13338:data<=16'd285;
      13339:data<=-16'd6234;
      13340:data<=-16'd5360;
      13341:data<=-16'd5215;
      13342:data<=-16'd5712;
      13343:data<=-16'd4854;
      13344:data<=-16'd4965;
      13345:data<=-16'd3850;
      13346:data<=-16'd2217;
      13347:data<=-16'd1521;
      13348:data<=-16'd740;
      13349:data<=-16'd1398;
      13350:data<=-16'd1917;
      13351:data<=-16'd1019;
      13352:data<=-16'd1336;
      13353:data<=-16'd1268;
      13354:data<=16'd749;
      13355:data<=16'd1256;
      13356:data<=-16'd9;
      13357:data<=16'd2103;
      13358:data<=16'd6930;
      13359:data<=16'd7547;
      13360:data<=16'd5661;
      13361:data<=16'd6331;
      13362:data<=16'd7206;
      13363:data<=16'd7686;
      13364:data<=16'd7941;
      13365:data<=16'd6478;
      13366:data<=16'd5865;
      13367:data<=16'd6235;
      13368:data<=16'd6100;
      13369:data<=16'd6190;
      13370:data<=16'd5949;
      13371:data<=16'd6871;
      13372:data<=16'd8199;
      13373:data<=16'd7345;
      13374:data<=16'd6860;
      13375:data<=16'd6382;
      13376:data<=16'd5800;
      13377:data<=16'd6839;
      13378:data<=16'd6398;
      13379:data<=16'd7181;
      13380:data<=16'd8805;
      13381:data<=16'd5838;
      13382:data<=16'd9116;
      13383:data<=16'd20089;
      13384:data<=16'd22651;
      13385:data<=16'd19948;
      13386:data<=16'd20024;
      13387:data<=16'd19575;
      13388:data<=16'd19977;
      13389:data<=16'd20262;
      13390:data<=16'd18105;
      13391:data<=16'd17129;
      13392:data<=16'd16988;
      13393:data<=16'd15985;
      13394:data<=16'd14850;
      13395:data<=16'd14722;
      13396:data<=16'd16098;
      13397:data<=16'd15716;
      13398:data<=16'd13988;
      13399:data<=16'd13913;
      13400:data<=16'd13283;
      13401:data<=16'd12308;
      13402:data<=16'd12038;
      13403:data<=16'd11130;
      13404:data<=16'd11097;
      13405:data<=16'd11508;
      13406:data<=16'd11145;
      13407:data<=16'd10701;
      13408:data<=16'd10038;
      13409:data<=16'd10477;
      13410:data<=16'd9333;
      13411:data<=16'd4901;
      13412:data<=16'd4153;
      13413:data<=16'd5979;
      13414:data<=16'd4895;
      13415:data<=16'd4469;
      13416:data<=16'd4639;
      13417:data<=16'd3418;
      13418:data<=16'd3093;
      13419:data<=16'd3090;
      13420:data<=16'd3130;
      13421:data<=16'd2634;
      13422:data<=16'd1113;
      13423:data<=16'd1251;
      13424:data<=16'd1301;
      13425:data<=16'd851;
      13426:data<=16'd1016;
      13427:data<=-16'd4857;
      13428:data<=-16'd14211;
      13429:data<=-16'd16869;
      13430:data<=-16'd16459;
      13431:data<=-16'd17202;
      13432:data<=-16'd16104;
      13433:data<=-16'd14942;
      13434:data<=-16'd15071;
      13435:data<=-16'd14334;
      13436:data<=-16'd13389;
      13437:data<=-16'd14123;
      13438:data<=-16'd15597;
      13439:data<=-16'd15409;
      13440:data<=-16'd14524;
      13441:data<=-16'd14701;
      13442:data<=-16'd14757;
      13443:data<=-16'd14358;
      13444:data<=-16'd13718;
      13445:data<=-16'd13602;
      13446:data<=-16'd14939;
      13447:data<=-16'd14980;
      13448:data<=-16'd13770;
      13449:data<=-16'd14043;
      13450:data<=-16'd13917;
      13451:data<=-16'd13353;
      13452:data<=-16'd13417;
      13453:data<=-16'd12457;
      13454:data<=-16'd12560;
      13455:data<=-16'd14366;
      13456:data<=-16'd14581;
      13457:data<=-16'd13552;
      13458:data<=-16'd12948;
      13459:data<=-16'd12903;
      13460:data<=-16'd12185;
      13461:data<=-16'd10919;
      13462:data<=-16'd11659;
      13463:data<=-16'd11755;
      13464:data<=-16'd8960;
      13465:data<=-16'd7450;
      13466:data<=-16'd7715;
      13467:data<=-16'd7985;
      13468:data<=-16'd7086;
      13469:data<=-16'd5365;
      13470:data<=-16'd6972;
      13471:data<=-16'd5586;
      13472:data<=16'd3912;
      13473:data<=16'd8293;
      13474:data<=16'd6064;
      13475:data<=16'd6492;
      13476:data<=16'd5771;
      13477:data<=16'd4958;
      13478:data<=16'd6680;
      13479:data<=16'd4948;
      13480:data<=16'd2687;
      13481:data<=16'd2714;
      13482:data<=16'd1949;
      13483:data<=16'd2359;
      13484:data<=16'd2813;
      13485:data<=16'd1938;
      13486:data<=16'd2094;
      13487:data<=16'd1398;
      13488:data<=-16'd30;
      13489:data<=-16'd308;
      13490:data<=-16'd453;
      13491:data<=-16'd338;
      13492:data<=-16'd626;
      13493:data<=-16'd1030;
      13494:data<=-16'd534;
      13495:data<=-16'd911;
      13496:data<=-16'd1680;
      13497:data<=-16'd2203;
      13498:data<=-16'd2842;
      13499:data<=-16'd2315;
      13500:data<=-16'd2003;
      13501:data<=-16'd2194;
      13502:data<=-16'd1683;
      13503:data<=-16'd2093;
      13504:data<=-16'd3065;
      13505:data<=-16'd4165;
      13506:data<=-16'd5154;
      13507:data<=-16'd4494;
      13508:data<=-16'd3908;
      13509:data<=-16'd3559;
      13510:data<=-16'd3495;
      13511:data<=-16'd4558;
      13512:data<=-16'd3800;
      13513:data<=-16'd4554;
      13514:data<=-16'd6548;
      13515:data<=-16'd3786;
      13516:data<=-16'd8291;
      13517:data<=-16'd22110;
      13518:data<=-16'd25784;
      13519:data<=-16'd22206;
      13520:data<=-16'd22183;
      13521:data<=-16'd21713;
      13522:data<=-16'd21679;
      13523:data<=-16'd21996;
      13524:data<=-16'd20371;
      13525:data<=-16'd19854;
      13526:data<=-16'd19097;
      13527:data<=-16'd17849;
      13528:data<=-16'd17329;
      13529:data<=-16'd16284;
      13530:data<=-16'd16897;
      13531:data<=-16'd17112;
      13532:data<=-16'd14916;
      13533:data<=-16'd14361;
      13534:data<=-16'd14242;
      13535:data<=-16'd13609;
      13536:data<=-16'd13564;
      13537:data<=-16'd12413;
      13538:data<=-16'd12405;
      13539:data<=-16'd13065;
      13540:data<=-16'd11658;
      13541:data<=-16'd11059;
      13542:data<=-16'd11059;
      13543:data<=-16'd10463;
      13544:data<=-16'd10161;
      13545:data<=-16'd9132;
      13546:data<=-16'd9056;
      13547:data<=-16'd9815;
      13548:data<=-16'd9074;
      13549:data<=-16'd8570;
      13550:data<=-16'd8026;
      13551:data<=-16'd6667;
      13552:data<=-16'd6055;
      13553:data<=-16'd5823;
      13554:data<=-16'd5615;
      13555:data<=-16'd5042;
      13556:data<=-16'd4353;
      13557:data<=-16'd3583;
      13558:data<=-16'd2267;
      13559:data<=-16'd2955;
      13560:data<=-16'd802;
      13561:data<=16'd8728;
      13562:data<=16'd14408;
      13563:data<=16'd14035;
      13564:data<=16'd15628;
      13565:data<=16'd15746;
      13566:data<=16'd14512;
      13567:data<=16'd14921;
      13568:data<=16'd13612;
      13569:data<=16'd13693;
      13570:data<=16'd16431;
      13571:data<=16'd17747;
      13572:data<=16'd18747;
      13573:data<=16'd19267;
      13574:data<=16'd18748;
      13575:data<=16'd18378;
      13576:data<=16'd17443;
      13577:data<=16'd16838;
      13578:data<=16'd16518;
      13579:data<=16'd16751;
      13580:data<=16'd18310;
      13581:data<=16'd17663;
      13582:data<=16'd16019;
      13583:data<=16'd16439;
      13584:data<=16'd16281;
      13585:data<=16'd15766;
      13586:data<=16'd15062;
      13587:data<=16'd13855;
      13588:data<=16'd14765;
      13589:data<=16'd15311;
      13590:data<=16'd14374;
      13591:data<=16'd14445;
      13592:data<=16'd13900;
      13593:data<=16'd13330;
      13594:data<=16'd13097;
      13595:data<=16'd11700;
      13596:data<=16'd11746;
      13597:data<=16'd13047;
      13598:data<=16'd13687;
      13599:data<=16'd13147;
      13600:data<=16'd11306;
      13601:data<=16'd11623;
      13602:data<=16'd11612;
      13603:data<=16'd9447;
      13604:data<=16'd11229;
      13605:data<=16'd8939;
      13606:data<=-16'd1833;
      13607:data<=-16'd5259;
      13608:data<=-16'd2443;
      13609:data<=-16'd3504;
      13610:data<=-16'd3215;
      13611:data<=-16'd2411;
      13612:data<=-16'd3864;
      13613:data<=-16'd2822;
      13614:data<=-16'd1193;
      13615:data<=-16'd694;
      13616:data<=-16'd70;
      13617:data<=-16'd604;
      13618:data<=-16'd578;
      13619:data<=-16'd335;
      13620:data<=-16'd1284;
      13621:data<=16'd58;
      13622:data<=16'd2015;
      13623:data<=16'd141;
      13624:data<=-16'd2663;
      13625:data<=-16'd2904;
      13626:data<=-16'd1798;
      13627:data<=-16'd1359;
      13628:data<=-16'd1838;
      13629:data<=-16'd1973;
      13630:data<=-16'd802;
      13631:data<=16'd488;
      13632:data<=16'd305;
      13633:data<=-16'd8;
      13634:data<=16'd652;
      13635:data<=16'd902;
      13636:data<=16'd916;
      13637:data<=16'd1231;
      13638:data<=16'd1864;
      13639:data<=16'd3300;
      13640:data<=16'd4041;
      13641:data<=16'd3889;
      13642:data<=16'd3830;
      13643:data<=16'd3143;
      13644:data<=16'd3125;
      13645:data<=16'd3425;
      13646:data<=16'd3422;
      13647:data<=16'd5530;
      13648:data<=16'd5774;
      13649:data<=16'd4851;
      13650:data<=16'd11949;
      13651:data<=16'd20174;
      13652:data<=16'd19916;
      13653:data<=16'd17881;
      13654:data<=16'd17491;
      13655:data<=16'd17475;
      13656:data<=16'd18457;
      13657:data<=16'd17735;
      13658:data<=16'd16302;
      13659:data<=16'd16316;
      13660:data<=16'd15888;
      13661:data<=16'd15414;
      13662:data<=16'd14804;
      13663:data<=16'd14140;
      13664:data<=16'd14966;
      13665:data<=16'd15126;
      13666:data<=16'd14084;
      13667:data<=16'd13453;
      13668:data<=16'd12748;
      13669:data<=16'd12243;
      13670:data<=16'd11535;
      13671:data<=16'd10886;
      13672:data<=16'd11580;
      13673:data<=16'd11832;
      13674:data<=16'd10933;
      13675:data<=16'd10149;
      13676:data<=16'd10922;
      13677:data<=16'd13370;
      13678:data<=16'd13107;
      13679:data<=16'd10980;
      13680:data<=16'd11917;
      13681:data<=16'd12414;
      13682:data<=16'd11007;
      13683:data<=16'd11132;
      13684:data<=16'd10771;
      13685:data<=16'd8942;
      13686:data<=16'd7868;
      13687:data<=16'd7846;
      13688:data<=16'd7318;
      13689:data<=16'd5633;
      13690:data<=16'd5526;
      13691:data<=16'd5538;
      13692:data<=16'd3933;
      13693:data<=16'd4723;
      13694:data<=16'd1583;
      13695:data<=-16'd9075;
      13696:data<=-16'd13899;
      13697:data<=-16'd12700;
      13698:data<=-16'd13976;
      13699:data<=-16'd14090;
      13700:data<=-16'd13515;
      13701:data<=-16'd14246;
      13702:data<=-16'd13283;
      13703:data<=-16'd12734;
      13704:data<=-16'd13097;
      13705:data<=-16'd13479;
      13706:data<=-16'd14842;
      13707:data<=-16'd14624;
      13708:data<=-16'd13579;
      13709:data<=-16'd13893;
      13710:data<=-16'd13982;
      13711:data<=-16'd13767;
      13712:data<=-16'd13241;
      13713:data<=-16'd13520;
      13714:data<=-16'd14959;
      13715:data<=-16'd14590;
      13716:data<=-16'd14058;
      13717:data<=-16'd14243;
      13718:data<=-16'd13279;
      13719:data<=-16'd13339;
      13720:data<=-16'd13403;
      13721:data<=-16'd12853;
      13722:data<=-16'd13799;
      13723:data<=-16'd13485;
      13724:data<=-16'd12907;
      13725:data<=-16'd13825;
      13726:data<=-16'd13483;
      13727:data<=-16'd13073;
      13728:data<=-16'd12054;
      13729:data<=-16'd11492;
      13730:data<=-16'd14938;
      13731:data<=-16'd16580;
      13732:data<=-16'd15641;
      13733:data<=-16'd16066;
      13734:data<=-16'd14956;
      13735:data<=-16'd14736;
      13736:data<=-16'd14663;
      13737:data<=-16'd12524;
      13738:data<=-16'd14337;
      13739:data<=-16'd11402;
      13740:data<=16'd105;
      13741:data<=16'd3002;
      13742:data<=16'd21;
      13743:data<=16'd1154;
      13744:data<=16'd417;
      13745:data<=-16'd56;
      13746:data<=16'd1550;
      13747:data<=16'd196;
      13748:data<=-16'd1251;
      13749:data<=-16'd1756;
      13750:data<=-16'd2094;
      13751:data<=-16'd1068;
      13752:data<=-16'd1280;
      13753:data<=-16'd1691;
      13754:data<=-16'd987;
      13755:data<=-16'd2162;
      13756:data<=-16'd3656;
      13757:data<=-16'd3539;
      13758:data<=-16'd3415;
      13759:data<=-16'd3445;
      13760:data<=-16'd3289;
      13761:data<=-16'd3280;
      13762:data<=-16'd3435;
      13763:data<=-16'd3571;
      13764:data<=-16'd4287;
      13765:data<=-16'd5356;
      13766:data<=-16'd5348;
      13767:data<=-16'd5178;
      13768:data<=-16'd5137;
      13769:data<=-16'd4610;
      13770:data<=-16'd4655;
      13771:data<=-16'd4287;
      13772:data<=-16'd4628;
      13773:data<=-16'd6869;
      13774:data<=-16'd7009;
      13775:data<=-16'd6431;
      13776:data<=-16'd6884;
      13777:data<=-16'd6088;
      13778:data<=-16'd6258;
      13779:data<=-16'd5538;
      13780:data<=-16'd4793;
      13781:data<=-16'd8417;
      13782:data<=-16'd7388;
      13783:data<=-16'd5136;
      13784:data<=-16'd13653;
      13785:data<=-16'd19394;
      13786:data<=-16'd16703;
      13787:data<=-16'd16416;
      13788:data<=-16'd16130;
      13789:data<=-16'd16010;
      13790:data<=-16'd17441;
      13791:data<=-16'd15791;
      13792:data<=-16'd15409;
      13793:data<=-16'd15964;
      13794:data<=-16'd14031;
      13795:data<=-16'd14038;
      13796:data<=-16'd13900;
      13797:data<=-16'd12727;
      13798:data<=-16'd13876;
      13799:data<=-16'd14061;
      13800:data<=-16'd13062;
      13801:data<=-16'd12628;
      13802:data<=-16'd12145;
      13803:data<=-16'd12041;
      13804:data<=-16'd10878;
      13805:data<=-16'd10615;
      13806:data<=-16'd12193;
      13807:data<=-16'd11294;
      13808:data<=-16'd9966;
      13809:data<=-16'd9893;
      13810:data<=-16'd8893;
      13811:data<=-16'd8282;
      13812:data<=-16'd7260;
      13813:data<=-16'd6493;
      13814:data<=-16'd7773;
      13815:data<=-16'd8084;
      13816:data<=-16'd7750;
      13817:data<=-16'd7492;
      13818:data<=-16'd6437;
      13819:data<=-16'd6228;
      13820:data<=-16'd5656;
      13821:data<=-16'd5142;
      13822:data<=-16'd5046;
      13823:data<=-16'd3392;
      13824:data<=-16'd3662;
      13825:data<=-16'd3621;
      13826:data<=-16'd1597;
      13827:data<=-16'd3568;
      13828:data<=16'd3;
      13829:data<=16'd11964;
      13830:data<=16'd15332;
      13831:data<=16'd13270;
      13832:data<=16'd14854;
      13833:data<=16'd14906;
      13834:data<=16'd15117;
      13835:data<=16'd14672;
      13836:data<=16'd10557;
      13837:data<=16'd9053;
      13838:data<=16'd9656;
      13839:data<=16'd10172;
      13840:data<=16'd12057;
      13841:data<=16'd11997;
      13842:data<=16'd11194;
      13843:data<=16'd11468;
      13844:data<=16'd10533;
      13845:data<=16'd10188;
      13846:data<=16'd10552;
      13847:data<=16'd11066;
      13848:data<=16'd12698;
      13849:data<=16'd12706;
      13850:data<=16'd11731;
      13851:data<=16'd11729;
      13852:data<=16'd11232;
      13853:data<=16'd10909;
      13854:data<=16'd10323;
      13855:data<=16'd9530;
      13856:data<=16'd10514;
      13857:data<=16'd11106;
      13858:data<=16'd10801;
      13859:data<=16'd10972;
      13860:data<=16'd10473;
      13861:data<=16'd10184;
      13862:data<=16'd9981;
      13863:data<=16'd8821;
      13864:data<=16'd8669;
      13865:data<=16'd9632;
      13866:data<=16'd10322;
      13867:data<=16'd10188;
      13868:data<=16'd9594;
      13869:data<=16'd9386;
      13870:data<=16'd8648;
      13871:data<=16'd8617;
      13872:data<=16'd8135;
      13873:data<=16'd1568;
      13874:data<=-16'd5271;
      13875:data<=-16'd4919;
      13876:data<=-16'd3559;
      13877:data<=-16'd3924;
      13878:data<=-16'd3654;
      13879:data<=-16'd4059;
      13880:data<=-16'd3535;
      13881:data<=-16'd1660;
      13882:data<=-16'd610;
      13883:data<=-16'd21;
      13884:data<=-16'd693;
      13885:data<=-16'd1425;
      13886:data<=-16'd177;
      13887:data<=-16'd32;
      13888:data<=-16'd375;
      13889:data<=16'd2904;
      13890:data<=16'd6678;
      13891:data<=16'd6607;
      13892:data<=16'd5368;
      13893:data<=16'd5714;
      13894:data<=16'd6134;
      13895:data<=16'd6205;
      13896:data<=16'd6067;
      13897:data<=16'd5582;
      13898:data<=16'd6784;
      13899:data<=16'd8188;
      13900:data<=16'd7614;
      13901:data<=16'd7720;
      13902:data<=16'd7539;
      13903:data<=16'd6360;
      13904:data<=16'd6957;
      13905:data<=16'd7095;
      13906:data<=16'd7242;
      13907:data<=16'd9273;
      13908:data<=16'd9318;
      13909:data<=16'd8590;
      13910:data<=16'd8769;
      13911:data<=16'd8176;
      13912:data<=16'd8431;
      13913:data<=16'd7994;
      13914:data<=16'd8204;
      13915:data<=16'd10566;
      13916:data<=16'd8959;
      13917:data<=16'd11189;
      13918:data<=16'd22324;
      13919:data<=16'd25519;
      13920:data<=16'd21303;
      13921:data<=16'd21346;
      13922:data<=16'd21218;
      13923:data<=16'd21290;
      13924:data<=16'd22635;
      13925:data<=16'd20676;
      13926:data<=16'd19452;
      13927:data<=16'd19261;
      13928:data<=16'd17861;
      13929:data<=16'd17914;
      13930:data<=16'd16810;
      13931:data<=16'd15717;
      13932:data<=16'd17614;
      13933:data<=16'd17479;
      13934:data<=16'd15753;
      13935:data<=16'd15447;
      13936:data<=16'd14916;
      13937:data<=16'd14587;
      13938:data<=16'd13826;
      13939:data<=16'd12824;
      13940:data<=16'd13587;
      13941:data<=16'd13209;
      13942:data<=16'd10326;
      13943:data<=16'd8019;
      13944:data<=16'd7447;
      13945:data<=16'd7204;
      13946:data<=16'd6152;
      13947:data<=16'd5946;
      13948:data<=16'd6796;
      13949:data<=16'd6595;
      13950:data<=16'd6256;
      13951:data<=16'd6061;
      13952:data<=16'd5470;
      13953:data<=16'd5392;
      13954:data<=16'd4955;
      13955:data<=16'd4328;
      13956:data<=16'd3771;
      13957:data<=16'd3008;
      13958:data<=16'd3206;
      13959:data<=16'd2085;
      13960:data<=16'd1253;
      13961:data<=16'd3051;
      13962:data<=-16'd2193;
      13963:data<=-16'd12841;
      13964:data<=-16'd15245;
      13965:data<=-16'd13796;
      13966:data<=-16'd14913;
      13967:data<=-16'd14733;
      13968:data<=-16'd14659;
      13969:data<=-16'd14860;
      13970:data<=-16'd13740;
      13971:data<=-16'd13274;
      13972:data<=-16'd12871;
      13973:data<=-16'd13421;
      13974:data<=-16'd14697;
      13975:data<=-16'd13709;
      13976:data<=-16'd13267;
      13977:data<=-16'd13896;
      13978:data<=-16'd12886;
      13979:data<=-16'd12296;
      13980:data<=-16'd12328;
      13981:data<=-16'd12483;
      13982:data<=-16'd13635;
      13983:data<=-16'd13600;
      13984:data<=-16'd12669;
      13985:data<=-16'd12493;
      13986:data<=-16'd11958;
      13987:data<=-16'd11367;
      13988:data<=-16'd10975;
      13989:data<=-16'd10702;
      13990:data<=-16'd11438;
      13991:data<=-16'd11819;
      13992:data<=-16'd10937;
      13993:data<=-16'd10598;
      13994:data<=-16'd10933;
      13995:data<=-16'd9436;
      13996:data<=-16'd6068;
      13997:data<=-16'd4417;
      13998:data<=-16'd5444;
      13999:data<=-16'd6925;
      14000:data<=-16'd7168;
      14001:data<=-16'd6197;
      14002:data<=-16'd6334;
      14003:data<=-16'd6517;
      14004:data<=-16'd5307;
      14005:data<=-16'd6308;
      14006:data<=-16'd4755;
      14007:data<=16'd3762;
      14008:data<=16'd8170;
      14009:data<=16'd6329;
      14010:data<=16'd6536;
      14011:data<=16'd6630;
      14012:data<=16'd5557;
      14013:data<=16'd5891;
      14014:data<=16'd5527;
      14015:data<=16'd4623;
      14016:data<=16'd3597;
      14017:data<=16'd2278;
      14018:data<=16'd2296;
      14019:data<=16'd2614;
      14020:data<=16'd2578;
      14021:data<=16'd2538;
      14022:data<=16'd2009;
      14023:data<=16'd1216;
      14024:data<=16'd24;
      14025:data<=16'd156;
      14026:data<=16'd1019;
      14027:data<=-16'd473;
      14028:data<=-16'd1037;
      14029:data<=-16'd47;
      14030:data<=-16'd773;
      14031:data<=-16'd1518;
      14032:data<=-16'd2558;
      14033:data<=-16'd3310;
      14034:data<=-16'd2646;
      14035:data<=-16'd3676;
      14036:data<=-16'd3683;
      14037:data<=-16'd2605;
      14038:data<=-16'd4106;
      14039:data<=-16'd3877;
      14040:data<=-16'd3826;
      14041:data<=-16'd6167;
      14042:data<=-16'd5659;
      14043:data<=-16'd5221;
      14044:data<=-16'd5233;
      14045:data<=-16'd4490;
      14046:data<=-16'd6243;
      14047:data<=-16'd5424;
      14048:data<=-16'd6091;
      14049:data<=-16'd11676;
      14050:data<=-16'd10446;
      14051:data<=-16'd12472;
      14052:data<=-16'd24641;
      14053:data<=-16'd26996;
      14054:data<=-16'd22889;
      14055:data<=-16'd23698;
      14056:data<=-16'd22803;
      14057:data<=-16'd22466;
      14058:data<=-16'd23143;
      14059:data<=-16'd21197;
      14060:data<=-16'd20961;
      14061:data<=-16'd20350;
      14062:data<=-16'd19121;
      14063:data<=-16'd19520;
      14064:data<=-16'd17617;
      14065:data<=-16'd17080;
      14066:data<=-16'd19027;
      14067:data<=-16'd17898;
      14068:data<=-16'd16719;
      14069:data<=-16'd16692;
      14070:data<=-16'd15681;
      14071:data<=-16'd15036;
      14072:data<=-16'd14111;
      14073:data<=-16'd14117;
      14074:data<=-16'd15417;
      14075:data<=-16'd14748;
      14076:data<=-16'd13468;
      14077:data<=-16'd13236;
      14078:data<=-16'd12786;
      14079:data<=-16'd11887;
      14080:data<=-16'd10793;
      14081:data<=-16'd10235;
      14082:data<=-16'd10220;
      14083:data<=-16'd10571;
      14084:data<=-16'd10793;
      14085:data<=-16'd9426;
      14086:data<=-16'd8167;
      14087:data<=-16'd8085;
      14088:data<=-16'd7732;
      14089:data<=-16'd7357;
      14090:data<=-16'd6416;
      14091:data<=-16'd5914;
      14092:data<=-16'd6062;
      14093:data<=-16'd4388;
      14094:data<=-16'd4241;
      14095:data<=-16'd2984;
      14096:data<=16'd5929;
      14097:data<=16'd12546;
      14098:data<=16'd12305;
      14099:data<=16'd13326;
      14100:data<=16'd13559;
      14101:data<=16'd13491;
      14102:data<=16'd16938;
      14103:data<=16'd17637;
      14104:data<=16'd15834;
      14105:data<=16'd15858;
      14106:data<=16'd15540;
      14107:data<=16'd15916;
      14108:data<=16'd17054;
      14109:data<=16'd16515;
      14110:data<=16'd15785;
      14111:data<=16'd15309;
      14112:data<=16'd15127;
      14113:data<=16'd15226;
      14114:data<=16'd14331;
      14115:data<=16'd14522;
      14116:data<=16'd15731;
      14117:data<=16'd15192;
      14118:data<=16'd14583;
      14119:data<=16'd14419;
      14120:data<=16'd13521;
      14121:data<=16'd13107;
      14122:data<=16'd12555;
      14123:data<=16'd11950;
      14124:data<=16'd13103;
      14125:data<=16'd13908;
      14126:data<=16'd12948;
      14127:data<=16'd12190;
      14128:data<=16'd11735;
      14129:data<=16'd11432;
      14130:data<=16'd11577;
      14131:data<=16'd10715;
      14132:data<=16'd10176;
      14133:data<=16'd11791;
      14134:data<=16'd11955;
      14135:data<=16'd10484;
      14136:data<=16'd10912;
      14137:data<=16'd10144;
      14138:data<=16'd8495;
      14139:data<=16'd9993;
      14140:data<=16'd6960;
      14141:data<=-16'd2437;
      14142:data<=-16'd5727;
      14143:data<=-16'd3615;
      14144:data<=-16'd4079;
      14145:data<=-16'd4168;
      14146:data<=-16'd3536;
      14147:data<=-16'd4331;
      14148:data<=-16'd3856;
      14149:data<=-16'd2570;
      14150:data<=-16'd1765;
      14151:data<=-16'd1384;
      14152:data<=-16'd1592;
      14153:data<=-16'd740;
      14154:data<=-16'd1410;
      14155:data<=-16'd5230;
      14156:data<=-16'd6226;
      14157:data<=-16'd4214;
      14158:data<=-16'd3366;
      14159:data<=-16'd2898;
      14160:data<=-16'd2895;
      14161:data<=-16'd3265;
      14162:data<=-16'd2657;
      14163:data<=-16'd2129;
      14164:data<=-16'd1588;
      14165:data<=-16'd676;
      14166:data<=-16'd89;
      14167:data<=16'd626;
      14168:data<=16'd1115;
      14169:data<=16'd763;
      14170:data<=16'd140;
      14171:data<=16'd405;
      14172:data<=16'd1401;
      14173:data<=16'd1407;
      14174:data<=16'd1792;
      14175:data<=16'd3195;
      14176:data<=16'd3102;
      14177:data<=16'd2729;
      14178:data<=16'd2899;
      14179:data<=16'd2711;
      14180:data<=16'd2854;
      14181:data<=16'd2390;
      14182:data<=16'd3216;
      14183:data<=16'd4948;
      14184:data<=16'd4517;
      14185:data<=16'd9547;
      14186:data<=16'd18592;
      14187:data<=16'd19311;
      14188:data<=16'd17450;
      14189:data<=16'd18281;
      14190:data<=16'd17079;
      14191:data<=16'd17453;
      14192:data<=16'd18225;
      14193:data<=16'd16170;
      14194:data<=16'd15449;
      14195:data<=16'd14892;
      14196:data<=16'd14413;
      14197:data<=16'd14592;
      14198:data<=16'd12801;
      14199:data<=16'd13063;
      14200:data<=16'd14783;
      14201:data<=16'd14023;
      14202:data<=16'd13782;
      14203:data<=16'd12853;
      14204:data<=16'd11442;
      14205:data<=16'd11885;
      14206:data<=16'd10689;
      14207:data<=16'd10994;
      14208:data<=16'd14678;
      14209:data<=16'd15289;
      14210:data<=16'd13822;
      14211:data<=16'd13180;
      14212:data<=16'd12428;
      14213:data<=16'd11862;
      14214:data<=16'd10637;
      14215:data<=16'd9950;
      14216:data<=16'd10836;
      14217:data<=16'd10860;
      14218:data<=16'd10082;
      14219:data<=16'd9247;
      14220:data<=16'd8507;
      14221:data<=16'd8596;
      14222:data<=16'd8552;
      14223:data<=16'd7482;
      14224:data<=16'd6285;
      14225:data<=16'd6545;
      14226:data<=16'd6237;
      14227:data<=16'd4306;
      14228:data<=16'd4934;
      14229:data<=16'd2420;
      14230:data<=-16'd7735;
      14231:data<=-16'd12555;
      14232:data<=-16'd10986;
      14233:data<=-16'd12525;
      14234:data<=-16'd13192;
      14235:data<=-16'd12331;
      14236:data<=-16'd12743;
      14237:data<=-16'd12020;
      14238:data<=-16'd12217;
      14239:data<=-16'd12507;
      14240:data<=-16'd11741;
      14241:data<=-16'd13050;
      14242:data<=-16'd13723;
      14243:data<=-16'd13567;
      14244:data<=-16'd14082;
      14245:data<=-16'd12880;
      14246:data<=-16'd12895;
      14247:data<=-16'd13703;
      14248:data<=-16'd12417;
      14249:data<=-16'd12998;
      14250:data<=-16'd14119;
      14251:data<=-16'd13156;
      14252:data<=-16'd12807;
      14253:data<=-16'd12430;
      14254:data<=-16'd11967;
      14255:data<=-16'd11899;
      14256:data<=-16'd10962;
      14257:data<=-16'd11130;
      14258:data<=-16'd12410;
      14259:data<=-16'd12354;
      14260:data<=-16'd11972;
      14261:data<=-16'd13300;
      14262:data<=-16'd15067;
      14263:data<=-16'd14451;
      14264:data<=-16'd13546;
      14265:data<=-16'd14148;
      14266:data<=-16'd14137;
      14267:data<=-16'd15233;
      14268:data<=-16'd16090;
      14269:data<=-16'd14233;
      14270:data<=-16'd14107;
      14271:data<=-16'd13474;
      14272:data<=-16'd11541;
      14273:data<=-16'd13156;
      14274:data<=-16'd9403;
      14275:data<=16'd593;
      14276:data<=16'd2807;
      14277:data<=16'd629;
      14278:data<=16'd1497;
      14279:data<=16'd1639;
      14280:data<=16'd1478;
      14281:data<=16'd1767;
      14282:data<=16'd1165;
      14283:data<=16'd514;
      14284:data<=-16'd651;
      14285:data<=-16'd1283;
      14286:data<=-16'd816;
      14287:data<=-16'd1033;
      14288:data<=-16'd1410;
      14289:data<=-16'd1066;
      14290:data<=-16'd361;
      14291:data<=-16'd945;
      14292:data<=-16'd3019;
      14293:data<=-16'd3322;
      14294:data<=-16'd2452;
      14295:data<=-16'd2641;
      14296:data<=-16'd2731;
      14297:data<=-16'd2963;
      14298:data<=-16'd3218;
      14299:data<=-16'd3412;
      14300:data<=-16'd4798;
      14301:data<=-16'd5518;
      14302:data<=-16'd5043;
      14303:data<=-16'd4726;
      14304:data<=-16'd4510;
      14305:data<=-16'd5165;
      14306:data<=-16'd5332;
      14307:data<=-16'd4613;
      14308:data<=-16'd5480;
      14309:data<=-16'd6534;
      14310:data<=-16'd6484;
      14311:data<=-16'd5523;
      14312:data<=-16'd4543;
      14313:data<=-16'd5598;
      14314:data<=-16'd4159;
      14315:data<=-16'd249;
      14316:data<=-16'd999;
      14317:data<=-16'd2187;
      14318:data<=-16'd3990;
      14319:data<=-16'd12690;
      14320:data<=-16'd18128;
      14321:data<=-16'd16409;
      14322:data<=-16'd16120;
      14323:data<=-16'd15716;
      14324:data<=-16'd15233;
      14325:data<=-16'd16712;
      14326:data<=-16'd15905;
      14327:data<=-16'd14522;
      14328:data<=-16'd14201;
      14329:data<=-16'd13060;
      14330:data<=-16'd12795;
      14331:data<=-16'd12358;
      14332:data<=-16'd11536;
      14333:data<=-16'd12474;
      14334:data<=-16'd12974;
      14335:data<=-16'd12552;
      14336:data<=-16'd12031;
      14337:data<=-16'd10937;
      14338:data<=-16'd10715;
      14339:data<=-16'd10366;
      14340:data<=-16'd8945;
      14341:data<=-16'd8671;
      14342:data<=-16'd9227;
      14343:data<=-16'd9324;
      14344:data<=-16'd8758;
      14345:data<=-16'd7671;
      14346:data<=-16'd7138;
      14347:data<=-16'd7015;
      14348:data<=-16'd6628;
      14349:data<=-16'd6114;
      14350:data<=-16'd6193;
      14351:data<=-16'd6931;
      14352:data<=-16'd6394;
      14353:data<=-16'd5426;
      14354:data<=-16'd5398;
      14355:data<=-16'd4730;
      14356:data<=-16'd4804;
      14357:data<=-16'd4648;
      14358:data<=-16'd2645;
      14359:data<=-16'd3031;
      14360:data<=-16'd2940;
      14361:data<=-16'd1369;
      14362:data<=-16'd3442;
      14363:data<=16'd928;
      14364:data<=16'd12618;
      14365:data<=16'd15239;
      14366:data<=16'd13411;
      14367:data<=16'd14196;
      14368:data<=16'd11361;
      14369:data<=16'd10088;
      14370:data<=16'd11714;
      14371:data<=16'd10460;
      14372:data<=16'd10487;
      14373:data<=16'd10942;
      14374:data<=16'd10088;
      14375:data<=16'd11881;
      14376:data<=16'd12531;
      14377:data<=16'd11489;
      14378:data<=16'd12378;
      14379:data<=16'd12269;
      14380:data<=16'd11655;
      14381:data<=16'd11664;
      14382:data<=16'd10677;
      14383:data<=16'd11280;
      14384:data<=16'd12687;
      14385:data<=16'd12160;
      14386:data<=16'd11656;
      14387:data<=16'd11414;
      14388:data<=16'd11036;
      14389:data<=16'd11251;
      14390:data<=16'd10950;
      14391:data<=16'd10533;
      14392:data<=16'd11156;
      14393:data<=16'd11573;
      14394:data<=16'd10994;
      14395:data<=16'd10598;
      14396:data<=16'd10737;
      14397:data<=16'd10217;
      14398:data<=16'd9447;
      14399:data<=16'd9652;
      14400:data<=16'd10440;
      14401:data<=16'd10953;
      14402:data<=16'd10613;
      14403:data<=16'd10419;
      14404:data<=16'd10434;
      14405:data<=16'd9353;
      14406:data<=16'd9520;
      14407:data<=16'd8737;
      14408:data<=16'd1789;
      14409:data<=-16'd4149;
      14410:data<=-16'd4015;
      14411:data<=-16'd4015;
      14412:data<=-16'd4168;
      14413:data<=-16'd2939;
      14414:data<=-16'd3068;
      14415:data<=-16'd3306;
      14416:data<=-16'd2561;
      14417:data<=-16'd1187;
      14418:data<=-16'd88;
      14419:data<=-16'd698;
      14420:data<=16'd262;
      14421:data<=16'd3257;
      14422:data<=16'd4253;
      14423:data<=16'd3865;
      14424:data<=16'd3328;
      14425:data<=16'd3797;
      14426:data<=16'd6020;
      14427:data<=16'd6514;
      14428:data<=16'd5520;
      14429:data<=16'd5510;
      14430:data<=16'd5600;
      14431:data<=16'd5835;
      14432:data<=16'd5815;
      14433:data<=16'd5985;
      14434:data<=16'd7338;
      14435:data<=16'd7677;
      14436:data<=16'd7506;
      14437:data<=16'd7567;
      14438:data<=16'd6711;
      14439:data<=16'd6584;
      14440:data<=16'd6419;
      14441:data<=16'd6170;
      14442:data<=16'd7661;
      14443:data<=16'd8059;
      14444:data<=16'd7700;
      14445:data<=16'd7900;
      14446:data<=16'd7253;
      14447:data<=16'd7806;
      14448:data<=16'd7638;
      14449:data<=16'd6322;
      14450:data<=16'd7470;
      14451:data<=16'd7207;
      14452:data<=16'd9865;
      14453:data<=16'd19776;
      14454:data<=16'd23093;
      14455:data<=16'd19772;
      14456:data<=16'd20175;
      14457:data<=16'd19666;
      14458:data<=16'd18769;
      14459:data<=16'd20451;
      14460:data<=16'd19878;
      14461:data<=16'd18703;
      14462:data<=16'd17770;
      14463:data<=16'd16089;
      14464:data<=16'd16362;
      14465:data<=16'd16143;
      14466:data<=16'd15138;
      14467:data<=16'd15755;
      14468:data<=16'd15790;
      14469:data<=16'd15532;
      14470:data<=16'd14725;
      14471:data<=16'd13065;
      14472:data<=16'd13355;
      14473:data<=16'd12129;
      14474:data<=16'd8035;
      14475:data<=16'd6898;
      14476:data<=16'd7877;
      14477:data<=16'd7389;
      14478:data<=16'd6766;
      14479:data<=16'd6886;
      14480:data<=16'd6551;
      14481:data<=16'd5627;
      14482:data<=16'd5486;
      14483:data<=16'd5659;
      14484:data<=16'd5850;
      14485:data<=16'd6689;
      14486:data<=16'd5780;
      14487:data<=16'd4085;
      14488:data<=16'd4138;
      14489:data<=16'd3680;
      14490:data<=16'd3651;
      14491:data<=16'd4038;
      14492:data<=16'd2737;
      14493:data<=16'd2772;
      14494:data<=16'd2123;
      14495:data<=16'd816;
      14496:data<=16'd2736;
      14497:data<=-16'd2306;
      14498:data<=-16'd13462;
      14499:data<=-16'd15130;
      14500:data<=-16'd13647;
      14501:data<=-16'd16198;
      14502:data<=-16'd15615;
      14503:data<=-16'd15012;
      14504:data<=-16'd16037;
      14505:data<=-16'd14791;
      14506:data<=-16'd14490;
      14507:data<=-16'd14327;
      14508:data<=-16'd13486;
      14509:data<=-16'd14930;
      14510:data<=-16'd15383;
      14511:data<=-16'd14484;
      14512:data<=-16'd14980;
      14513:data<=-16'd14847;
      14514:data<=-16'd14155;
      14515:data<=-16'd13691;
      14516:data<=-16'd13086;
      14517:data<=-16'd13782;
      14518:data<=-16'd14369;
      14519:data<=-16'd13511;
      14520:data<=-16'd13176;
      14521:data<=-16'd13206;
      14522:data<=-16'd12844;
      14523:data<=-16'd12504;
      14524:data<=-16'd12116;
      14525:data<=-16'd12580;
      14526:data<=-16'd12737;
      14527:data<=-16'd10073;
      14528:data<=-16'd7730;
      14529:data<=-16'd8073;
      14530:data<=-16'd7685;
      14531:data<=-16'd6909;
      14532:data<=-16'd7247;
      14533:data<=-16'd7018;
      14534:data<=-16'd8025;
      14535:data<=-16'd9364;
      14536:data<=-16'd8202;
      14537:data<=-16'd8179;
      14538:data<=-16'd8132;
      14539:data<=-16'd6736;
      14540:data<=-16'd8331;
      14541:data<=-16'd5506;
      14542:data<=16'd4299;
      14543:data<=16'd7729;
      14544:data<=16'd5733;
      14545:data<=16'd6041;
      14546:data<=16'd5770;
      14547:data<=16'd5353;
      14548:data<=16'd5533;
      14549:data<=16'd4760;
      14550:data<=16'd4353;
      14551:data<=16'd3087;
      14552:data<=16'd1888;
      14553:data<=16'd2209;
      14554:data<=16'd1697;
      14555:data<=16'd1642;
      14556:data<=16'd1877;
      14557:data<=16'd1283;
      14558:data<=16'd1688;
      14559:data<=16'd370;
      14560:data<=-16'd2118;
      14561:data<=-16'd2112;
      14562:data<=-16'd2099;
      14563:data<=-16'd2027;
      14564:data<=-16'd1586;
      14565:data<=-16'd2147;
      14566:data<=-16'd1442;
      14567:data<=-16'd1648;
      14568:data<=-16'd3527;
      14569:data<=-16'd3509;
      14570:data<=-16'd3559;
      14571:data<=-16'd3539;
      14572:data<=-16'd3181;
      14573:data<=-16'd4564;
      14574:data<=-16'd3853;
      14575:data<=-16'd2676;
      14576:data<=-16'd4740;
      14577:data<=-16'd5694;
      14578:data<=-16'd5385;
      14579:data<=-16'd5278;
      14580:data<=-16'd6119;
      14581:data<=-16'd9132;
      14582:data<=-16'd9204;
      14583:data<=-16'd8287;
      14584:data<=-16'd9891;
      14585:data<=-16'd8758;
      14586:data<=-16'd12193;
      14587:data<=-16'd22651;
      14588:data<=-16'd25402;
      14589:data<=-16'd22876;
      14590:data<=-16'd22776;
      14591:data<=-16'd21343;
      14592:data<=-16'd21205;
      14593:data<=-16'd22254;
      14594:data<=-16'd21062;
      14595:data<=-16'd20824;
      14596:data<=-16'd20118;
      14597:data<=-16'd18556;
      14598:data<=-16'd18930;
      14599:data<=-16'd18096;
      14600:data<=-16'd16671;
      14601:data<=-16'd17218;
      14602:data<=-16'd17394;
      14603:data<=-16'd16924;
      14604:data<=-16'd15881;
      14605:data<=-16'd14486;
      14606:data<=-16'd14651;
      14607:data<=-16'd14495;
      14608:data<=-16'd13129;
      14609:data<=-16'd13377;
      14610:data<=-16'd14378;
      14611:data<=-16'd13752;
      14612:data<=-16'd12707;
      14613:data<=-16'd12126;
      14614:data<=-16'd11074;
      14615:data<=-16'd10287;
      14616:data<=-16'd10199;
      14617:data<=-16'd10149;
      14618:data<=-16'd10939;
      14619:data<=-16'd11192;
      14620:data<=-16'd9721;
      14621:data<=-16'd9127;
      14622:data<=-16'd8853;
      14623:data<=-16'd7920;
      14624:data<=-16'd7583;
      14625:data<=-16'd6435;
      14626:data<=-16'd5894;
      14627:data<=-16'd6517;
      14628:data<=-16'd5172;
      14629:data<=-16'd4796;
      14630:data<=-16'd3196;
      14631:data<=16'd5362;
      14632:data<=16'd11949;
      14633:data<=16'd12745;
      14634:data<=16'd15637;
      14635:data<=16'd17970;
      14636:data<=16'd16816;
      14637:data<=16'd16725;
      14638:data<=16'd17098;
      14639:data<=16'd16536;
      14640:data<=16'd15687;
      14641:data<=16'd14519;
      14642:data<=16'd14786;
      14643:data<=16'd15852;
      14644:data<=16'd15632;
      14645:data<=16'd15335;
      14646:data<=16'd15488;
      14647:data<=16'd15374;
      14648:data<=16'd15012;
      14649:data<=16'd14075;
      14650:data<=16'd13259;
      14651:data<=16'd13908;
      14652:data<=16'd15097;
      14653:data<=16'd15252;
      14654:data<=16'd14892;
      14655:data<=16'd14387;
      14656:data<=16'd13441;
      14657:data<=16'd13012;
      14658:data<=16'd12828;
      14659:data<=16'd12578;
      14660:data<=16'd13418;
      14661:data<=16'd13687;
      14662:data<=16'd12901;
      14663:data<=16'd13004;
      14664:data<=16'd12405;
      14665:data<=16'd11267;
      14666:data<=16'd11133;
      14667:data<=16'd10704;
      14668:data<=16'd11213;
      14669:data<=16'd11724;
      14670:data<=16'd10589;
      14671:data<=16'd11100;
      14672:data<=16'd10863;
      14673:data<=16'd9667;
      14674:data<=16'd11450;
      14675:data<=16'd7095;
      14676:data<=-16'd3359;
      14677:data<=-16'd5444;
      14678:data<=-16'd3011;
      14679:data<=-16'd3582;
      14680:data<=-16'd3145;
      14681:data<=-16'd2732;
      14682:data<=-16'd2917;
      14683:data<=-16'd2775;
      14684:data<=-16'd2814;
      14685:data<=-16'd349;
      14686:data<=-16'd50;
      14687:data<=-16'd4152;
      14688:data<=-16'd4858;
      14689:data<=-16'd4097;
      14690:data<=-16'd4869;
      14691:data<=-16'd4055;
      14692:data<=-16'd3798;
      14693:data<=-16'd2955;
      14694:data<=-16'd796;
      14695:data<=-16'd1139;
      14696:data<=-16'd1171;
      14697:data<=-16'd361;
      14698:data<=-16'd717;
      14699:data<=-16'd164;
      14700:data<=-16'd346;
      14701:data<=-16'd552;
      14702:data<=16'd1110;
      14703:data<=16'd1410;
      14704:data<=16'd1425;
      14705:data<=16'd1759;
      14706:data<=16'd1074;
      14707:data<=16'd1471;
      14708:data<=16'd1303;
      14709:data<=16'd946;
      14710:data<=16'd2669;
      14711:data<=16'd3184;
      14712:data<=16'd3230;
      14713:data<=16'd3739;
      14714:data<=16'd2972;
      14715:data<=16'd2995;
      14716:data<=16'd2628;
      14717:data<=16'd2241;
      14718:data<=16'd3530;
      14719:data<=16'd4109;
      14720:data<=16'd9777;
      14721:data<=16'd19385;
      14722:data<=16'd20515;
      14723:data<=16'd18023;
      14724:data<=16'd18307;
      14725:data<=16'd16894;
      14726:data<=16'd16724;
      14727:data<=16'd17579;
      14728:data<=16'd16093;
      14729:data<=16'd15662;
      14730:data<=16'd15311;
      14731:data<=16'd14387;
      14732:data<=16'd14622;
      14733:data<=16'd13840;
      14734:data<=16'd13306;
      14735:data<=16'd13875;
      14736:data<=16'd13813;
      14737:data<=16'd13584;
      14738:data<=16'd12383;
      14739:data<=16'd12595;
      14740:data<=16'd15708;
      14741:data<=16'd16020;
      14742:data<=16'd14198;
      14743:data<=16'd15006;
      14744:data<=16'd16201;
      14745:data<=16'd15559;
      14746:data<=16'd14223;
      14747:data<=16'd13411;
      14748:data<=16'd12971;
      14749:data<=16'd12044;
      14750:data<=16'd11427;
      14751:data<=16'd11588;
      14752:data<=16'd12028;
      14753:data<=16'd12070;
      14754:data<=16'd11130;
      14755:data<=16'd10546;
      14756:data<=16'd10293;
      14757:data<=16'd9502;
      14758:data<=16'd8839;
      14759:data<=16'd7747;
      14760:data<=16'd7147;
      14761:data<=16'd6901;
      14762:data<=16'd5891;
      14763:data<=16'd6852;
      14764:data<=16'd3927;
      14765:data<=-16'd7221;
      14766:data<=-16'd12709;
      14767:data<=-16'd9940;
      14768:data<=-16'd10176;
      14769:data<=-16'd11527;
      14770:data<=-16'd11541;
      14771:data<=-16'd12129;
      14772:data<=-16'd11174;
      14773:data<=-16'd10827;
      14774:data<=-16'd11210;
      14775:data<=-16'd9467;
      14776:data<=-16'd8950;
      14777:data<=-16'd10147;
      14778:data<=-16'd10484;
      14779:data<=-16'd10749;
      14780:data<=-16'd10748;
      14781:data<=-16'd10252;
      14782:data<=-16'd9926;
      14783:data<=-16'd9586;
      14784:data<=-16'd9509;
      14785:data<=-16'd10120;
      14786:data<=-16'd11271;
      14787:data<=-16'd11488;
      14788:data<=-16'd10568;
      14789:data<=-16'd10461;
      14790:data<=-16'd10419;
      14791:data<=-16'd9445;
      14792:data<=-16'd9518;
      14793:data<=-16'd11979;
      14794:data<=-16'd15130;
      14795:data<=-16'd15706;
      14796:data<=-16'd14800;
      14797:data<=-16'd14768;
      14798:data<=-16'd13900;
      14799:data<=-16'd13265;
      14800:data<=-16'd13170;
      14801:data<=-16'd11972;
      14802:data<=-16'd13113;
      14803:data<=-16'd14466;
      14804:data<=-16'd12945;
      14805:data<=-16'd13092;
      14806:data<=-16'd12464;
      14807:data<=-16'd11262;
      14808:data<=-16'd13436;
      14809:data<=-16'd8916;
      14810:data<=16'd1048;
      14811:data<=16'd2215;
      14812:data<=-16'd523;
      14813:data<=-16'd293;
      14814:data<=-16'd587;
      14815:data<=-16'd466;
      14816:data<=16'd49;
      14817:data<=16'd41;
      14818:data<=-16'd21;
      14819:data<=-16'd1941;
      14820:data<=-16'd3055;
      14821:data<=-16'd1938;
      14822:data<=-16'd2149;
      14823:data<=-16'd2496;
      14824:data<=-16'd1785;
      14825:data<=-16'd1618;
      14826:data<=-16'd1897;
      14827:data<=-16'd3052;
      14828:data<=-16'd4003;
      14829:data<=-16'd3518;
      14830:data<=-16'd3442;
      14831:data<=-16'd3694;
      14832:data<=-16'd3456;
      14833:data<=-16'd3327;
      14834:data<=-16'd2877;
      14835:data<=-16'd2910;
      14836:data<=-16'd4138;
      14837:data<=-16'd4934;
      14838:data<=-16'd4746;
      14839:data<=-16'd3974;
      14840:data<=-16'd3289;
      14841:data<=-16'd3601;
      14842:data<=-16'd3707;
      14843:data<=-16'd3565;
      14844:data<=-16'd5033;
      14845:data<=-16'd5389;
      14846:data<=-16'd2403;
      14847:data<=-16'd494;
      14848:data<=-16'd785;
      14849:data<=16'd35;
      14850:data<=16'd509;
      14851:data<=-16'd185;
      14852:data<=-16'd117;
      14853:data<=-16'd2752;
      14854:data<=-16'd9884;
      14855:data<=-16'd14863;
      14856:data<=-16'd14593;
      14857:data<=-16'd13496;
      14858:data<=-16'd13062;
      14859:data<=-16'd11906;
      14860:data<=-16'd11932;
      14861:data<=-16'd13113;
      14862:data<=-16'd12366;
      14863:data<=-16'd11292;
      14864:data<=-16'd11453;
      14865:data<=-16'd10578;
      14866:data<=-16'd9829;
      14867:data<=-16'd10073;
      14868:data<=-16'd9647;
      14869:data<=-16'd10178;
      14870:data<=-16'd11066;
      14871:data<=-16'd10100;
      14872:data<=-16'd9505;
      14873:data<=-16'd9332;
      14874:data<=-16'd8511;
      14875:data<=-16'd8439;
      14876:data<=-16'd8126;
      14877:data<=-16'd7964;
      14878:data<=-16'd9050;
      14879:data<=-16'd8848;
      14880:data<=-16'd7853;
      14881:data<=-16'd7550;
      14882:data<=-16'd6969;
      14883:data<=-16'd6965;
      14884:data<=-16'd6858;
      14885:data<=-16'd6337;
      14886:data<=-16'd7174;
      14887:data<=-16'd7092;
      14888:data<=-16'd5973;
      14889:data<=-16'd6037;
      14890:data<=-16'd5371;
      14891:data<=-16'd4880;
      14892:data<=-16'd5192;
      14893:data<=-16'd4167;
      14894:data<=-16'd3836;
      14895:data<=-16'd3298;
      14896:data<=-16'd2384;
      14897:data<=-16'd4247;
      14898:data<=-16'd1077;
      14899:data<=16'd7902;
      14900:data<=16'd9065;
      14901:data<=16'd5802;
      14902:data<=16'd7576;
      14903:data<=16'd8866;
      14904:data<=16'd8075;
      14905:data<=16'd8385;
      14906:data<=16'd8351;
      14907:data<=16'd8360;
      14908:data<=16'd8175;
      14909:data<=16'd7288;
      14910:data<=16'd8099;
      14911:data<=16'd9592;
      14912:data<=16'd9668;
      14913:data<=16'd9441;
      14914:data<=16'd9359;
      14915:data<=16'd9068;
      14916:data<=16'd8895;
      14917:data<=16'd8743;
      14918:data<=16'd8660;
      14919:data<=16'd9426;
      14920:data<=16'd10417;
      14921:data<=16'd10387;
      14922:data<=16'd10040;
      14923:data<=16'd9527;
      14924:data<=16'd8848;
      14925:data<=16'd9001;
      14926:data<=16'd8880;
      14927:data<=16'd9003;
      14928:data<=16'd10342;
      14929:data<=16'd10088;
      14930:data<=16'd9488;
      14931:data<=16'd10187;
      14932:data<=16'd9538;
      14933:data<=16'd9165;
      14934:data<=16'd9266;
      14935:data<=16'd8513;
      14936:data<=16'd9975;
      14937:data<=16'd10892;
      14938:data<=16'd9588;
      14939:data<=16'd10035;
      14940:data<=16'd9720;
      14941:data<=16'd9179;
      14942:data<=16'd9156;
      14943:data<=16'd2846;
      14944:data<=-16'd3949;
      14945:data<=-16'd3266;
      14946:data<=-16'd2020;
      14947:data<=-16'd2558;
      14948:data<=-16'd2152;
      14949:data<=-16'd1821;
      14950:data<=-16'd1472;
      14951:data<=-16'd1697;
      14952:data<=-16'd370;
      14953:data<=16'd4005;
      14954:data<=16'd5862;
      14955:data<=16'd4825;
      14956:data<=16'd4611;
      14957:data<=16'd4488;
      14958:data<=16'd4220;
      14959:data<=16'd3707;
      14960:data<=16'd3926;
      14961:data<=16'd5958;
      14962:data<=16'd6300;
      14963:data<=16'd5204;
      14964:data<=16'd5538;
      14965:data<=16'd5313;
      14966:data<=16'd4535;
      14967:data<=16'd4498;
      14968:data<=16'd4258;
      14969:data<=16'd4889;
      14970:data<=16'd6414;
      14971:data<=16'd6693;
      14972:data<=16'd5940;
      14973:data<=16'd5607;
      14974:data<=16'd5664;
      14975:data<=16'd5333;
      14976:data<=16'd5065;
      14977:data<=16'd5486;
      14978:data<=16'd6472;
      14979:data<=16'd7259;
      14980:data<=16'd6375;
      14981:data<=16'd5579;
      14982:data<=16'd6125;
      14983:data<=16'd5069;
      14984:data<=16'd4523;
      14985:data<=16'd5419;
      14986:data<=16'd4043;
      14987:data<=16'd7089;
      14988:data<=16'd16480;
      14989:data<=16'd19843;
      14990:data<=16'd17517;
      14991:data<=16'd17209;
      14992:data<=16'd16487;
      14993:data<=16'd15115;
      14994:data<=16'd15303;
      14995:data<=16'd15323;
      14996:data<=16'd14762;
      14997:data<=16'd14110;
      14998:data<=16'd13591;
      14999:data<=16'd12962;
      15000:data<=16'd11967;
      15001:data<=16'd11721;
      15002:data<=16'd11771;
      15003:data<=16'd12308;
      15004:data<=16'd13426;
      15005:data<=16'd11386;
      15006:data<=16'd7324;
      15007:data<=16'd6065;
      15008:data<=16'd6297;
      15009:data<=16'd5762;
      15010:data<=16'd5096;
      15011:data<=16'd5119;
      15012:data<=16'd5814;
      15013:data<=16'd5868;
      15014:data<=16'd5470;
      15015:data<=16'd5110;
      15016:data<=16'd4463;
      15017:data<=16'd4479;
      15018:data<=16'd4149;
      15019:data<=16'd3407;
      15020:data<=16'd4255;
      15021:data<=16'd4555;
      15022:data<=16'd3885;
      15023:data<=16'd3527;
      15024:data<=16'd1859;
      15025:data<=16'd1321;
      15026:data<=16'd2413;
      15027:data<=16'd1804;
      15028:data<=16'd1633;
      15029:data<=16'd1318;
      15030:data<=16'd419;
      15031:data<=16'd2102;
      15032:data<=-16'd1497;
      15033:data<=-16'd11770;
      15034:data<=-16'd14750;
      15035:data<=-16'd12000;
      15036:data<=-16'd12900;
      15037:data<=-16'd14149;
      15038:data<=-16'd14208;
      15039:data<=-16'd14085;
      15040:data<=-16'd12692;
      15041:data<=-16'd12633;
      15042:data<=-16'd13106;
      15043:data<=-16'd11937;
      15044:data<=-16'd12504;
      15045:data<=-16'd14366;
      15046:data<=-16'd14135;
      15047:data<=-16'd13333;
      15048:data<=-16'd13491;
      15049:data<=-16'd13505;
      15050:data<=-16'd12894;
      15051:data<=-16'd12135;
      15052:data<=-16'd11903;
      15053:data<=-16'd12636;
      15054:data<=-16'd13597;
      15055:data<=-16'd13297;
      15056:data<=-16'd12475;
      15057:data<=-16'd12659;
      15058:data<=-16'd11618;
      15059:data<=-16'd8187;
      15060:data<=-16'd6294;
      15061:data<=-16'd7507;
      15062:data<=-16'd8784;
      15063:data<=-16'd8774;
      15064:data<=-16'd8282;
      15065:data<=-16'd7835;
      15066:data<=-16'd7958;
      15067:data<=-16'd8020;
      15068:data<=-16'd7388;
      15069:data<=-16'd7938;
      15070:data<=-16'd9289;
      15071:data<=-16'd9016;
      15072:data<=-16'd8772;
      15073:data<=-16'd9012;
      15074:data<=-16'd8513;
      15075:data<=-16'd8893;
      15076:data<=-16'd6200;
      15077:data<=16'd1682;
      15078:data<=16'd5160;
      15079:data<=16'd3030;
      15080:data<=16'd2878;
      15081:data<=16'd3156;
      15082:data<=16'd2228;
      15083:data<=16'd2112;
      15084:data<=16'd1756;
      15085:data<=16'd1498;
      15086:data<=16'd1027;
      15087:data<=-16'd406;
      15088:data<=-16'd699;
      15089:data<=-16'd529;
      15090:data<=-16'd819;
      15091:data<=-16'd839;
      15092:data<=-16'd1104;
      15093:data<=-16'd546;
      15094:data<=-16'd384;
      15095:data<=-16'd2508;
      15096:data<=-16'd3489;
      15097:data<=-16'd2952;
      15098:data<=-16'd3107;
      15099:data<=-16'd2858;
      15100:data<=-16'd2781;
      15101:data<=-16'd3149;
      15102:data<=-16'd2878;
      15103:data<=-16'd3143;
      15104:data<=-16'd4070;
      15105:data<=-16'd4710;
      15106:data<=-16'd4443;
      15107:data<=-16'd3497;
      15108:data<=-16'd3849;
      15109:data<=-16'd4444;
      15110:data<=-16'd3858;
      15111:data<=-16'd5187;
      15112:data<=-16'd8863;
      15113:data<=-16'd10843;
      15114:data<=-16'd9832;
      15115:data<=-16'd9195;
      15116:data<=-16'd9997;
      15117:data<=-16'd8975;
      15118:data<=-16'd7978;
      15119:data<=-16'd8863;
      15120:data<=-16'd8334;
      15121:data<=-16'd11788;
      15122:data<=-16'd21030;
      15123:data<=-16'd23560;
      15124:data<=-16'd20243;
      15125:data<=-16'd20474;
      15126:data<=-16'd20010;
      15127:data<=-16'd17794;
      15128:data<=-16'd18389;
      15129:data<=-16'd19009;
      15130:data<=-16'd18472;
      15131:data<=-16'd17816;
      15132:data<=-16'd16186;
      15133:data<=-16'd15656;
      15134:data<=-16'd16114;
      15135:data<=-16'd14986;
      15136:data<=-16'd14343;
      15137:data<=-16'd15211;
      15138:data<=-16'd14960;
      15139:data<=-16'd13951;
      15140:data<=-16'd13482;
      15141:data<=-16'd12680;
      15142:data<=-16'd11838;
      15143:data<=-16'd11342;
      15144:data<=-16'd10769;
      15145:data<=-16'd11001;
      15146:data<=-16'd11442;
      15147:data<=-16'd10906;
      15148:data<=-16'd10320;
      15149:data<=-16'd9582;
      15150:data<=-16'd8980;
      15151:data<=-16'd9031;
      15152:data<=-16'd7962;
      15153:data<=-16'd7219;
      15154:data<=-16'd8216;
      15155:data<=-16'd7900;
      15156:data<=-16'd6795;
      15157:data<=-16'd6537;
      15158:data<=-16'd5900;
      15159:data<=-16'd5633;
      15160:data<=-16'd5421;
      15161:data<=-16'd4320;
      15162:data<=-16'd3773;
      15163:data<=-16'd3679;
      15164:data<=-16'd3204;
      15165:data<=16'd405;
      15166:data<=16'd9085;
      15167:data<=16'd15731;
      15168:data<=16'd15659;
      15169:data<=16'd14633;
      15170:data<=16'd15778;
      15171:data<=16'd16662;
      15172:data<=16'd15969;
      15173:data<=16'd14763;
      15174:data<=16'd14543;
      15175:data<=16'd14759;
      15176:data<=16'd14521;
      15177:data<=16'd13905;
      15178:data<=16'd13882;
      15179:data<=16'd15462;
      15180:data<=16'd16113;
      15181:data<=16'd14885;
      15182:data<=16'd14700;
      15183:data<=16'd14795;
      15184:data<=16'd14179;
      15185:data<=16'd13861;
      15186:data<=16'd13468;
      15187:data<=16'd14258;
      15188:data<=16'd15305;
      15189:data<=16'd14480;
      15190:data<=16'd14016;
      15191:data<=16'd13773;
      15192:data<=16'd13127;
      15193:data<=16'd13292;
      15194:data<=16'd12706;
      15195:data<=16'd12877;
      15196:data<=16'd14346;
      15197:data<=16'd13535;
      15198:data<=16'd12384;
      15199:data<=16'd12164;
      15200:data<=16'd11593;
      15201:data<=16'd11580;
      15202:data<=16'd10718;
      15203:data<=16'd10909;
      15204:data<=16'd13057;
      15205:data<=16'd12387;
      15206:data<=16'd11558;
      15207:data<=16'd11708;
      15208:data<=16'd10548;
      15209:data<=16'd11662;
      15210:data<=16'd8639;
      15211:data<=-16'd967;
      15212:data<=-16'd3369;
      15213:data<=-16'd435;
      15214:data<=-16'd766;
      15215:data<=-16'd408;
      15216:data<=16'd143;
      15217:data<=-16'd575;
      15218:data<=-16'd1801;
      15219:data<=-16'd4411;
      15220:data<=-16'd3976;
      15221:data<=-16'd1735;
      15222:data<=-16'd2111;
      15223:data<=-16'd1632;
      15224:data<=-16'd1096;
      15225:data<=-16'd1598;
      15226:data<=-16'd1046;
      15227:data<=-16'd1665;
      15228:data<=-16'd1248;
      15229:data<=16'd1116;
      15230:data<=16'd1101;
      15231:data<=16'd996;
      15232:data<=16'd1618;
      15233:data<=16'd1154;
      15234:data<=16'd1324;
      15235:data<=16'd819;
      15236:data<=16'd367;
      15237:data<=16'd2052;
      15238:data<=16'd3301;
      15239:data<=16'd3676;
      15240:data<=16'd2978;
      15241:data<=16'd1855;
      15242:data<=16'd2961;
      15243:data<=16'd3388;
      15244:data<=16'd2546;
      15245:data<=16'd3557;
      15246:data<=16'd4620;
      15247:data<=16'd4968;
      15248:data<=16'd4864;
      15249:data<=16'd4388;
      15250:data<=16'd4951;
      15251:data<=16'd4766;
      15252:data<=16'd4446;
      15253:data<=16'd4910;
      15254:data<=16'd4525;
      15255:data<=16'd9374;
      15256:data<=16'd18671;
      15257:data<=16'd20591;
      15258:data<=16'd17509;
      15259:data<=16'd17064;
      15260:data<=16'd16745;
      15261:data<=16'd15749;
      15262:data<=16'd15794;
      15263:data<=16'd16316;
      15264:data<=16'd16349;
      15265:data<=16'd15244;
      15266:data<=16'd13940;
      15267:data<=16'd13480;
      15268:data<=16'd13788;
      15269:data<=16'd13388;
      15270:data<=16'd12417;
      15271:data<=16'd14653;
      15272:data<=16'd17596;
      15273:data<=16'd16475;
      15274:data<=16'd15277;
      15275:data<=16'd15481;
      15276:data<=16'd14713;
      15277:data<=16'd14269;
      15278:data<=16'd13708;
      15279:data<=16'd13491;
      15280:data<=16'd14531;
      15281:data<=16'd14230;
      15282:data<=16'd13204;
      15283:data<=16'd12495;
      15284:data<=16'd11515;
      15285:data<=16'd11408;
      15286:data<=16'd11024;
      15287:data<=16'd10301;
      15288:data<=16'd10619;
      15289:data<=16'd10331;
      15290:data<=16'd9629;
      15291:data<=16'd9172;
      15292:data<=16'd8531;
      15293:data<=16'd8241;
      15294:data<=16'd7538;
      15295:data<=16'd6884;
      15296:data<=16'd6096;
      15297:data<=16'd5012;
      15298:data<=16'd5971;
      15299:data<=16'd3233;
      15300:data<=-16'd5755;
      15301:data<=-16'd10131;
      15302:data<=-16'd9395;
      15303:data<=-16'd10166;
      15304:data<=-16'd10507;
      15305:data<=-16'd10590;
      15306:data<=-16'd10836;
      15307:data<=-16'd9882;
      15308:data<=-16'd10028;
      15309:data<=-16'd10454;
      15310:data<=-16'd9867;
      15311:data<=-16'd9435;
      15312:data<=-16'd9450;
      15313:data<=-16'd10953;
      15314:data<=-16'd11823;
      15315:data<=-16'd10934;
      15316:data<=-16'd11179;
      15317:data<=-16'd10988;
      15318:data<=-16'd10046;
      15319:data<=-16'd10100;
      15320:data<=-16'd10113;
      15321:data<=-16'd11603;
      15322:data<=-16'd12483;
      15323:data<=-16'd10801;
      15324:data<=-16'd12337;
      15325:data<=-16'd15488;
      15326:data<=-16'd15588;
      15327:data<=-16'd14815;
      15328:data<=-16'd13671;
      15329:data<=-16'd13966;
      15330:data<=-16'd15693;
      15331:data<=-16'd14860;
      15332:data<=-16'd14125;
      15333:data<=-16'd14302;
      15334:data<=-16'd13045;
      15335:data<=-16'd12581;
      15336:data<=-16'd12311;
      15337:data<=-16'd12381;
      15338:data<=-16'd13433;
      15339:data<=-16'd12818;
      15340:data<=-16'd13010;
      15341:data<=-16'd13160;
      15342:data<=-16'd11600;
      15343:data<=-16'd12710;
      15344:data<=-16'd9042;
      15345:data<=16'd1019;
      15346:data<=16'd2649;
      15347:data<=-16'd337;
      15348:data<=16'd981;
      15349:data<=16'd523;
      15350:data<=-16'd502;
      15351:data<=16'd52;
      15352:data<=-16'd264;
      15353:data<=16'd770;
      15354:data<=16'd86;
      15355:data<=-16'd2676;
      15356:data<=-16'd2231;
      15357:data<=-16'd1765;
      15358:data<=-16'd2224;
      15359:data<=-16'd1624;
      15360:data<=-16'd2150;
      15361:data<=-16'd1797;
      15362:data<=-16'd1574;
      15363:data<=-16'd4024;
      15364:data<=-16'd4300;
      15365:data<=-16'd3149;
      15366:data<=-16'd3465;
      15367:data<=-16'd2796;
      15368:data<=-16'd2698;
      15369:data<=-16'd3066;
      15370:data<=-16'd2030;
      15371:data<=-16'd2978;
      15372:data<=-16'd4992;
      15373:data<=-16'd4840;
      15374:data<=-16'd4124;
      15375:data<=-16'd3949;
      15376:data<=-16'd4202;
      15377:data<=-16'd2872;
      15378:data<=16'd626;
      15379:data<=16'd970;
      15380:data<=-16'd1541;
      15381:data<=-16'd1497;
      15382:data<=-16'd804;
      15383:data<=-16'd1336;
      15384:data<=-16'd1178;
      15385:data<=-16'd1594;
      15386:data<=-16'd1902;
      15387:data<=-16'd773;
      15388:data<=-16'd3703;
      15389:data<=-16'd11817;
      15390:data<=-16'd16750;
      15391:data<=-16'd16099;
      15392:data<=-16'd15053;
      15393:data<=-16'd14712;
      15394:data<=-16'd13605;
      15395:data<=-16'd12533;
      15396:data<=-16'd12427;
      15397:data<=-16'd13207;
      15398:data<=-16'd13872;
      15399:data<=-16'd13345;
      15400:data<=-16'd12066;
      15401:data<=-16'd11354;
      15402:data<=-16'd11301;
      15403:data<=-16'd10709;
      15404:data<=-16'd10340;
      15405:data<=-16'd11191;
      15406:data<=-16'd11100;
      15407:data<=-16'd10097;
      15408:data<=-16'd10105;
      15409:data<=-16'd9814;
      15410:data<=-16'd9059;
      15411:data<=-16'd8625;
      15412:data<=-16'd8144;
      15413:data<=-16'd9138;
      15414:data<=-16'd10408;
      15415:data<=-16'd9241;
      15416:data<=-16'd7962;
      15417:data<=-16'd8144;
      15418:data<=-16'd8225;
      15419:data<=-16'd7313;
      15420:data<=-16'd5941;
      15421:data<=-16'd6223;
      15422:data<=-16'd7345;
      15423:data<=-16'd6799;
      15424:data<=-16'd5981;
      15425:data<=-16'd5817;
      15426:data<=-16'd5679;
      15427:data<=-16'd5192;
      15428:data<=-16'd3927;
      15429:data<=-16'd3475;
      15430:data<=-16'd3953;
      15431:data<=-16'd5621;
      15432:data<=-16'd8502;
      15433:data<=-16'd4352;
      15434:data<=16'd6126;
      15435:data<=16'd9139;
      15436:data<=16'd6845;
      15437:data<=16'd8240;
      15438:data<=16'd9476;
      15439:data<=16'd9218;
      15440:data<=16'd9685;
      15441:data<=16'd9520;
      15442:data<=16'd9467;
      15443:data<=16'd9559;
      15444:data<=16'd8824;
      15445:data<=16'd8361;
      15446:data<=16'd8810;
      15447:data<=16'd9961;
      15448:data<=16'd10440;
      15449:data<=16'd10099;
      15450:data<=16'd10184;
      15451:data<=16'd9932;
      15452:data<=16'd9802;
      15453:data<=16'd10035;
      15454:data<=16'd9753;
      15455:data<=16'd10704;
      15456:data<=16'd11732;
      15457:data<=16'd11025;
      15458:data<=16'd10912;
      15459:data<=16'd10898;
      15460:data<=16'd10202;
      15461:data<=16'd10006;
      15462:data<=16'd9888;
      15463:data<=16'd10830;
      15464:data<=16'd12284;
      15465:data<=16'd12440;
      15466:data<=16'd12182;
      15467:data<=16'd11339;
      15468:data<=16'd10997;
      15469:data<=16'd11391;
      15470:data<=16'd10169;
      15471:data<=16'd10204;
      15472:data<=16'd11724;
      15473:data<=16'd11521;
      15474:data<=16'd11644;
      15475:data<=16'd11044;
      15476:data<=16'd10081;
      15477:data<=16'd10448;
      15478:data<=16'd4739;
      15479:data<=-16'd3292;
      15480:data<=-16'd2908;
      15481:data<=-16'd1028;
      15482:data<=-16'd1949;
      15483:data<=-16'd922;
      15484:data<=16'd6;
      15485:data<=16'd576;
      15486:data<=16'd1263;
      15487:data<=16'd434;
      15488:data<=16'd1280;
      15489:data<=16'd3139;
      15490:data<=16'd3037;
      15491:data<=16'd3052;
      15492:data<=16'd3230;
      15493:data<=16'd2866;
      15494:data<=16'd2576;
      15495:data<=16'd2003;
      15496:data<=16'd2689;
      15497:data<=16'd4331;
      15498:data<=16'd4360;
      15499:data<=16'd3855;
      15500:data<=16'd4065;
      15501:data<=16'd4076;
      15502:data<=16'd3588;
      15503:data<=16'd2732;
      15504:data<=16'd2500;
      15505:data<=16'd3718;
      15506:data<=16'd4792;
      15507:data<=16'd4576;
      15508:data<=16'd4170;
      15509:data<=16'd3859;
      15510:data<=16'd3570;
      15511:data<=16'd3695;
      15512:data<=16'd3236;
      15513:data<=16'd3266;
      15514:data<=16'd5213;
      15515:data<=16'd5911;
      15516:data<=16'd5336;
      15517:data<=16'd5491;
      15518:data<=16'd4461;
      15519:data<=16'd4114;
      15520:data<=16'd4505;
      15521:data<=16'd3045;
      15522:data<=16'd7071;
      15523:data<=16'd16264;
      15524:data<=16'd18774;
      15525:data<=16'd16889;
      15526:data<=16'd16810;
      15527:data<=16'd15931;
      15528:data<=16'd14894;
      15529:data<=16'd14525;
      15530:data<=16'd14230;
      15531:data<=16'd14971;
      15532:data<=16'd14833;
      15533:data<=16'd13737;
      15534:data<=16'd13182;
      15535:data<=16'd12375;
      15536:data<=16'd11476;
      15537:data<=16'd9708;
      15538:data<=16'd8302;
      15539:data<=16'd9674;
      15540:data<=16'd10138;
      15541:data<=16'd8537;
      15542:data<=16'd7633;
      15543:data<=16'd6921;
      15544:data<=16'd6862;
      15545:data<=16'd6898;
      15546:data<=16'd6220;
      15547:data<=16'd7148;
      15548:data<=16'd7577;
      15549:data<=16'd6208;
      15550:data<=16'd6155;
      15551:data<=16'd6267;
      15552:data<=16'd5620;
      15553:data<=16'd5080;
      15554:data<=16'd4303;
      15555:data<=16'd4499;
      15556:data<=16'd4657;
      15557:data<=16'd4179;
      15558:data<=16'd4758;
      15559:data<=16'd4626;
      15560:data<=16'd3867;
      15561:data<=16'd3250;
      15562:data<=16'd1838;
      15563:data<=16'd2017;
      15564:data<=16'd2015;
      15565:data<=16'd978;
      15566:data<=16'd2320;
      15567:data<=-16'd1548;
      15568:data<=-16'd11414;
      15569:data<=-16'd13693;
      15570:data<=-16'd11056;
      15571:data<=-16'd12436;
      15572:data<=-16'd14011;
      15573:data<=-16'd14169;
      15574:data<=-16'd14113;
      15575:data<=-16'd13640;
      15576:data<=-16'd13879;
      15577:data<=-16'd13438;
      15578:data<=-16'd12160;
      15579:data<=-16'd11987;
      15580:data<=-16'd12731;
      15581:data<=-16'd13946;
      15582:data<=-16'd14304;
      15583:data<=-16'd13532;
      15584:data<=-16'd13080;
      15585:data<=-16'd12684;
      15586:data<=-16'd12367;
      15587:data<=-16'd11917;
      15588:data<=-16'd11785;
      15589:data<=-16'd13088;
      15590:data<=-16'd12695;
      15591:data<=-16'd10520;
      15592:data<=-16'd10267;
      15593:data<=-16'd10511;
      15594:data<=-16'd10307;
      15595:data<=-16'd10067;
      15596:data<=-16'd9332;
      15597:data<=-16'd10196;
      15598:data<=-16'd11462;
      15599:data<=-16'd11000;
      15600:data<=-16'd10436;
      15601:data<=-16'd9677;
      15602:data<=-16'd9420;
      15603:data<=-16'd9633;
      15604:data<=-16'd8596;
      15605:data<=-16'd8824;
      15606:data<=-16'd10050;
      15607:data<=-16'd9878;
      15608:data<=-16'd9441;
      15609:data<=-16'd8950;
      15610:data<=-16'd9629;
      15611:data<=-16'd7830;
      15612:data<=16'd798;
      15613:data<=16'd5504;
      15614:data<=16'd2523;
      15615:data<=16'd2033;
      15616:data<=16'd2864;
      15617:data<=16'd2312;
      15618:data<=16'd2776;
      15619:data<=16'd2059;
      15620:data<=16'd2015;
      15621:data<=16'd3181;
      15622:data<=16'd1594;
      15623:data<=-16'd121;
      15624:data<=-16'd253;
      15625:data<=-16'd115;
      15626:data<=16'd314;
      15627:data<=-16'd393;
      15628:data<=-16'd509;
      15629:data<=16'd652;
      15630:data<=-16'd425;
      15631:data<=-16'd2323;
      15632:data<=-16'd2819;
      15633:data<=-16'd2816;
      15634:data<=-16'd2452;
      15635:data<=-16'd2403;
      15636:data<=-16'd2460;
      15637:data<=-16'd2024;
      15638:data<=-16'd2278;
      15639:data<=-16'd3369;
      15640:data<=-16'd4017;
      15641:data<=-16'd3362;
      15642:data<=-16'd3118;
      15643:data<=-16'd4552;
      15644:data<=-16'd5409;
      15645:data<=-16'd5372;
      15646:data<=-16'd5256;
      15647:data<=-16'd5462;
      15648:data<=-16'd6910;
      15649:data<=-16'd6893;
      15650:data<=-16'd5982;
      15651:data<=-16'd6951;
      15652:data<=-16'd6478;
      15653:data<=-16'd5940;
      15654:data<=-16'd5868;
      15655:data<=-16'd3374;
      15656:data<=-16'd7897;
      15657:data<=-16'd18403;
      15658:data<=-16'd19996;
      15659:data<=-16'd17540;
      15660:data<=-16'd18269;
      15661:data<=-16'd17229;
      15662:data<=-16'd16117;
      15663:data<=-16'd16172;
      15664:data<=-16'd15926;
      15665:data<=-16'd16607;
      15666:data<=-16'd15805;
      15667:data<=-16'd14090;
      15668:data<=-16'd13800;
      15669:data<=-16'd13300;
      15670:data<=-16'd12833;
      15671:data<=-16'd12138;
      15672:data<=-16'd11624;
      15673:data<=-16'd12589;
      15674:data<=-16'd12357;
      15675:data<=-16'd11427;
      15676:data<=-16'd11171;
      15677:data<=-16'd10113;
      15678:data<=-16'd9542;
      15679:data<=-16'd8713;
      15680:data<=-16'd7802;
      15681:data<=-16'd9465;
      15682:data<=-16'd10029;
      15683:data<=-16'd8699;
      15684:data<=-16'd8695;
      15685:data<=-16'd8125;
      15686:data<=-16'd7169;
      15687:data<=-16'd6675;
      15688:data<=-16'd5441;
      15689:data<=-16'd5486;
      15690:data<=-16'd6434;
      15691:data<=-16'd6238;
      15692:data<=-16'd5783;
      15693:data<=-16'd5318;
      15694:data<=-16'd4933;
      15695:data<=-16'd4303;
      15696:data<=-16'd2914;
      15697:data<=-16'd1306;
      15698:data<=-16'd3;
      15699:data<=-16'd832;
      15700:data<=-16'd544;
      15701:data<=16'd6454;
      15702:data<=16'd13624;
      15703:data<=16'd14252;
      15704:data<=16'd13048;
      15705:data<=16'd13326;
      15706:data<=16'd14207;
      15707:data<=16'd14833;
      15708:data<=16'd14689;
      15709:data<=16'd14354;
      15710:data<=16'd13581;
      15711:data<=16'd13214;
      15712:data<=16'd13579;
      15713:data<=16'd12907;
      15714:data<=16'd13179;
      15715:data<=16'd14781;
      15716:data<=16'd14862;
      15717:data<=16'd14445;
      15718:data<=16'd13762;
      15719:data<=16'd13018;
      15720:data<=16'd13553;
      15721:data<=16'd13135;
      15722:data<=16'd12948;
      15723:data<=16'd14298;
      15724:data<=16'd13755;
      15725:data<=16'd13113;
      15726:data<=16'd13573;
      15727:data<=16'd12715;
      15728:data<=16'd12607;
      15729:data<=16'd12875;
      15730:data<=16'd12041;
      15731:data<=16'd12348;
      15732:data<=16'd12833;
      15733:data<=16'd12710;
      15734:data<=16'd12387;
      15735:data<=16'd11241;
      15736:data<=16'd11265;
      15737:data<=16'd11394;
      15738:data<=16'd9890;
      15739:data<=16'd9976;
      15740:data<=16'd11309;
      15741:data<=16'd11679;
      15742:data<=16'd10912;
      15743:data<=16'd9797;
      15744:data<=16'd10804;
      15745:data<=16'd8355;
      15746:data<=-16'd1108;
      15747:data<=-16'd5004;
      15748:data<=-16'd1387;
      15749:data<=-16'd1400;
      15750:data<=-16'd3057;
      15751:data<=-16'd2955;
      15752:data<=-16'd3617;
      15753:data<=-16'd3071;
      15754:data<=-16'd2394;
      15755:data<=-16'd3243;
      15756:data<=-16'd2397;
      15757:data<=-16'd691;
      15758:data<=-16'd271;
      15759:data<=-16'd440;
      15760:data<=-16'd638;
      15761:data<=-16'd126;
      15762:data<=-16'd67;
      15763:data<=-16'd858;
      15764:data<=16'd86;
      15765:data<=16'd1712;
      15766:data<=16'd1880;
      15767:data<=16'd1859;
      15768:data<=16'd1779;
      15769:data<=16'd1369;
      15770:data<=16'd1532;
      15771:data<=16'd1647;
      15772:data<=16'd1657;
      15773:data<=16'd2557;
      15774:data<=16'd3260;
      15775:data<=16'd3248;
      15776:data<=16'd3712;
      15777:data<=16'd3685;
      15778:data<=16'd2940;
      15779:data<=16'd3146;
      15780:data<=16'd3133;
      15781:data<=16'd3159;
      15782:data<=16'd4821;
      15783:data<=16'd5372;
      15784:data<=16'd4918;
      15785:data<=16'd5195;
      15786:data<=16'd4317;
      15787:data<=16'd4123;
      15788:data<=16'd4146;
      15789:data<=16'd2722;
      15790:data<=16'd8135;
      15791:data<=16'd18137;
      15792:data<=16'd19576;
      15793:data<=16'd16727;
      15794:data<=16'd16971;
      15795:data<=16'd16308;
      15796:data<=16'd15027;
      15797:data<=16'd14945;
      15798:data<=16'd14985;
      15799:data<=16'd15609;
      15800:data<=16'd15179;
      15801:data<=16'd13353;
      15802:data<=16'd12856;
      15803:data<=16'd13869;
      15804:data<=16'd14624;
      15805:data<=16'd13750;
      15806:data<=16'd12834;
      15807:data<=16'd13875;
      15808:data<=16'd14697;
      15809:data<=16'd13802;
      15810:data<=16'd12355;
      15811:data<=16'd11594;
      15812:data<=16'd11477;
      15813:data<=16'd10410;
      15814:data<=16'd10034;
      15815:data<=16'd11330;
      15816:data<=16'd10824;
      15817:data<=16'd9875;
      15818:data<=16'd10370;
      15819:data<=16'd9506;
      15820:data<=16'd8128;
      15821:data<=16'd7409;
      15822:data<=16'd6974;
      15823:data<=16'd8014;
      15824:data<=16'd8595;
      15825:data<=16'd7598;
      15826:data<=16'd7047;
      15827:data<=16'd6959;
      15828:data<=16'd6777;
      15829:data<=16'd5993;
      15830:data<=16'd4966;
      15831:data<=16'd4296;
      15832:data<=16'd3853;
      15833:data<=16'd4696;
      15834:data<=16'd2033;
      15835:data<=-16'd6707;
      15836:data<=-16'd10966;
      15837:data<=-16'd9368;
      15838:data<=-16'd9935;
      15839:data<=-16'd10824;
      15840:data<=-16'd11392;
      15841:data<=-16'd12501;
      15842:data<=-16'd11468;
      15843:data<=-16'd11009;
      15844:data<=-16'd11474;
      15845:data<=-16'd10941;
      15846:data<=-16'd11007;
      15847:data<=-16'd10571;
      15848:data<=-16'd10950;
      15849:data<=-16'd12756;
      15850:data<=-16'd12508;
      15851:data<=-16'd12424;
      15852:data<=-16'd12689;
      15853:data<=-16'd11514;
      15854:data<=-16'd11603;
      15855:data<=-16'd11568;
      15856:data<=-16'd12014;
      15857:data<=-16'd14610;
      15858:data<=-16'd14888;
      15859:data<=-16'd14195;
      15860:data<=-16'd14267;
      15861:data<=-16'd12954;
      15862:data<=-16'd12919;
      15863:data<=-16'd12994;
      15864:data<=-16'd11768;
      15865:data<=-16'd12477;
      15866:data<=-16'd13204;
      15867:data<=-16'd12995;
      15868:data<=-16'd12568;
      15869:data<=-16'd11406;
      15870:data<=-16'd11627;
      15871:data<=-16'd11315;
      15872:data<=-16'd10158;
      15873:data<=-16'd11264;
      15874:data<=-16'd11864;
      15875:data<=-16'd12146;
      15876:data<=-16'd12231;
      15877:data<=-16'd10815;
      15878:data<=-16'd12057;
      15879:data<=-16'd8842;
      15880:data<=16'd1820;
      15881:data<=16'd3876;
      15882:data<=-16'd472;
      15883:data<=16'd502;
      15884:data<=16'd1113;
      15885:data<=16'd478;
      15886:data<=16'd1122;
      15887:data<=16'd100;
      15888:data<=16'd180;
      15889:data<=16'd801;
      15890:data<=-16'd901;
      15891:data<=-16'd1654;
      15892:data<=-16'd1580;
      15893:data<=-16'd1897;
      15894:data<=-16'd1369;
      15895:data<=-16'd1111;
      15896:data<=-16'd1060;
      15897:data<=-16'd496;
      15898:data<=-16'd1107;
      15899:data<=-16'd3039;
      15900:data<=-16'd3927;
      15901:data<=-16'd3201;
      15902:data<=-16'd2839;
      15903:data<=-16'd2949;
      15904:data<=-16'd2755;
      15905:data<=-16'd2989;
      15906:data<=-16'd3560;
      15907:data<=-16'd4728;
      15908:data<=-16'd5838;
      15909:data<=-16'd4751;
      15910:data<=-16'd3099;
      15911:data<=-16'd2866;
      15912:data<=-16'd3171;
      15913:data<=-16'd3055;
      15914:data<=-16'd2115;
      15915:data<=-16'd2543;
      15916:data<=-16'd4287;
      15917:data<=-16'd4273;
      15918:data<=-16'd4231;
      15919:data<=-16'd4488;
      15920:data<=-16'd3905;
      15921:data<=-16'd4206;
      15922:data<=-16'd2995;
      15923:data<=-16'd3774;
      15924:data<=-16'd12319;
      15925:data<=-16'd18283;
      15926:data<=-16'd17095;
      15927:data<=-16'd17001;
      15928:data<=-16'd16960;
      15929:data<=-16'd15582;
      15930:data<=-16'd15158;
      15931:data<=-16'd14422;
      15932:data<=-16'd15118;
      15933:data<=-16'd15973;
      15934:data<=-16'd14160;
      15935:data<=-16'd13368;
      15936:data<=-16'd13514;
      15937:data<=-16'd12859;
      15938:data<=-16'd12742;
      15939:data<=-16'd12126;
      15940:data<=-16'd12032;
      15941:data<=-16'd13086;
      15942:data<=-16'd12880;
      15943:data<=-16'd12017;
      15944:data<=-16'd11038;
      15945:data<=-16'd10414;
      15946:data<=-16'd10366;
      15947:data<=-16'd9034;
      15948:data<=-16'd8940;
      15949:data<=-16'd10800;
      15950:data<=-16'd10589;
      15951:data<=-16'd9697;
      15952:data<=-16'd9435;
      15953:data<=-16'd8492;
      15954:data<=-16'd7827;
      15955:data<=-16'd6993;
      15956:data<=-16'd6555;
      15957:data<=-16'd7407;
      15958:data<=-16'd7724;
      15959:data<=-16'd7650;
      15960:data<=-16'd7080;
      15961:data<=-16'd6193;
      15962:data<=-16'd6610;
      15963:data<=-16'd7100;
      15964:data<=-16'd7330;
      15965:data<=-16'd6711;
      15966:data<=-16'd5711;
      15967:data<=-16'd7127;
      15968:data<=-16'd3714;
      15969:data<=16'd6149;
      15970:data<=16'd9071;
      15971:data<=16'd7084;
      15972:data<=16'd8525;
      15973:data<=16'd8802;
      15974:data<=16'd8910;
      15975:data<=16'd10348;
      15976:data<=16'd9406;
      15977:data<=16'd8860;
      15978:data<=16'd9204;
      15979:data<=16'd8893;
      15980:data<=16'd9004;
      15981:data<=16'd8414;
      15982:data<=16'd9133;
      15983:data<=16'd11009;
      15984:data<=16'd10551;
      15985:data<=16'd10361;
      15986:data<=16'd10449;
      15987:data<=16'd9483;
      15988:data<=16'd9577;
      15989:data<=16'd8763;
      15990:data<=16'd8431;
      15991:data<=16'd10810;
      15992:data<=16'd11342;
      15993:data<=16'd10499;
      15994:data<=16'd10481;
      15995:data<=16'd9973;
      15996:data<=16'd9865;
      15997:data<=16'd9106;
      15998:data<=16'd8323;
      15999:data<=16'd9991;
      16000:data<=16'd10954;
      16001:data<=16'd10420;
      16002:data<=16'd10058;
      16003:data<=16'd9365;
      16004:data<=16'd9436;
      16005:data<=16'd9251;
      16006:data<=16'd8150;
      16007:data<=16'd8416;
      16008:data<=16'd9429;
      16009:data<=16'd10132;
      16010:data<=16'd9477;
      16011:data<=16'd8636;
      16012:data<=16'd9464;
      16013:data<=16'd4582;
      16014:data<=-16'd4948;
      16015:data<=-16'd5548;
      16016:data<=-16'd866;
      16017:data<=-16'd349;
      16018:data<=-16'd349;
      16019:data<=-16'd123;
      16020:data<=-16'd558;
      16021:data<=-16'd32;
      16022:data<=-16'd517;
      16023:data<=-16'd617;
      16024:data<=16'd1321;
      16025:data<=16'd2303;
      16026:data<=16'd1911;
      16027:data<=16'd1148;
      16028:data<=16'd858;
      16029:data<=16'd1598;
      16030:data<=16'd1521;
      16031:data<=16'd995;
      16032:data<=16'd2036;
      16033:data<=16'd3739;
      16034:data<=16'd4431;
      16035:data<=16'd3946;
      16036:data<=16'd3519;
      16037:data<=16'd3451;
      16038:data<=16'd2723;
      16039:data<=16'd2071;
      16040:data<=16'd2905;
      16041:data<=16'd4675;
      16042:data<=16'd5457;
      16043:data<=16'd5133;
      16044:data<=16'd5036;
      16045:data<=16'd4540;
      16046:data<=16'd4027;
      16047:data<=16'd4156;
      16048:data<=16'd3573;
      16049:data<=16'd4030;
      16050:data<=16'd5577;
      16051:data<=16'd5598;
      16052:data<=16'd5762;
      16053:data<=16'd5745;
      16054:data<=16'd5227;
      16055:data<=16'd5075;
      16056:data<=16'd2945;
      16057:data<=16'd5974;
      16058:data<=16'd16575;
      16059:data<=16'd20113;
      16060:data<=16'd17547;
      16061:data<=16'd18117;
      16062:data<=16'd17250;
      16063:data<=16'd15835;
      16064:data<=16'd15722;
      16065:data<=16'd14454;
      16066:data<=16'd15669;
      16067:data<=16'd16575;
      16068:data<=16'd14125;
      16069:data<=16'd12701;
      16070:data<=16'd11611;
      16071:data<=16'd11192;
      16072:data<=16'd11314;
      16073:data<=16'd9403;
      16074:data<=16'd9535;
      16075:data<=16'd10780;
      16076:data<=16'd9993;
      16077:data<=16'd10182;
      16078:data<=16'd9451;
      16079:data<=16'd7938;
      16080:data<=16'd8188;
      16081:data<=16'd7641;
      16082:data<=16'd7964;
      16083:data<=16'd9153;
      16084:data<=16'd8387;
      16085:data<=16'd8126;
      16086:data<=16'd7844;
      16087:data<=16'd7018;
      16088:data<=16'd6818;
      16089:data<=16'd5644;
      16090:data<=16'd5844;
      16091:data<=16'd7250;
      16092:data<=16'd6886;
      16093:data<=16'd6660;
      16094:data<=16'd5935;
      16095:data<=16'd5210;
      16096:data<=16'd5718;
      16097:data<=16'd4698;
      16098:data<=16'd4493;
      16099:data<=16'd4681;
      16100:data<=16'd3648;
      16101:data<=16'd5218;
      16102:data<=16'd1654;
      16103:data<=-16'd8781;
      16104:data<=-16'd11588;
      16105:data<=-16'd9136;
      16106:data<=-16'd9693;
      16107:data<=-16'd9809;
      16108:data<=-16'd10349;
      16109:data<=-16'd11218;
      16110:data<=-16'd10534;
      16111:data<=-16'd10777;
      16112:data<=-16'd10618;
      16113:data<=-16'd10014;
      16114:data<=-16'd9909;
      16115:data<=-16'd8866;
      16116:data<=-16'd9784;
      16117:data<=-16'd11770;
      16118:data<=-16'd11273;
      16119:data<=-16'd10730;
      16120:data<=-16'd10351;
      16121:data<=-16'd9339;
      16122:data<=-16'd8314;
      16123:data<=-16'd6554;
      16124:data<=-16'd6734;
      16125:data<=-16'd8758;
      16126:data<=-16'd8910;
      16127:data<=-16'd8658;
      16128:data<=-16'd8699;
      16129:data<=-16'd8137;
      16130:data<=-16'd7912;
      16131:data<=-16'd7169;
      16132:data<=-16'd6946;
      16133:data<=-16'd8455;
      16134:data<=-16'd9027;
      16135:data<=-16'd8307;
      16136:data<=-16'd7812;
      16137:data<=-16'd7732;
      16138:data<=-16'd7912;
      16139:data<=-16'd7351;
      16140:data<=-16'd6307;
      16141:data<=-16'd6687;
      16142:data<=-16'd8334;
      16143:data<=-16'd8352;
      16144:data<=-16'd7010;
      16145:data<=-16'd8055;
      16146:data<=-16'd6874;
      16147:data<=16'd1528;
      16148:data<=16'd7617;
      16149:data<=16'd6423;
      16150:data<=16'd4777;
      16151:data<=16'd3798;
      16152:data<=16'd3013;
      16153:data<=16'd3624;
      16154:data<=16'd3541;
      16155:data<=16'd3341;
      16156:data<=16'd3635;
      16157:data<=16'd2805;
      16158:data<=16'd1545;
      16159:data<=16'd479;
      16160:data<=16'd473;
      16161:data<=16'd1351;
      16162:data<=16'd1014;
      16163:data<=16'd431;
      16164:data<=16'd676;
      16165:data<=16'd992;
      16166:data<=16'd200;
      16167:data<=-16'd2134;
      16168:data<=-16'd2378;
      16169:data<=-16'd823;
      16170:data<=-16'd1351;
      16171:data<=-16'd1401;
      16172:data<=-16'd608;
      16173:data<=-16'd864;
      16174:data<=-16'd883;
      16175:data<=-16'd3043;
      16176:data<=-16'd5937;
      16177:data<=-16'd5410;
      16178:data<=-16'd4605;
      16179:data<=-16'd4541;
      16180:data<=-16'd4266;
      16181:data<=-16'd4118;
      16182:data<=-16'd3330;
      16183:data<=-16'd4435;
      16184:data<=-16'd5826;
      16185:data<=-16'd4902;
      16186:data<=-16'd5283;
      16187:data<=-16'd4958;
      16188:data<=-16'd4162;
      16189:data<=-16'd4948;
      16190:data<=-16'd2645;
      16191:data<=-16'd5633;
      16192:data<=-16'd16853;
      16193:data<=-16'd19725;
      16194:data<=-16'd16917;
      16195:data<=-16'd17673;
      16196:data<=-16'd16313;
      16197:data<=-16'd14932;
      16198:data<=-16'd14894;
      16199:data<=-16'd13443;
      16200:data<=-16'd14557;
      16201:data<=-16'd15481;
      16202:data<=-16'd14142;
      16203:data<=-16'd13894;
      16204:data<=-16'd12734;
      16205:data<=-16'd11982;
      16206:data<=-16'd12143;
      16207:data<=-16'd10630;
      16208:data<=-16'd10937;
      16209:data<=-16'd12085;
      16210:data<=-16'd11253;
      16211:data<=-16'd10586;
      16212:data<=-16'd9371;
      16213:data<=-16'd8865;
      16214:data<=-16'd9494;
      16215:data<=-16'd8281;
      16216:data<=-16'd8197;
      16217:data<=-16'd9547;
      16218:data<=-16'd9336;
      16219:data<=-16'd9204;
      16220:data<=-16'd8560;
      16221:data<=-16'd7344;
      16222:data<=-16'd6893;
      16223:data<=-16'd5938;
      16224:data<=-16'd6062;
      16225:data<=-16'd7066;
      16226:data<=-16'd6996;
      16227:data<=-16'd7109;
      16228:data<=-16'd5720;
      16229:data<=-16'd3294;
      16230:data<=-16'd3008;
      16231:data<=-16'd2969;
      16232:data<=-16'd2558;
      16233:data<=-16'd2146;
      16234:data<=-16'd1773;
      16235:data<=-16'd1632;
      16236:data<=16'd3642;
      16237:data<=16'd11455;
      16238:data<=16'd12475;
      16239:data<=16'd11206;
      16240:data<=16'd11944;
      16241:data<=16'd11591;
      16242:data<=16'd12199;
      16243:data<=16'd12995;
      16244:data<=16'd12296;
      16245:data<=16'd12508;
      16246:data<=16'd11993;
      16247:data<=16'd10930;
      16248:data<=16'd11130;
      16249:data<=16'd11189;
      16250:data<=16'd12088;
      16251:data<=16'd13004;
      16252:data<=16'd12281;
      16253:data<=16'd11941;
      16254:data<=16'd11643;
      16255:data<=16'd11192;
      16256:data<=16'd10834;
      16257:data<=16'd9693;
      16258:data<=16'd10445;
      16259:data<=16'd12248;
      16260:data<=16'd11735;
      16261:data<=16'd11132;
      16262:data<=16'd11074;
      16263:data<=16'd10840;
      16264:data<=16'd10821;
      16265:data<=16'd9508;
      16266:data<=16'd9068;
      16267:data<=16'd10887;
      16268:data<=16'd11060;
      16269:data<=16'd10090;
      16270:data<=16'd10367;
      16271:data<=16'd10345;
      16272:data<=16'd9630;
      16273:data<=16'd9286;
      16274:data<=16'd9010;
      16275:data<=16'd9048;
      16276:data<=16'd10241;
      16277:data<=16'd10329;
      16278:data<=16'd8912;
      16279:data<=16'd9471;
      16280:data<=16'd6968;
      16281:data<=-16'd2494;
      16282:data<=-16'd8193;
      16283:data<=-16'd6699;
      16284:data<=-16'd5303;
      16285:data<=-16'd4499;
      16286:data<=-16'd4175;
      16287:data<=-16'd4564;
      16288:data<=-16'd3727;
      16289:data<=-16'd3852;
      16290:data<=-16'd4422;
      16291:data<=-16'd3016;
      16292:data<=-16'd1830;
      16293:data<=-16'd1348;
      16294:data<=-16'd1010;
      16295:data<=-16'd1307;
      16296:data<=-16'd1513;
      16297:data<=-16'd1486;
      16298:data<=-16'd1290;
      16299:data<=-16'd1392;
      16300:data<=-16'd966;
      16301:data<=16'd1224;
      16302:data<=16'd2108;
      16303:data<=16'd1169;
      16304:data<=16'd925;
      16305:data<=16'd711;
      16306:data<=16'd789;
      16307:data<=16'd587;
      16308:data<=16'd221;
      16309:data<=16'd2265;
      16310:data<=16'd3500;
      16311:data<=16'd3015;
      16312:data<=16'd3615;
      16313:data<=16'd2817;
      16314:data<=16'd2070;
      16315:data<=16'd2470;
      16316:data<=16'd1610;
      16317:data<=16'd2972;
      16318:data<=16'd4434;
      16319:data<=16'd3077;
      16320:data<=16'd3436;
      16321:data<=16'd3303;
      16322:data<=16'd2968;
      16323:data<=16'd3879;
      16324:data<=16'd1425;
      16325:data<=16'd4860;
      16326:data<=16'd16096;
      16327:data<=16'd18542;
      16328:data<=16'd15396;
      16329:data<=16'd15955;
      16330:data<=16'd15449;
      16331:data<=16'd14504;
      16332:data<=16'd14002;
      16333:data<=16'd13035;
      16334:data<=16'd14425;
      16335:data<=16'd15726;
      16336:data<=16'd15722;
      16337:data<=16'd15239;
      16338:data<=16'd13380;
      16339:data<=16'd13065;
      16340:data<=16'd13321;
      16341:data<=16'd12170;
      16342:data<=16'd12402;
      16343:data<=16'd12537;
      16344:data<=16'd11972;
      16345:data<=16'd11841;
      16346:data<=16'd10719;
      16347:data<=16'd10331;
      16348:data<=16'd9976;
      16349:data<=16'd8642;
      16350:data<=16'd9400;
      16351:data<=16'd10125;
      16352:data<=16'd9741;
      16353:data<=16'd9873;
      16354:data<=16'd8661;
      16355:data<=16'd7812;
      16356:data<=16'd7523;
      16357:data<=16'd5823;
      16358:data<=16'd5999;
      16359:data<=16'd7421;
      16360:data<=16'd7694;
      16361:data<=16'd7679;
      16362:data<=16'd6455;
      16363:data<=16'd5450;
      16364:data<=16'd5492;
      16365:data<=16'd4886;
      16366:data<=16'd4290;
      16367:data<=16'd3594;
      16368:data<=16'd3771;
      16369:data<=16'd2038;
      16370:data<=-16'd6152;
      16371:data<=-16'd11785;
      16372:data<=-16'd10607;
      16373:data<=-16'd10643;
      16374:data<=-16'd10699;
      16375:data<=-16'd10343;
      16376:data<=-16'd12319;
      16377:data<=-16'd12260;
      16378:data<=-16'd11533;
      16379:data<=-16'd12008;
      16380:data<=-16'd11041;
      16381:data<=-16'd10919;
      16382:data<=-16'd10937;
      16383:data<=-16'd10367;
      16384:data<=-16'd11929;
      16385:data<=-16'd12609;
      16386:data<=-16'd12073;
      16387:data<=-16'd12759;
      16388:data<=-16'd12874;
      16389:data<=-16'd12819;
      16390:data<=-16'd12624;
      16391:data<=-16'd11837;
      16392:data<=-16'd12551;
      16393:data<=-16'd13658;
      16394:data<=-16'd13850;
      16395:data<=-16'd13621;
      16396:data<=-16'd12979;
      16397:data<=-16'd12922;
      16398:data<=-16'd12666;
      16399:data<=-16'd11618;
      16400:data<=-16'd11424;
      16401:data<=-16'd12087;
      16402:data<=-16'd13001;
      16403:data<=-16'd13089;
      16404:data<=-16'd12310;
      16405:data<=-16'd12158;
      16406:data<=-16'd11809;
      16407:data<=-16'd11392;
      16408:data<=-16'd11227;
      16409:data<=-16'd11036;
      16410:data<=-16'd12352;
      16411:data<=-16'd11981;
      16412:data<=-16'd10188;
      16413:data<=-16'd11790;
      16414:data<=-16'd8619;
      16415:data<=16'd1149;
      16416:data<=16'd4250;
      16417:data<=16'd2220;
      16418:data<=16'd2059;
      16419:data<=16'd933;
      16420:data<=16'd488;
      16421:data<=16'd1439;
      16422:data<=16'd540;
      16423:data<=16'd80;
      16424:data<=16'd751;
      16425:data<=16'd27;
      16426:data<=-16'd1515;
      16427:data<=-16'd2314;
      16428:data<=-16'd2083;
      16429:data<=-16'd1727;
      16430:data<=-16'd1844;
      16431:data<=-16'd2015;
      16432:data<=-16'd1636;
      16433:data<=-16'd1221;
      16434:data<=-16'd2746;
      16435:data<=-16'd4813;
      16436:data<=-16'd4513;
      16437:data<=-16'd3506;
      16438:data<=-16'd3259;
      16439:data<=-16'd3574;
      16440:data<=-16'd3694;
      16441:data<=-16'd1691;
      16442:data<=-16'd646;
      16443:data<=-16'd2886;
      16444:data<=-16'd3894;
      16445:data<=-16'd3421;
      16446:data<=-16'd3671;
      16447:data<=-16'd3491;
      16448:data<=-16'd3280;
      16449:data<=-16'd2787;
      16450:data<=-16'd2426;
      16451:data<=-16'd3738;
      16452:data<=-16'd4300;
      16453:data<=-16'd4081;
      16454:data<=-16'd4467;
      16455:data<=-16'd3874;
      16456:data<=-16'd3606;
      16457:data<=-16'd3312;
      16458:data<=-16'd3500;
      16459:data<=-16'd10019;
      16460:data<=-16'd17697;
      16461:data<=-16'd18064;
      16462:data<=-16'd16763;
      16463:data<=-16'd17183;
      16464:data<=-16'd16205;
      16465:data<=-16'd15168;
      16466:data<=-16'd14554;
      16467:data<=-16'd14213;
      16468:data<=-16'd14989;
      16469:data<=-16'd14842;
      16470:data<=-16'd13705;
      16471:data<=-16'd13185;
      16472:data<=-16'd12656;
      16473:data<=-16'd11887;
      16474:data<=-16'd11116;
      16475:data<=-16'd10886;
      16476:data<=-16'd11461;
      16477:data<=-16'd11759;
      16478:data<=-16'd11626;
      16479:data<=-16'd10892;
      16480:data<=-16'd9777;
      16481:data<=-16'd9511;
      16482:data<=-16'd8943;
      16483:data<=-16'd8023;
      16484:data<=-16'd8592;
      16485:data<=-16'd9300;
      16486:data<=-16'd9182;
      16487:data<=-16'd8948;
      16488:data<=-16'd8111;
      16489:data<=-16'd7266;
      16490:data<=-16'd7016;
      16491:data<=-16'd6613;
      16492:data<=-16'd6470;
      16493:data<=-16'd7432;
      16494:data<=-16'd8526;
      16495:data<=-16'd8431;
      16496:data<=-16'd8144;
      16497:data<=-16'd7944;
      16498:data<=-16'd7103;
      16499:data<=-16'd7074;
      16500:data<=-16'd6304;
      16501:data<=-16'd4855;
      16502:data<=-16'd6291;
      16503:data<=-16'd2905;
      16504:data<=16'd7272;
      16505:data<=16'd10217;
      16506:data<=16'd8328;
      16507:data<=16'd10143;
      16508:data<=16'd9626;
      16509:data<=16'd9145;
      16510:data<=16'd11771;
      16511:data<=16'd11104;
      16512:data<=16'd10231;
      16513:data<=16'd11115;
      16514:data<=16'd10149;
      16515:data<=16'd9741;
      16516:data<=16'd9515;
      16517:data<=16'd9327;
      16518:data<=16'd11213;
      16519:data<=16'd11677;
      16520:data<=16'd10962;
      16521:data<=16'd11112;
      16522:data<=16'd10634;
      16523:data<=16'd10615;
      16524:data<=16'd10205;
      16525:data<=16'd9086;
      16526:data<=16'd10255;
      16527:data<=16'd11637;
      16528:data<=16'd11544;
      16529:data<=16'd11436;
      16530:data<=16'd10865;
      16531:data<=16'd10539;
      16532:data<=16'd10540;
      16533:data<=16'd9808;
      16534:data<=16'd9734;
      16535:data<=16'd10985;
      16536:data<=16'd11982;
      16537:data<=16'd11364;
      16538:data<=16'd10466;
      16539:data<=16'd10348;
      16540:data<=16'd9599;
      16541:data<=16'd9386;
      16542:data<=16'd9966;
      16543:data<=16'd10275;
      16544:data<=16'd11664;
      16545:data<=16'd11035;
      16546:data<=16'd9420;
      16547:data<=16'd11526;
      16548:data<=16'd8443;
      16549:data<=-16'd872;
      16550:data<=-16'd3080;
      16551:data<=-16'd329;
      16552:data<=16'd402;
      16553:data<=16'd917;
      16554:data<=16'd529;
      16555:data<=16'd143;
      16556:data<=16'd813;
      16557:data<=16'd607;
      16558:data<=16'd640;
      16559:data<=16'd1483;
      16560:data<=16'd3054;
      16561:data<=16'd4338;
      16562:data<=16'd3347;
      16563:data<=16'd2758;
      16564:data<=16'd3259;
      16565:data<=16'd3254;
      16566:data<=16'd3673;
      16567:data<=16'd3460;
      16568:data<=16'd3997;
      16569:data<=16'd5800;
      16570:data<=16'd5324;
      16571:data<=16'd5016;
      16572:data<=16'd5491;
      16573:data<=16'd4522;
      16574:data<=16'd4763;
      16575:data<=16'd4617;
      16576:data<=16'd3940;
      16577:data<=16'd5879;
      16578:data<=16'd6815;
      16579:data<=16'd6358;
      16580:data<=16'd6328;
      16581:data<=16'd5335;
      16582:data<=16'd5036;
      16583:data<=16'd4681;
      16584:data<=16'd4422;
      16585:data<=16'd6226;
      16586:data<=16'd6507;
      16587:data<=16'd5976;
      16588:data<=16'd6300;
      16589:data<=16'd5697;
      16590:data<=16'd5733;
      16591:data<=16'd4455;
      16592:data<=16'd5762;
      16593:data<=16'd15555;
      16594:data<=16'd21140;
      16595:data<=16'd18742;
      16596:data<=16'd18666;
      16597:data<=16'd17858;
      16598:data<=16'd16095;
      16599:data<=16'd16927;
      16600:data<=16'd15364;
      16601:data<=16'd13782;
      16602:data<=16'd14721;
      16603:data<=16'd14273;
      16604:data<=16'd13227;
      16605:data<=16'd12041;
      16606:data<=16'd11309;
      16607:data<=16'd11630;
      16608:data<=16'd10516;
      16609:data<=16'd10072;
      16610:data<=16'd10937;
      16611:data<=16'd10625;
      16612:data<=16'd10843;
      16613:data<=16'd10642;
      16614:data<=16'd9315;
      16615:data<=16'd9289;
      16616:data<=16'd8648;
      16617:data<=16'd7244;
      16618:data<=16'd7638;
      16619:data<=16'd8584;
      16620:data<=16'd8710;
      16621:data<=16'd8134;
      16622:data<=16'd7504;
      16623:data<=16'd7225;
      16624:data<=16'd6801;
      16625:data<=16'd6419;
      16626:data<=16'd6191;
      16627:data<=16'd6768;
      16628:data<=16'd7715;
      16629:data<=16'd7115;
      16630:data<=16'd6649;
      16631:data<=16'd6455;
      16632:data<=16'd5294;
      16633:data<=16'd5773;
      16634:data<=16'd5415;
      16635:data<=16'd3654;
      16636:data<=16'd5025;
      16637:data<=16'd1668;
      16638:data<=-16'd8384;
      16639:data<=-16'd11353;
      16640:data<=-16'd9159;
      16641:data<=-16'd10210;
      16642:data<=-16'd10100;
      16643:data<=-16'd9925;
      16644:data<=-16'd12389;
      16645:data<=-16'd12637;
      16646:data<=-16'd11724;
      16647:data<=-16'd11858;
      16648:data<=-16'd10985;
      16649:data<=-16'd10342;
      16650:data<=-16'd10034;
      16651:data<=-16'd9658;
      16652:data<=-16'd11213;
      16653:data<=-16'd11653;
      16654:data<=-16'd9479;
      16655:data<=-16'd8965;
      16656:data<=-16'd9010;
      16657:data<=-16'd7931;
      16658:data<=-16'd8046;
      16659:data<=-16'd8052;
      16660:data<=-16'd8072;
      16661:data<=-16'd9448;
      16662:data<=-16'd9382;
      16663:data<=-16'd8830;
      16664:data<=-16'd9216;
      16665:data<=-16'd8542;
      16666:data<=-16'd8357;
      16667:data<=-16'd8310;
      16668:data<=-16'd7630;
      16669:data<=-16'd9247;
      16670:data<=-16'd9999;
      16671:data<=-16'd8502;
      16672:data<=-16'd8909;
      16673:data<=-16'd8921;
      16674:data<=-16'd8229;
      16675:data<=-16'd8940;
      16676:data<=-16'd8555;
      16677:data<=-16'd9183;
      16678:data<=-16'd10358;
      16679:data<=-16'd8869;
      16680:data<=-16'd9341;
      16681:data<=-16'd8093;
      16682:data<=16'd5;
      16683:data<=16'd4992;
      16684:data<=16'd4617;
      16685:data<=16'd4643;
      16686:data<=16'd3269;
      16687:data<=16'd2035;
      16688:data<=16'd2925;
      16689:data<=16'd3080;
      16690:data<=16'd2890;
      16691:data<=16'd2732;
      16692:data<=16'd2476;
      16693:data<=16'd1977;
      16694:data<=-16'd230;
      16695:data<=-16'd1372;
      16696:data<=-16'd531;
      16697:data<=-16'd508;
      16698:data<=-16'd429;
      16699:data<=-16'd778;
      16700:data<=-16'd1560;
      16701:data<=-16'd966;
      16702:data<=-16'd1882;
      16703:data<=-16'd3885;
      16704:data<=-16'd3894;
      16705:data<=-16'd3635;
      16706:data<=-16'd3770;
      16707:data<=-16'd4766;
      16708:data<=-16'd6050;
      16709:data<=-16'd4958;
      16710:data<=-16'd4561;
      16711:data<=-16'd6243;
      16712:data<=-16'd6626;
      16713:data<=-16'd6282;
      16714:data<=-16'd5714;
      16715:data<=-16'd5154;
      16716:data<=-16'd5125;
      16717:data<=-16'd4311;
      16718:data<=-16'd4683;
      16719:data<=-16'd5930;
      16720:data<=-16'd5791;
      16721:data<=-16'd6117;
      16722:data<=-16'd5547;
      16723:data<=-16'd4987;
      16724:data<=-16'd5943;
      16725:data<=-16'd4120;
      16726:data<=-16'd6927;
      16727:data<=-16'd17569;
      16728:data<=-16'd20745;
      16729:data<=-16'd17873;
      16730:data<=-16'd18777;
      16731:data<=-16'd18230;
      16732:data<=-16'd16775;
      16733:data<=-16'd16744;
      16734:data<=-16'd15039;
      16735:data<=-16'd15531;
      16736:data<=-16'd17500;
      16737:data<=-16'd16463;
      16738:data<=-16'd15244;
      16739:data<=-16'd14446;
      16740:data<=-16'd13540;
      16741:data<=-16'd13468;
      16742:data<=-16'd12565;
      16743:data<=-16'd11755;
      16744:data<=-16'd12363;
      16745:data<=-16'd12839;
      16746:data<=-16'd12587;
      16747:data<=-16'd11359;
      16748:data<=-16'd10123;
      16749:data<=-16'd10040;
      16750:data<=-16'd9627;
      16751:data<=-16'd8519;
      16752:data<=-16'd8523;
      16753:data<=-16'd9735;
      16754:data<=-16'd9949;
      16755:data<=-16'd8997;
      16756:data<=-16'd8684;
      16757:data<=-16'd8106;
      16758:data<=-16'd7016;
      16759:data<=-16'd6388;
      16760:data<=-16'd5277;
      16761:data<=-16'd5281;
      16762:data<=-16'd6213;
      16763:data<=-16'd5054;
      16764:data<=-16'd4554;
      16765:data<=-16'd5184;
      16766:data<=-16'd4109;
      16767:data<=-16'd3503;
      16768:data<=-16'd3215;
      16769:data<=-16'd3039;
      16770:data<=-16'd3186;
      16771:data<=16'd2743;
      16772:data<=16'd11094;
      16773:data<=16'd11524;
      16774:data<=16'd9715;
      16775:data<=16'd11195;
      16776:data<=16'd11326;
      16777:data<=16'd11347;
      16778:data<=16'd12922;
      16779:data<=16'd13038;
      16780:data<=16'd12489;
      16781:data<=16'd12389;
      16782:data<=16'd11844;
      16783:data<=16'd11323;
      16784:data<=16'd10806;
      16785:data<=16'd10784;
      16786:data<=16'd12239;
      16787:data<=16'd13214;
      16788:data<=16'd12543;
      16789:data<=16'd11888;
      16790:data<=16'd11712;
      16791:data<=16'd11699;
      16792:data<=16'd11145;
      16793:data<=16'd9906;
      16794:data<=16'd10470;
      16795:data<=16'd12034;
      16796:data<=16'd11744;
      16797:data<=16'd11229;
      16798:data<=16'd10622;
      16799:data<=16'd9734;
      16800:data<=16'd10390;
      16801:data<=16'd9823;
      16802:data<=16'd8834;
      16803:data<=16'd10613;
      16804:data<=16'd10765;
      16805:data<=16'd10058;
      16806:data<=16'd11215;
      16807:data<=16'd10100;
      16808:data<=16'd9059;
      16809:data<=16'd9458;
      16810:data<=16'd8608;
      16811:data<=16'd10378;
      16812:data<=16'd11189;
      16813:data<=16'd8152;
      16814:data<=16'd8498;
      16815:data<=16'd5871;
      16816:data<=-16'd3617;
      16817:data<=-16'd7503;
      16818:data<=-16'd6393;
      16819:data<=-16'd6184;
      16820:data<=-16'd4452;
      16821:data<=-16'd3871;
      16822:data<=-16'd4796;
      16823:data<=-16'd4215;
      16824:data<=-16'd3870;
      16825:data<=-16'd3644;
      16826:data<=-16'd3573;
      16827:data<=-16'd3271;
      16828:data<=-16'd963;
      16829:data<=-16'd135;
      16830:data<=-16'd1102;
      16831:data<=-16'd890;
      16832:data<=-16'd1027;
      16833:data<=-16'd1004;
      16834:data<=-16'd717;
      16835:data<=-16'd1131;
      16836:data<=16'd434;
      16837:data<=16'd2188;
      16838:data<=16'd1839;
      16839:data<=16'd1838;
      16840:data<=16'd1723;
      16841:data<=16'd1307;
      16842:data<=16'd1307;
      16843:data<=16'd967;
      16844:data<=16'd1707;
      16845:data<=16'd2883;
      16846:data<=16'd3263;
      16847:data<=16'd3588;
      16848:data<=16'd2816;
      16849:data<=16'd2488;
      16850:data<=16'd2769;
      16851:data<=16'd1574;
      16852:data<=16'd2366;
      16853:data<=16'd4064;
      16854:data<=16'd3512;
      16855:data<=16'd3868;
      16856:data<=16'd3486;
      16857:data<=16'd2443;
      16858:data<=16'd2910;
      16859:data<=16'd1253;
      16860:data<=16'd4623;
      16861:data<=16'd15399;
      16862:data<=16'd18412;
      16863:data<=16'd15873;
      16864:data<=16'd16780;
      16865:data<=16'd15383;
      16866:data<=16'd14383;
      16867:data<=16'd16609;
      16868:data<=16'd15867;
      16869:data<=16'd15226;
      16870:data<=16'd16333;
      16871:data<=16'd15380;
      16872:data<=16'd14615;
      16873:data<=16'd14424;
      16874:data<=16'd13509;
      16875:data<=16'd12531;
      16876:data<=16'd11233;
      16877:data<=16'd11543;
      16878:data<=16'd12850;
      16879:data<=16'd12269;
      16880:data<=16'd11539;
      16881:data<=16'd10927;
      16882:data<=16'd9799;
      16883:data<=16'd9797;
      16884:data<=16'd9298;
      16885:data<=16'd8146;
      16886:data<=16'd8939;
      16887:data<=16'd9865;
      16888:data<=16'd9260;
      16889:data<=16'd8464;
      16890:data<=16'd7708;
      16891:data<=16'd7333;
      16892:data<=16'd7157;
      16893:data<=16'd6012;
      16894:data<=16'd5588;
      16895:data<=16'd6919;
      16896:data<=16'd7404;
      16897:data<=16'd6807;
      16898:data<=16'd6481;
      16899:data<=16'd5903;
      16900:data<=16'd5677;
      16901:data<=16'd5426;
      16902:data<=16'd4443;
      16903:data<=16'd4593;
      16904:data<=16'd2347;
      16905:data<=-16'd5335;
      16906:data<=-16'd10402;
      16907:data<=-16'd9773;
      16908:data<=-16'd9711;
      16909:data<=-16'd10129;
      16910:data<=-16'd9274;
      16911:data<=-16'd9859;
      16912:data<=-16'd11445;
      16913:data<=-16'd11715;
      16914:data<=-16'd10986;
      16915:data<=-16'd10510;
      16916:data<=-16'd10584;
      16917:data<=-16'd10167;
      16918:data<=-16'd9395;
      16919:data<=-16'd10399;
      16920:data<=-16'd12925;
      16921:data<=-16'd13894;
      16922:data<=-16'd13051;
      16923:data<=-16'd12748;
      16924:data<=-16'd12766;
      16925:data<=-16'd11987;
      16926:data<=-16'd10986;
      16927:data<=-16'd10836;
      16928:data<=-16'd12185;
      16929:data<=-16'd13057;
      16930:data<=-16'd12413;
      16931:data<=-16'd12361;
      16932:data<=-16'd11788;
      16933:data<=-16'd10583;
      16934:data<=-16'd10912;
      16935:data<=-16'd10308;
      16936:data<=-16'd10099;
      16937:data<=-16'd12425;
      16938:data<=-16'd12129;
      16939:data<=-16'd10680;
      16940:data<=-16'd11215;
      16941:data<=-16'd10273;
      16942:data<=-16'd9873;
      16943:data<=-16'd10196;
      16944:data<=-16'd9297;
      16945:data<=-16'd10997;
      16946:data<=-16'd11411;
      16947:data<=-16'd9571;
      16948:data<=-16'd11465;
      16949:data<=-16'd7971;
      16950:data<=16'd2378;
      16951:data<=16'd4817;
      16952:data<=16'd2638;
      16953:data<=16'd3397;
      16954:data<=16'd2177;
      16955:data<=16'd823;
      16956:data<=16'd1536;
      16957:data<=16'd980;
      16958:data<=16'd986;
      16959:data<=16'd2099;
      16960:data<=16'd1823;
      16961:data<=16'd585;
      16962:data<=-16'd735;
      16963:data<=-16'd1210;
      16964:data<=-16'd822;
      16965:data<=-16'd904;
      16966:data<=-16'd1177;
      16967:data<=-16'd954;
      16968:data<=-16'd469;
      16969:data<=-16'd926;
      16970:data<=-16'd2840;
      16971:data<=-16'd3888;
      16972:data<=-16'd2928;
      16973:data<=-16'd1160;
      16974:data<=16'd152;
      16975:data<=-16'd347;
      16976:data<=-16'd1037;
      16977:data<=-16'd323;
      16978:data<=-16'd802;
      16979:data<=-16'd2349;
      16980:data<=-16'd2716;
      16981:data<=-16'd2657;
      16982:data<=-16'd2473;
      16983:data<=-16'd2165;
      16984:data<=-16'd1792;
      16985:data<=-16'd1240;
      16986:data<=-16'd2023;
      16987:data<=-16'd3069;
      16988:data<=-16'd2860;
      16989:data<=-16'd3015;
      16990:data<=-16'd2955;
      16991:data<=-16'd2532;
      16992:data<=-16'd2417;
      16993:data<=-16'd2742;
      16994:data<=-16'd8255;
      16995:data<=-16'd16199;
      16996:data<=-16'd17029;
      16997:data<=-16'd15276;
      16998:data<=-16'd15920;
      16999:data<=-16'd14522;
      17000:data<=-16'd13368;
      17001:data<=-16'd13479;
      17002:data<=-16'd12011;
      17003:data<=-16'd12569;
      17004:data<=-16'd14211;
      17005:data<=-16'd13110;
      17006:data<=-16'd11899;
      17007:data<=-16'd11338;
      17008:data<=-16'd10707;
      17009:data<=-16'd10511;
      17010:data<=-16'd9917;
      17011:data<=-16'd9873;
      17012:data<=-16'd10540;
      17013:data<=-16'd10366;
      17014:data<=-16'd9894;
      17015:data<=-16'd9085;
      17016:data<=-16'd7909;
      17017:data<=-16'd7382;
      17018:data<=-16'd7057;
      17019:data<=-16'd7080;
      17020:data<=-16'd7762;
      17021:data<=-16'd8229;
      17022:data<=-16'd8476;
      17023:data<=-16'd7975;
      17024:data<=-16'd6446;
      17025:data<=-16'd6401;
      17026:data<=-16'd7774;
      17027:data<=-16'd7357;
      17028:data<=-16'd6905;
      17029:data<=-16'd8423;
      17030:data<=-16'd8355;
      17031:data<=-16'd7307;
      17032:data<=-16'd7603;
      17033:data<=-16'd6802;
      17034:data<=-16'd6175;
      17035:data<=-16'd6096;
      17036:data<=-16'd4778;
      17037:data<=-16'd5380;
      17038:data<=-16'd2554;
      17039:data<=16'd7080;
      17040:data<=16'd10357;
      17041:data<=16'd7762;
      17042:data<=16'd9163;
      17043:data<=16'd9132;
      17044:data<=16'd7735;
      17045:data<=16'd9718;
      17046:data<=16'd10436;
      17047:data<=16'd10214;
      17048:data<=16'd10607;
      17049:data<=16'd9787;
      17050:data<=16'd9771;
      17051:data<=16'd9649;
      17052:data<=16'd8728;
      17053:data<=16'd9658;
      17054:data<=16'd11000;
      17055:data<=16'd11373;
      17056:data<=16'd10981;
      17057:data<=16'd10114;
      17058:data<=16'd10143;
      17059:data<=16'd10064;
      17060:data<=16'd9503;
      17061:data<=16'd9855;
      17062:data<=16'd10625;
      17063:data<=16'd11233;
      17064:data<=16'd11242;
      17065:data<=16'd11148;
      17066:data<=16'd11270;
      17067:data<=16'd10399;
      17068:data<=16'd9773;
      17069:data<=16'd9687;
      17070:data<=16'd9677;
      17071:data<=16'd10941;
      17072:data<=16'd11100;
      17073:data<=16'd10343;
      17074:data<=16'd10760;
      17075:data<=16'd9973;
      17076:data<=16'd9547;
      17077:data<=16'd9858;
      17078:data<=16'd9740;
      17079:data<=16'd12684;
      17080:data<=16'd13623;
      17081:data<=16'd11395;
      17082:data<=16'd12881;
      17083:data<=16'd9059;
      17084:data<=-16'd916;
      17085:data<=-16'd2641;
      17086:data<=-16'd449;
      17087:data<=-16'd823;
      17088:data<=16'd349;
      17089:data<=16'd1283;
      17090:data<=16'd1301;
      17091:data<=16'd1084;
      17092:data<=16'd238;
      17093:data<=16'd948;
      17094:data<=16'd1362;
      17095:data<=16'd1489;
      17096:data<=16'd3159;
      17097:data<=16'd3392;
      17098:data<=16'd2889;
      17099:data<=16'd2769;
      17100:data<=16'd2320;
      17101:data<=16'd3016;
      17102:data<=16'd3004;
      17103:data<=16'd2975;
      17104:data<=16'd4884;
      17105:data<=16'd5118;
      17106:data<=16'd4628;
      17107:data<=16'd5015;
      17108:data<=16'd4408;
      17109:data<=16'd4435;
      17110:data<=16'd4117;
      17111:data<=16'd3062;
      17112:data<=16'd4425;
      17113:data<=16'd5927;
      17114:data<=16'd5915;
      17115:data<=16'd5859;
      17116:data<=16'd5439;
      17117:data<=16'd5074;
      17118:data<=16'd4502;
      17119:data<=16'd3971;
      17120:data<=16'd4543;
      17121:data<=16'd5260;
      17122:data<=16'd5853;
      17123:data<=16'd5494;
      17124:data<=16'd4993;
      17125:data<=16'd5623;
      17126:data<=16'd4223;
      17127:data<=16'd5421;
      17128:data<=16'd13820;
      17129:data<=16'd18848;
      17130:data<=16'd17735;
      17131:data<=16'd17623;
      17132:data<=16'd16363;
      17133:data<=16'd13717;
      17134:data<=16'd13282;
      17135:data<=16'd12690;
      17136:data<=16'd11326;
      17137:data<=16'd11561;
      17138:data<=16'd12703;
      17139:data<=16'd12229;
      17140:data<=16'd10493;
      17141:data<=16'd10146;
      17142:data<=16'd10157;
      17143:data<=16'd9109;
      17144:data<=16'd8587;
      17145:data<=16'd8907;
      17146:data<=16'd9793;
      17147:data<=16'd9994;
      17148:data<=16'd8661;
      17149:data<=16'd7931;
      17150:data<=16'd7500;
      17151:data<=16'd6792;
      17152:data<=16'd6987;
      17153:data<=16'd6792;
      17154:data<=16'd6777;
      17155:data<=16'd7498;
      17156:data<=16'd7083;
      17157:data<=16'd6583;
      17158:data<=16'd5868;
      17159:data<=16'd4899;
      17160:data<=16'd5345;
      17161:data<=16'd4716;
      17162:data<=16'd4084;
      17163:data<=16'd5706;
      17164:data<=16'd5485;
      17165:data<=16'd4467;
      17166:data<=16'd4763;
      17167:data<=16'd4029;
      17168:data<=16'd4035;
      17169:data<=16'd3720;
      17170:data<=16'd2576;
      17171:data<=16'd4050;
      17172:data<=16'd496;
      17173:data<=-16'd9392;
      17174:data<=-16'd12105;
      17175:data<=-16'd9903;
      17176:data<=-16'd11176;
      17177:data<=-16'd10966;
      17178:data<=-16'd9683;
      17179:data<=-16'd11223;
      17180:data<=-16'd11909;
      17181:data<=-16'd11232;
      17182:data<=-16'd10950;
      17183:data<=-16'd10674;
      17184:data<=-16'd10763;
      17185:data<=-16'd9462;
      17186:data<=-16'd7109;
      17187:data<=-16'd7721;
      17188:data<=-16'd9647;
      17189:data<=-16'd9632;
      17190:data<=-16'd9380;
      17191:data<=-16'd9376;
      17192:data<=-16'd8771;
      17193:data<=-16'd8414;
      17194:data<=-16'd8002;
      17195:data<=-16'd7905;
      17196:data<=-16'd9524;
      17197:data<=-16'd10736;
      17198:data<=-16'd10013;
      17199:data<=-16'd9608;
      17200:data<=-16'd9620;
      17201:data<=-16'd8990;
      17202:data<=-16'd8725;
      17203:data<=-16'd8599;
      17204:data<=-16'd8546;
      17205:data<=-16'd9482;
      17206:data<=-16'd10149;
      17207:data<=-16'd9770;
      17208:data<=-16'd9232;
      17209:data<=-16'd9031;
      17210:data<=-16'd9010;
      17211:data<=-16'd8464;
      17212:data<=-16'd8836;
      17213:data<=-16'd10387;
      17214:data<=-16'd10140;
      17215:data<=-16'd9890;
      17216:data<=-16'd8965;
      17217:data<=-16'd1741;
      17218:data<=16'd5222;
      17219:data<=16'd4890;
      17220:data<=16'd3419;
      17221:data<=16'd2887;
      17222:data<=16'd1864;
      17223:data<=16'd1970;
      17224:data<=16'd1436;
      17225:data<=16'd737;
      17226:data<=16'd1021;
      17227:data<=16'd429;
      17228:data<=16'd529;
      17229:data<=16'd447;
      17230:data<=-16'd1579;
      17231:data<=-16'd2320;
      17232:data<=-16'd2100;
      17233:data<=-16'd2002;
      17234:data<=-16'd1381;
      17235:data<=-16'd1924;
      17236:data<=-16'd2053;
      17237:data<=-16'd1882;
      17238:data<=-16'd4595;
      17239:data<=-16'd6789;
      17240:data<=-16'd6567;
      17241:data<=-16'd6669;
      17242:data<=-16'd6441;
      17243:data<=-16'd5779;
      17244:data<=-16'd5812;
      17245:data<=-16'd6012;
      17246:data<=-16'd6443;
      17247:data<=-16'd7150;
      17248:data<=-16'd7526;
      17249:data<=-16'd7087;
      17250:data<=-16'd6419;
      17251:data<=-16'd6112;
      17252:data<=-16'd5485;
      17253:data<=-16'd5310;
      17254:data<=-16'd5974;
      17255:data<=-16'd6501;
      17256:data<=-16'd6751;
      17257:data<=-16'd5846;
      17258:data<=-16'd5680;
      17259:data<=-16'd6522;
      17260:data<=-16'd4508;
      17261:data<=-16'd6663;
      17262:data<=-16'd16551;
      17263:data<=-16'd20926;
      17264:data<=-16'd19077;
      17265:data<=-16'd19364;
      17266:data<=-16'd18421;
      17267:data<=-16'd16675;
      17268:data<=-16'd17026;
      17269:data<=-16'd16104;
      17270:data<=-16'd14992;
      17271:data<=-16'd15432;
      17272:data<=-16'd15670;
      17273:data<=-16'd15218;
      17274:data<=-16'd14116;
      17275:data<=-16'd13242;
      17276:data<=-16'd12402;
      17277:data<=-16'd11239;
      17278:data<=-16'd11045;
      17279:data<=-16'd11053;
      17280:data<=-16'd11203;
      17281:data<=-16'd11476;
      17282:data<=-16'd10345;
      17283:data<=-16'd9532;
      17284:data<=-16'd9226;
      17285:data<=-16'd8202;
      17286:data<=-16'd8046;
      17287:data<=-16'd8134;
      17288:data<=-16'd8294;
      17289:data<=-16'd8956;
      17290:data<=-16'd8388;
      17291:data<=-16'd7386;
      17292:data<=-16'd5962;
      17293:data<=-16'd4478;
      17294:data<=-16'd4758;
      17295:data<=-16'd4096;
      17296:data<=-16'd3554;
      17297:data<=-16'd5215;
      17298:data<=-16'd5078;
      17299:data<=-16'd4684;
      17300:data<=-16'd5080;
      17301:data<=-16'd3926;
      17302:data<=-16'd4167;
      17303:data<=-16'd3932;
      17304:data<=-16'd2776;
      17305:data<=-16'd3706;
      17306:data<=16'd1368;
      17307:data<=16'd10672;
      17308:data<=16'd11837;
      17309:data<=16'd9764;
      17310:data<=16'd10499;
      17311:data<=16'd10134;
      17312:data<=16'd9784;
      17313:data<=16'd10862;
      17314:data<=16'd11559;
      17315:data<=16'd11430;
      17316:data<=16'd10903;
      17317:data<=16'd10800;
      17318:data<=16'd10654;
      17319:data<=16'd10243;
      17320:data<=16'd9928;
      17321:data<=16'd9897;
      17322:data<=16'd11279;
      17323:data<=16'd12148;
      17324:data<=16'd11116;
      17325:data<=16'd10501;
      17326:data<=16'd9881;
      17327:data<=16'd9288;
      17328:data<=16'd9514;
      17329:data<=16'd9421;
      17330:data<=16'd10278;
      17331:data<=16'd10998;
      17332:data<=16'd10058;
      17333:data<=16'd10014;
      17334:data<=16'd9781;
      17335:data<=16'd8934;
      17336:data<=16'd8948;
      17337:data<=16'd8369;
      17338:data<=16'd9048;
      17339:data<=16'd10608;
      17340:data<=16'd10058;
      17341:data<=16'd9703;
      17342:data<=16'd9392;
      17343:data<=16'd8931;
      17344:data<=16'd9085;
      17345:data<=16'd7083;
      17346:data<=16'd6614;
      17347:data<=16'd8414;
      17348:data<=16'd7768;
      17349:data<=16'd8426;
      17350:data<=16'd6266;
      17351:data<=-16'd3131;
      17352:data<=-16'd7092;
      17353:data<=-16'd5210;
      17354:data<=-16'd5709;
      17355:data<=-16'd4526;
      17356:data<=-16'd3019;
      17357:data<=-16'd3677;
      17358:data<=-16'd2881;
      17359:data<=-16'd2755;
      17360:data<=-16'd2977;
      17361:data<=-16'd1902;
      17362:data<=-16'd2129;
      17363:data<=-16'd1571;
      17364:data<=16'd53;
      17365:data<=16'd170;
      17366:data<=16'd575;
      17367:data<=16'd1010;
      17368:data<=16'd764;
      17369:data<=16'd958;
      17370:data<=16'd805;
      17371:data<=16'd1535;
      17372:data<=16'd3532;
      17373:data<=16'd3964;
      17374:data<=16'd3083;
      17375:data<=16'd2617;
      17376:data<=16'd2849;
      17377:data<=16'd3145;
      17378:data<=16'd2784;
      17379:data<=16'd3072;
      17380:data<=16'd4296;
      17381:data<=16'd4789;
      17382:data<=16'd4690;
      17383:data<=16'd4378;
      17384:data<=16'd3751;
      17385:data<=16'd3516;
      17386:data<=16'd3758;
      17387:data<=16'd3720;
      17388:data<=16'd3629;
      17389:data<=16'd4836;
      17390:data<=16'd5580;
      17391:data<=16'd4087;
      17392:data<=16'd4388;
      17393:data<=16'd5218;
      17394:data<=16'd2675;
      17395:data<=16'd5823;
      17396:data<=16'd16128;
      17397:data<=16'd19754;
      17398:data<=16'd18107;
      17399:data<=16'd19511;
      17400:data<=16'd19237;
      17401:data<=16'd17192;
      17402:data<=16'd17291;
      17403:data<=16'd16230;
      17404:data<=16'd14942;
      17405:data<=16'd15919;
      17406:data<=16'd15952;
      17407:data<=16'd14933;
      17408:data<=16'd14325;
      17409:data<=16'd13271;
      17410:data<=16'd12690;
      17411:data<=16'd12563;
      17412:data<=16'd11837;
      17413:data<=16'd11815;
      17414:data<=16'd12267;
      17415:data<=16'd11673;
      17416:data<=16'd10749;
      17417:data<=16'd9958;
      17418:data<=16'd9157;
      17419:data<=16'd8622;
      17420:data<=16'd8084;
      17421:data<=16'd8349;
      17422:data<=16'd9359;
      17423:data<=16'd8848;
      17424:data<=16'd7788;
      17425:data<=16'd7952;
      17426:data<=16'd7736;
      17427:data<=16'd7194;
      17428:data<=16'd7068;
      17429:data<=16'd6739;
      17430:data<=16'd7048;
      17431:data<=16'd7377;
      17432:data<=16'd6771;
      17433:data<=16'd6626;
      17434:data<=16'd6631;
      17435:data<=16'd6260;
      17436:data<=16'd5567;
      17437:data<=16'd4639;
      17438:data<=16'd5341;
      17439:data<=16'd3844;
      17440:data<=-16'd3838;
      17441:data<=-16'd9570;
      17442:data<=-16'd9157;
      17443:data<=-16'd8698;
      17444:data<=-16'd9010;
      17445:data<=-16'd8783;
      17446:data<=-16'd9232;
      17447:data<=-16'd9605;
      17448:data<=-16'd9855;
      17449:data<=-16'd10094;
      17450:data<=-16'd9899;
      17451:data<=-16'd10194;
      17452:data<=-16'd10693;
      17453:data<=-16'd10683;
      17454:data<=-16'd10493;
      17455:data<=-16'd11012;
      17456:data<=-16'd12386;
      17457:data<=-16'd12384;
      17458:data<=-16'd11268;
      17459:data<=-16'd11326;
      17460:data<=-16'd11362;
      17461:data<=-16'd10686;
      17462:data<=-16'd9988;
      17463:data<=-16'd9785;
      17464:data<=-16'd10978;
      17465:data<=-16'd11644;
      17466:data<=-16'd11028;
      17467:data<=-16'd10671;
      17468:data<=-16'd10026;
      17469:data<=-16'd10147;
      17470:data<=-16'd10381;
      17471:data<=-16'd9007;
      17472:data<=-16'd9589;
      17473:data<=-16'd11147;
      17474:data<=-16'd10584;
      17475:data<=-16'd10246;
      17476:data<=-16'd9579;
      17477:data<=-16'd9107;
      17478:data<=-16'd9505;
      17479:data<=-16'd8035;
      17480:data<=-16'd8614;
      17481:data<=-16'd10701;
      17482:data<=-16'd9964;
      17483:data<=-16'd10968;
      17484:data<=-16'd8194;
      17485:data<=16'd1862;
      17486:data<=16'd4940;
      17487:data<=16'd2726;
      17488:data<=16'd3933;
      17489:data<=16'd2384;
      17490:data<=16'd332;
      17491:data<=16'd1503;
      17492:data<=16'd946;
      17493:data<=16'd644;
      17494:data<=16'd1101;
      17495:data<=16'd406;
      17496:data<=16'd772;
      17497:data<=-16'd62;
      17498:data<=-16'd1902;
      17499:data<=-16'd1642;
      17500:data<=-16'd1480;
      17501:data<=-16'd1310;
      17502:data<=-16'd1134;
      17503:data<=-16'd2237;
      17504:data<=-16'd1418;
      17505:data<=-16'd79;
      17506:data<=-16'd1459;
      17507:data<=-16'd2235;
      17508:data<=-16'd1679;
      17509:data<=-16'd1917;
      17510:data<=-16'd2123;
      17511:data<=-16'd1756;
      17512:data<=-16'd1340;
      17513:data<=-16'd1739;
      17514:data<=-16'd2936;
      17515:data<=-16'd3286;
      17516:data<=-16'd3055;
      17517:data<=-16'd3309;
      17518:data<=-16'd3250;
      17519:data<=-16'd2996;
      17520:data<=-16'd3110;
      17521:data<=-16'd2742;
      17522:data<=-16'd2760;
      17523:data<=-16'd4214;
      17524:data<=-16'd4370;
      17525:data<=-16'd3071;
      17526:data<=-16'd3620;
      17527:data<=-16'd3735;
      17528:data<=-16'd3018;
      17529:data<=-16'd8031;
      17530:data<=-16'd15637;
      17531:data<=-16'd16779;
      17532:data<=-16'd14502;
      17533:data<=-16'd14064;
      17534:data<=-16'd13248;
      17535:data<=-16'd11811;
      17536:data<=-16'd11320;
      17537:data<=-16'd10487;
      17538:data<=-16'd9949;
      17539:data<=-16'd11097;
      17540:data<=-16'd11385;
      17541:data<=-16'd10081;
      17542:data<=-16'd9787;
      17543:data<=-16'd9747;
      17544:data<=-16'd8990;
      17545:data<=-16'd8865;
      17546:data<=-16'd8563;
      17547:data<=-16'd8244;
      17548:data<=-16'd8827;
      17549:data<=-16'd8526;
      17550:data<=-16'd7803;
      17551:data<=-16'd7733;
      17552:data<=-16'd7062;
      17553:data<=-16'd6219;
      17554:data<=-16'd5645;
      17555:data<=-16'd5645;
      17556:data<=-16'd6608;
      17557:data<=-16'd6551;
      17558:data<=-16'd5836;
      17559:data<=-16'd5753;
      17560:data<=-16'd5300;
      17561:data<=-16'd5553;
      17562:data<=-16'd5900;
      17563:data<=-16'd4828;
      17564:data<=-16'd4817;
      17565:data<=-16'd5720;
      17566:data<=-16'd5786;
      17567:data<=-16'd5325;
      17568:data<=-16'd4482;
      17569:data<=-16'd4663;
      17570:data<=-16'd4528;
      17571:data<=-16'd3383;
      17572:data<=-16'd4332;
      17573:data<=-16'd1977;
      17574:data<=16'd5981;
      17575:data<=16'd9107;
      17576:data<=16'd7447;
      17577:data<=16'd7794;
      17578:data<=16'd8053;
      17579:data<=16'd7609;
      17580:data<=16'd7726;
      17581:data<=16'd7923;
      17582:data<=16'd8815;
      17583:data<=16'd9034;
      17584:data<=16'd8369;
      17585:data<=16'd8119;
      17586:data<=16'd8066;
      17587:data<=16'd8599;
      17588:data<=16'd8328;
      17589:data<=16'd7749;
      17590:data<=16'd9467;
      17591:data<=16'd10322;
      17592:data<=16'd9279;
      17593:data<=16'd9113;
      17594:data<=16'd8789;
      17595:data<=16'd8258;
      17596:data<=16'd7858;
      17597:data<=16'd7691;
      17598:data<=16'd9025;
      17599:data<=16'd9024;
      17600:data<=16'd7799;
      17601:data<=16'd8467;
      17602:data<=16'd8596;
      17603:data<=16'd8175;
      17604:data<=16'd8222;
      17605:data<=16'd7488;
      17606:data<=16'd8437;
      17607:data<=16'd9799;
      17608:data<=16'd9318;
      17609:data<=16'd9292;
      17610:data<=16'd8737;
      17611:data<=16'd8549;
      17612:data<=16'd9277;
      17613:data<=16'd8002;
      17614:data<=16'd8614;
      17615:data<=16'd10383;
      17616:data<=16'd9359;
      17617:data<=16'd9896;
      17618:data<=16'd7001;
      17619:data<=-16'd1480;
      17620:data<=-16'd3099;
      17621:data<=-16'd889;
      17622:data<=-16'd1970;
      17623:data<=-16'd387;
      17624:data<=16'd1368;
      17625:data<=16'd411;
      17626:data<=16'd977;
      17627:data<=16'd1075;
      17628:data<=16'd658;
      17629:data<=16'd1375;
      17630:data<=16'd1093;
      17631:data<=16'd1368;
      17632:data<=16'd2370;
      17633:data<=16'd2238;
      17634:data<=16'd2252;
      17635:data<=16'd2223;
      17636:data<=16'd2105;
      17637:data<=16'd2261;
      17638:data<=16'd2003;
      17639:data<=16'd3005;
      17640:data<=16'd4798;
      17641:data<=16'd5245;
      17642:data<=16'd5338;
      17643:data<=16'd5236;
      17644:data<=16'd5127;
      17645:data<=16'd5418;
      17646:data<=16'd4601;
      17647:data<=16'd4419;
      17648:data<=16'd6390;
      17649:data<=16'd7015;
      17650:data<=16'd5903;
      17651:data<=16'd5800;
      17652:data<=16'd5808;
      17653:data<=16'd5084;
      17654:data<=16'd4683;
      17655:data<=16'd4168;
      17656:data<=16'd4384;
      17657:data<=16'd5885;
      17658:data<=16'd5768;
      17659:data<=16'd5159;
      17660:data<=16'd5818;
      17661:data<=16'd4616;
      17662:data<=16'd5318;
      17663:data<=16'd11552;
      17664:data<=16'd15590;
      17665:data<=16'd15429;
      17666:data<=16'd15474;
      17667:data<=16'd15023;
      17668:data<=16'd14411;
      17669:data<=16'd13735;
      17670:data<=16'd12075;
      17671:data<=16'd11468;
      17672:data<=16'd11488;
      17673:data<=16'd11605;
      17674:data<=16'd12057;
      17675:data<=16'd11370;
      17676:data<=16'd11188;
      17677:data<=16'd11260;
      17678:data<=16'd10014;
      17679:data<=16'd9650;
      17680:data<=16'd8916;
      17681:data<=16'd8041;
      17682:data<=16'd9467;
      17683:data<=16'd9468;
      17684:data<=16'd8047;
      17685:data<=16'd7897;
      17686:data<=16'd7219;
      17687:data<=16'd6590;
      17688:data<=16'd6188;
      17689:data<=16'd6056;
      17690:data<=16'd7192;
      17691:data<=16'd6501;
      17692:data<=16'd5234;
      17693:data<=16'd5648;
      17694:data<=16'd4679;
      17695:data<=16'd3923;
      17696:data<=16'd4058;
      17697:data<=16'd3462;
      17698:data<=16'd4469;
      17699:data<=16'd5168;
      17700:data<=16'd4293;
      17701:data<=16'd3883;
      17702:data<=16'd3175;
      17703:data<=16'd3580;
      17704:data<=16'd3356;
      17705:data<=16'd1668;
      17706:data<=16'd3231;
      17707:data<=16'd957;
      17708:data<=-16'd7715;
      17709:data<=-16'd10058;
      17710:data<=-16'd8108;
      17711:data<=-16'd9257;
      17712:data<=-16'd9209;
      17713:data<=-16'd8334;
      17714:data<=-16'd8919;
      17715:data<=-16'd9465;
      17716:data<=-16'd9843;
      17717:data<=-16'd9589;
      17718:data<=-16'd9529;
      17719:data<=-16'd9867;
      17720:data<=-16'd9897;
      17721:data<=-16'd10146;
      17722:data<=-16'd9244;
      17723:data<=-16'd9097;
      17724:data<=-16'd11186;
      17725:data<=-16'd11236;
      17726:data<=-16'd10464;
      17727:data<=-16'd10898;
      17728:data<=-16'd10407;
      17729:data<=-16'd10278;
      17730:data<=-16'd9988;
      17731:data<=-16'd9567;
      17732:data<=-16'd11129;
      17733:data<=-16'd11309;
      17734:data<=-16'd10298;
      17735:data<=-16'd10581;
      17736:data<=-16'd9987;
      17737:data<=-16'd9721;
      17738:data<=-16'd10187;
      17739:data<=-16'd9958;
      17740:data<=-16'd10736;
      17741:data<=-16'd11089;
      17742:data<=-16'd10525;
      17743:data<=-16'd10443;
      17744:data<=-16'd9767;
      17745:data<=-16'd10066;
      17746:data<=-16'd10334;
      17747:data<=-16'd8868;
      17748:data<=-16'd9468;
      17749:data<=-16'd10889;
      17750:data<=-16'd11077;
      17751:data<=-16'd10387;
      17752:data<=-16'd5122;
      17753:data<=16'd411;
      17754:data<=16'd355;
      17755:data<=16'd114;
      17756:data<=16'd306;
      17757:data<=-16'd1789;
      17758:data<=-16'd2544;
      17759:data<=-16'd1918;
      17760:data<=-16'd2217;
      17761:data<=-16'd2746;
      17762:data<=-16'd2728;
      17763:data<=-16'd2205;
      17764:data<=-16'd2457;
      17765:data<=-16'd3171;
      17766:data<=-16'd3504;
      17767:data<=-16'd4482;
      17768:data<=-16'd4723;
      17769:data<=-16'd3914;
      17770:data<=-16'd4152;
      17771:data<=-16'd4049;
      17772:data<=-16'd3397;
      17773:data<=-16'd4454;
      17774:data<=-16'd5990;
      17775:data<=-16'd6173;
      17776:data<=-16'd5838;
      17777:data<=-16'd5849;
      17778:data<=-16'd5718;
      17779:data<=-16'd5470;
      17780:data<=-16'd5539;
      17781:data<=-16'd5530;
      17782:data<=-16'd6109;
      17783:data<=-16'd6881;
      17784:data<=-16'd6341;
      17785:data<=-16'd6088;
      17786:data<=-16'd6122;
      17787:data<=-16'd5603;
      17788:data<=-16'd5761;
      17789:data<=-16'd4931;
      17790:data<=-16'd4817;
      17791:data<=-16'd7165;
      17792:data<=-16'd6608;
      17793:data<=-16'd5601;
      17794:data<=-16'd6733;
      17795:data<=-16'd4857;
      17796:data<=-16'd6564;
      17797:data<=-16'd14254;
      17798:data<=-16'd16874;
      17799:data<=-16'd16233;
      17800:data<=-16'd16675;
      17801:data<=-16'd15250;
      17802:data<=-16'd14358;
      17803:data<=-16'd13612;
      17804:data<=-16'd12003;
      17805:data<=-16'd12349;
      17806:data<=-16'd12477;
      17807:data<=-16'd12410;
      17808:data<=-16'd13215;
      17809:data<=-16'd12628;
      17810:data<=-16'd12251;
      17811:data<=-16'd11585;
      17812:data<=-16'd9824;
      17813:data<=-16'd9670;
      17814:data<=-16'd9204;
      17815:data<=-16'd8751;
      17816:data<=-16'd10044;
      17817:data<=-16'd9755;
      17818:data<=-16'd8784;
      17819:data<=-16'd8401;
      17820:data<=-16'd7471;
      17821:data<=-16'd7321;
      17822:data<=-16'd6601;
      17823:data<=-16'd6181;
      17824:data<=-16'd7783;
      17825:data<=-16'd7571;
      17826:data<=-16'd6620;
      17827:data<=-16'd6862;
      17828:data<=-16'd6179;
      17829:data<=-16'd5859;
      17830:data<=-16'd5194;
      17831:data<=-16'd4267;
      17832:data<=-16'd5435;
      17833:data<=-16'd5755;
      17834:data<=-16'd5533;
      17835:data<=-16'd5850;
      17836:data<=-16'd4637;
      17837:data<=-16'd4620;
      17838:data<=-16'd4444;
      17839:data<=-16'd3109;
      17840:data<=-16'd4197;
      17841:data<=-16'd516;
      17842:data<=16'd8006;
      17843:data<=16'd9368;
      17844:data<=16'd7495;
      17845:data<=16'd8699;
      17846:data<=16'd8346;
      17847:data<=16'd7242;
      17848:data<=16'd8012;
      17849:data<=16'd9168;
      17850:data<=16'd9539;
      17851:data<=16'd9056;
      17852:data<=16'd9036;
      17853:data<=16'd9162;
      17854:data<=16'd9022;
      17855:data<=16'd9006;
      17856:data<=16'd8223;
      17857:data<=16'd8708;
      17858:data<=16'd10329;
      17859:data<=16'd9925;
      17860:data<=16'd9682;
      17861:data<=16'd10105;
      17862:data<=16'd9511;
      17863:data<=16'd9353;
      17864:data<=16'd8945;
      17865:data<=16'd9045;
      17866:data<=16'd10696;
      17867:data<=16'd11039;
      17868:data<=16'd10686;
      17869:data<=16'd10610;
      17870:data<=16'd10219;
      17871:data<=16'd10379;
      17872:data<=16'd9794;
      17873:data<=16'd9737;
      17874:data<=16'd11264;
      17875:data<=16'd11106;
      17876:data<=16'd10989;
      17877:data<=16'd11500;
      17878:data<=16'd10322;
      17879:data<=16'd10155;
      17880:data<=16'd10399;
      17881:data<=16'd9831;
      17882:data<=16'd10292;
      17883:data<=16'd10484;
      17884:data<=16'd11314;
      17885:data<=16'd10081;
      17886:data<=16'd2957;
      17887:data<=-16'd1083;
      17888:data<=16'd143;
      17889:data<=-16'd723;
      17890:data<=-16'd503;
      17891:data<=16'd1698;
      17892:data<=16'd1729;
      17893:data<=16'd1912;
      17894:data<=16'd2601;
      17895:data<=16'd2648;
      17896:data<=16'd2952;
      17897:data<=16'd2734;
      17898:data<=16'd2698;
      17899:data<=16'd3527;
      17900:data<=16'd4416;
      17901:data<=16'd4937;
      17902:data<=16'd4275;
      17903:data<=16'd3968;
      17904:data<=16'd4833;
      17905:data<=16'd4576;
      17906:data<=16'd4047;
      17907:data<=16'd5136;
      17908:data<=16'd6563;
      17909:data<=16'd6704;
      17910:data<=16'd6128;
      17911:data<=16'd6149;
      17912:data<=16'd5735;
      17913:data<=16'd5156;
      17914:data<=16'd5885;
      17915:data<=16'd6131;
      17916:data<=16'd6234;
      17917:data<=16'd6874;
      17918:data<=16'd6320;
      17919:data<=16'd6328;
      17920:data<=16'd6473;
      17921:data<=16'd5492;
      17922:data<=16'd5785;
      17923:data<=16'd5662;
      17924:data<=16'd5911;
      17925:data<=16'd7840;
      17926:data<=16'd6616;
      17927:data<=16'd6029;
      17928:data<=16'd7451;
      17929:data<=16'd4916;
      17930:data<=16'd6913;
      17931:data<=16'd14897;
      17932:data<=16'd16854;
      17933:data<=16'd16607;
      17934:data<=16'd17728;
      17935:data<=16'd15697;
      17936:data<=16'd14492;
      17937:data<=16'd14540;
      17938:data<=16'd13330;
      17939:data<=16'd12927;
      17940:data<=16'd12574;
      17941:data<=16'd12969;
      17942:data<=16'd13990;
      17943:data<=16'd12971;
      17944:data<=16'd11894;
      17945:data<=16'd11135;
      17946:data<=16'd10278;
      17947:data<=16'd10425;
      17948:data<=16'd9526;
      17949:data<=16'd9028;
      17950:data<=16'd10270;
      17951:data<=16'd10328;
      17952:data<=16'd10032;
      17953:data<=16'd9473;
      17954:data<=16'd8185;
      17955:data<=16'd8034;
      17956:data<=16'd7605;
      17957:data<=16'd7685;
      17958:data<=16'd9033;
      17959:data<=16'd8526;
      17960:data<=16'd7984;
      17961:data<=16'd8091;
      17962:data<=16'd6822;
      17963:data<=16'd6445;
      17964:data<=16'd6391;
      17965:data<=16'd5785;
      17966:data<=16'd6470;
      17967:data<=16'd6695;
      17968:data<=16'd5965;
      17969:data<=16'd5609;
      17970:data<=16'd5612;
      17971:data<=16'd5661;
      17972:data<=16'd4449;
      17973:data<=16'd3861;
      17974:data<=16'd3240;
      17975:data<=-16'd2370;
      17976:data<=-16'd7837;
      17977:data<=-16'd7970;
      17978:data<=-16'd7639;
      17979:data<=-16'd7858;
      17980:data<=-16'd7336;
      17981:data<=-16'd7133;
      17982:data<=-16'd7385;
      17983:data<=-16'd8878;
      17984:data<=-16'd9812;
      17985:data<=-16'd9033;
      17986:data<=-16'd8799;
      17987:data<=-16'd8743;
      17988:data<=-16'd8812;
      17989:data<=-16'd8736;
      17990:data<=-16'd7973;
      17991:data<=-16'd9124;
      17992:data<=-16'd10334;
      17993:data<=-16'd9790;
      17994:data<=-16'd9950;
      17995:data<=-16'd9329;
      17996:data<=-16'd8583;
      17997:data<=-16'd9022;
      17998:data<=-16'd8310;
      17999:data<=-16'd8881;
      18000:data<=-16'd10343;
      18001:data<=-16'd9934;
      18002:data<=-16'd10329;
      18003:data<=-16'd10351;
      18004:data<=-16'd9787;
      18005:data<=-16'd10360;
      18006:data<=-16'd9036;
      18007:data<=-16'd8748;
      18008:data<=-16'd11018;
      18009:data<=-16'd11016;
      18010:data<=-16'd10686;
      18011:data<=-16'd10775;
      18012:data<=-16'd10016;
      18013:data<=-16'd10058;
      18014:data<=-16'd9213;
      18015:data<=-16'd9210;
      18016:data<=-16'd10502;
      18017:data<=-16'd10096;
      18018:data<=-16'd11069;
      18019:data<=-16'd8557;
      18020:data<=16'd56;
      18021:data<=16'd2344;
      18022:data<=16'd437;
      18023:data<=16'd1780;
      18024:data<=16'd334;
      18025:data<=-16'd1912;
      18026:data<=-16'd1491;
      18027:data<=-16'd1882;
      18028:data<=-16'd1362;
      18029:data<=-16'd643;
      18030:data<=-16'd1360;
      18031:data<=-16'd1102;
      18032:data<=-16'd1353;
      18033:data<=-16'd2649;
      18034:data<=-16'd3551;
      18035:data<=-16'd4241;
      18036:data<=-16'd4079;
      18037:data<=-16'd3912;
      18038:data<=-16'd3908;
      18039:data<=-16'd3386;
      18040:data<=-16'd3671;
      18041:data<=-16'd4229;
      18042:data<=-16'd4821;
      18043:data<=-16'd5545;
      18044:data<=-16'd5154;
      18045:data<=-16'd5143;
      18046:data<=-16'd5521;
      18047:data<=-16'd4757;
      18048:data<=-16'd4081;
      18049:data<=-16'd3956;
      18050:data<=-16'd5033;
      18051:data<=-16'd6203;
      18052:data<=-16'd5166;
      18053:data<=-16'd4502;
      18054:data<=-16'd4698;
      18055:data<=-16'd4266;
      18056:data<=-16'd4284;
      18057:data<=-16'd3832;
      18058:data<=-16'd4570;
      18059:data<=-16'd6622;
      18060:data<=-16'd5738;
      18061:data<=-16'd4995;
      18062:data<=-16'd5206;
      18063:data<=-16'd4416;
      18064:data<=-16'd8930;
      18065:data<=-16'd15669;
      18066:data<=-16'd16628;
      18067:data<=-16'd16331;
      18068:data<=-16'd16656;
      18069:data<=-16'd15594;
      18070:data<=-16'd14839;
      18071:data<=-16'd13961;
      18072:data<=-16'd13453;
      18073:data<=-16'd13136;
      18074:data<=-16'd11944;
      18075:data<=-16'd12518;
      18076:data<=-16'd13456;
      18077:data<=-16'd12516;
      18078:data<=-16'd11779;
      18079:data<=-16'd10916;
      18080:data<=-16'd10094;
      18081:data<=-16'd9903;
      18082:data<=-16'd9283;
      18083:data<=-16'd9787;
      18084:data<=-16'd10869;
      18085:data<=-16'd10525;
      18086:data<=-16'd9714;
      18087:data<=-16'd8695;
      18088:data<=-16'd8210;
      18089:data<=-16'd8244;
      18090:data<=-16'd7579;
      18091:data<=-16'd7844;
      18092:data<=-16'd8657;
      18093:data<=-16'd8583;
      18094:data<=-16'd8549;
      18095:data<=-16'd7873;
      18096:data<=-16'd7090;
      18097:data<=-16'd6918;
      18098:data<=-16'd6323;
      18099:data<=-16'd6548;
      18100:data<=-16'd6943;
      18101:data<=-16'd6548;
      18102:data<=-16'd6570;
      18103:data<=-16'd5823;
      18104:data<=-16'd5366;
      18105:data<=-16'd5462;
      18106:data<=-16'd4270;
      18107:data<=-16'd4726;
      18108:data<=-16'd2933;
      18109:data<=16'd4679;
      18110:data<=16'd7843;
      18111:data<=16'd6355;
      18112:data<=16'd7812;
      18113:data<=16'd8358;
      18114:data<=16'd7307;
      18115:data<=16'd7185;
      18116:data<=16'd6749;
      18117:data<=16'd7840;
      18118:data<=16'd9074;
      18119:data<=16'd8440;
      18120:data<=16'd8237;
      18121:data<=16'd8078;
      18122:data<=16'd8204;
      18123:data<=16'd8225;
      18124:data<=16'd7159;
      18125:data<=16'd8285;
      18126:data<=16'd9734;
      18127:data<=16'd8974;
      18128:data<=16'd9297;
      18129:data<=16'd9556;
      18130:data<=16'd8925;
      18131:data<=16'd8853;
      18132:data<=16'd8364;
      18133:data<=16'd9209;
      18134:data<=16'd10554;
      18135:data<=16'd10257;
      18136:data<=16'd10360;
      18137:data<=16'd9693;
      18138:data<=16'd8824;
      18139:data<=16'd9585;
      18140:data<=16'd9256;
      18141:data<=16'd9462;
      18142:data<=16'd10593;
      18143:data<=16'd10138;
      18144:data<=16'd10386;
      18145:data<=16'd9902;
      18146:data<=16'd8652;
      18147:data<=16'd9855;
      18148:data<=16'd9885;
      18149:data<=16'd9301;
      18150:data<=16'd10155;
      18151:data<=16'd10008;
      18152:data<=16'd10815;
      18153:data<=16'd8263;
      18154:data<=16'd220;
      18155:data<=-16'd2226;
      18156:data<=-16'd667;
      18157:data<=-16'd1767;
      18158:data<=-16'd429;
      18159:data<=16'd2020;
      18160:data<=16'd2208;
      18161:data<=16'd2312;
      18162:data<=16'd1815;
      18163:data<=16'd1971;
      18164:data<=16'd2455;
      18165:data<=16'd928;
      18166:data<=16'd734;
      18167:data<=16'd2505;
      18168:data<=16'd3544;
      18169:data<=16'd4029;
      18170:data<=16'd3647;
      18171:data<=16'd2740;
      18172:data<=16'd2369;
      18173:data<=16'd2384;
      18174:data<=16'd2845;
      18175:data<=16'd3338;
      18176:data<=16'd4023;
      18177:data<=16'd4804;
      18178:data<=16'd4360;
      18179:data<=16'd3541;
      18180:data<=16'd3720;
      18181:data<=16'd4161;
      18182:data<=16'd3983;
      18183:data<=16'd4118;
      18184:data<=16'd5190;
      18185:data<=16'd5081;
      18186:data<=16'd4270;
      18187:data<=16'd4652;
      18188:data<=16'd4193;
      18189:data<=16'd3521;
      18190:data<=16'd3847;
      18191:data<=16'd3488;
      18192:data<=16'd3915;
      18193:data<=16'd4446;
      18194:data<=16'd4014;
      18195:data<=16'd4496;
      18196:data<=16'd3357;
      18197:data<=16'd3991;
      18198:data<=16'd10762;
      18199:data<=16'd14495;
      18200:data<=16'd13944;
      18201:data<=16'd15314;
      18202:data<=16'd15015;
      18203:data<=16'd13493;
      18204:data<=16'd13244;
      18205:data<=16'd12058;
      18206:data<=16'd11676;
      18207:data<=16'd11327;
      18208:data<=16'd10155;
      18209:data<=16'd11267;
      18210:data<=16'd12405;
      18211:data<=16'd11990;
      18212:data<=16'd11195;
      18213:data<=16'd9788;
      18214:data<=16'd9221;
      18215:data<=16'd8617;
      18216:data<=16'd8193;
      18217:data<=16'd9894;
      18218:data<=16'd10125;
      18219:data<=16'd8860;
      18220:data<=16'd8516;
      18221:data<=16'd7570;
      18222:data<=16'd7486;
      18223:data<=16'd7608;
      18224:data<=16'd6708;
      18225:data<=16'd7815;
      18226:data<=16'd8337;
      18227:data<=16'd7030;
      18228:data<=16'd7033;
      18229:data<=16'd6514;
      18230:data<=16'd5749;
      18231:data<=16'd5782;
      18232:data<=16'd5009;
      18233:data<=16'd5257;
      18234:data<=16'd6264;
      18235:data<=16'd6595;
      18236:data<=16'd6716;
      18237:data<=16'd5841;
      18238:data<=16'd5553;
      18239:data<=16'd5335;
      18240:data<=16'd4452;
      18241:data<=16'd5471;
      18242:data<=16'd2414;
      18243:data<=-16'd5820;
      18244:data<=-16'd8663;
      18245:data<=-16'd7708;
      18246:data<=-16'd8436;
      18247:data<=-16'd8301;
      18248:data<=-16'd7777;
      18249:data<=-16'd7233;
      18250:data<=-16'd7380;
      18251:data<=-16'd9310;
      18252:data<=-16'd9318;
      18253:data<=-16'd8416;
      18254:data<=-16'd8843;
      18255:data<=-16'd8692;
      18256:data<=-16'd9027;
      18257:data<=-16'd8901;
      18258:data<=-16'd7934;
      18259:data<=-16'd9025;
      18260:data<=-16'd9809;
      18261:data<=-16'd9665;
      18262:data<=-16'd9935;
      18263:data<=-16'd9135;
      18264:data<=-16'd9726;
      18265:data<=-16'd10875;
      18266:data<=-16'd9244;
      18267:data<=-16'd8590;
      18268:data<=-16'd9544;
      18269:data<=-16'd9765;
      18270:data<=-16'd10266;
      18271:data<=-16'd10372;
      18272:data<=-16'd10078;
      18273:data<=-16'd9683;
      18274:data<=-16'd8680;
      18275:data<=-16'd8980;
      18276:data<=-16'd9999;
      18277:data<=-16'd10119;
      18278:data<=-16'd9900;
      18279:data<=-16'd8997;
      18280:data<=-16'd8569;
      18281:data<=-16'd9139;
      18282:data<=-16'd9268;
      18283:data<=-16'd9256;
      18284:data<=-16'd9151;
      18285:data<=-16'd10014;
      18286:data<=-16'd10190;
      18287:data<=-16'd4599;
      18288:data<=16'd1650;
      18289:data<=16'd2106;
      18290:data<=16'd1495;
      18291:data<=16'd1633;
      18292:data<=16'd388;
      18293:data<=-16'd587;
      18294:data<=-16'd852;
      18295:data<=-16'd813;
      18296:data<=-16'd459;
      18297:data<=-16'd285;
      18298:data<=-16'd112;
      18299:data<=-16'd403;
      18300:data<=-16'd1074;
      18301:data<=-16'd1738;
      18302:data<=-16'd2519;
      18303:data<=-16'd2544;
      18304:data<=-16'd2566;
      18305:data<=-16'd2928;
      18306:data<=-16'd2312;
      18307:data<=-16'd2005;
      18308:data<=-16'd2390;
      18309:data<=-16'd2864;
      18310:data<=-16'd3973;
      18311:data<=-16'd4044;
      18312:data<=-16'd3298;
      18313:data<=-16'd3466;
      18314:data<=-16'd3398;
      18315:data<=-16'd3022;
      18316:data<=-16'd2717;
      18317:data<=-16'd3125;
      18318:data<=-16'd4710;
      18319:data<=-16'd4780;
      18320:data<=-16'd4112;
      18321:data<=-16'd4540;
      18322:data<=-16'd4124;
      18323:data<=-16'd3802;
      18324:data<=-16'd3653;
      18325:data<=-16'd3400;
      18326:data<=-16'd4678;
      18327:data<=-16'd4323;
      18328:data<=-16'd3654;
      18329:data<=-16'd4689;
      18330:data<=-16'd2722;
      18331:data<=-16'd4369;
      18332:data<=-16'd12469;
      18333:data<=-16'd14815;
      18334:data<=-16'd13667;
      18335:data<=-16'd14951;
      18336:data<=-16'd14051;
      18337:data<=-16'd13054;
      18338:data<=-16'd12598;
      18339:data<=-16'd11118;
      18340:data<=-16'd11386;
      18341:data<=-16'd10495;
      18342:data<=-16'd9502;
      18343:data<=-16'd11577;
      18344:data<=-16'd11521;
      18345:data<=-16'd9973;
      18346:data<=-16'd9767;
      18347:data<=-16'd9303;
      18348:data<=-16'd9445;
      18349:data<=-16'd8678;
      18350:data<=-16'd8073;
      18351:data<=-16'd10184;
      18352:data<=-16'd10326;
      18353:data<=-16'd9095;
      18354:data<=-16'd9036;
      18355:data<=-16'd7559;
      18356:data<=-16'd7235;
      18357:data<=-16'd7985;
      18358:data<=-16'd6708;
      18359:data<=-16'd6801;
      18360:data<=-16'd8005;
      18361:data<=-16'd7221;
      18362:data<=-16'd6150;
      18363:data<=-16'd6423;
      18364:data<=-16'd6936;
      18365:data<=-16'd5615;
      18366:data<=-16'd4504;
      18367:data<=-16'd5598;
      18368:data<=-16'd5844;
      18369:data<=-16'd5981;
      18370:data<=-16'd6246;
      18371:data<=-16'd4484;
      18372:data<=-16'd4091;
      18373:data<=-16'd4196;
      18374:data<=-16'd3738;
      18375:data<=-16'd5406;
      18376:data<=-16'd1541;
      18377:data<=16'd7383;
      18378:data<=16'd8924;
      18379:data<=16'd7228;
      18380:data<=16'd8740;
      18381:data<=16'd8625;
      18382:data<=16'd7424;
      18383:data<=16'd7254;
      18384:data<=16'd7357;
      18385:data<=16'd7815;
      18386:data<=16'd7812;
      18387:data<=16'd8422;
      18388:data<=16'd9317;
      18389:data<=16'd8890;
      18390:data<=16'd8724;
      18391:data<=16'd8093;
      18392:data<=16'd7535;
      18393:data<=16'd9210;
      18394:data<=16'd9903;
      18395:data<=16'd9696;
      18396:data<=16'd10705;
      18397:data<=16'd10329;
      18398:data<=16'd9577;
      18399:data<=16'd9796;
      18400:data<=16'd9200;
      18401:data<=16'd9479;
      18402:data<=16'd10919;
      18403:data<=16'd11251;
      18404:data<=16'd10731;
      18405:data<=16'd10264;
      18406:data<=16'd10674;
      18407:data<=16'd10945;
      18408:data<=16'd9914;
      18409:data<=16'd10031;
      18410:data<=16'd11013;
      18411:data<=16'd10383;
      18412:data<=16'd9887;
      18413:data<=16'd10205;
      18414:data<=16'd9624;
      18415:data<=16'd9150;
      18416:data<=16'd9424;
      18417:data<=16'd9072;
      18418:data<=16'd9541;
      18419:data<=16'd11679;
      18420:data<=16'd9750;
      18421:data<=16'd2494;
      18422:data<=-16'd1368;
      18423:data<=-16'd399;
      18424:data<=-16'd931;
      18425:data<=-16'd1751;
      18426:data<=16'd358;
      18427:data<=16'd2998;
      18428:data<=16'd3647;
      18429:data<=16'd2861;
      18430:data<=16'd3072;
      18431:data<=16'd3949;
      18432:data<=16'd3062;
      18433:data<=16'd1892;
      18434:data<=16'd2605;
      18435:data<=16'd4347;
      18436:data<=16'd5140;
      18437:data<=16'd4094;
      18438:data<=16'd3592;
      18439:data<=16'd4461;
      18440:data<=16'd4084;
      18441:data<=16'd3086;
      18442:data<=16'd3298;
      18443:data<=16'd4123;
      18444:data<=16'd5018;
      18445:data<=16'd5483;
      18446:data<=16'd5486;
      18447:data<=16'd5359;
      18448:data<=16'd5221;
      18449:data<=16'd5072;
      18450:data<=16'd4288;
      18451:data<=16'd4531;
      18452:data<=16'd6454;
      18453:data<=16'd6589;
      18454:data<=16'd5539;
      18455:data<=16'd5573;
      18456:data<=16'd5143;
      18457:data<=16'd3936;
      18458:data<=16'd2641;
      18459:data<=16'd3256;
      18460:data<=16'd5721;
      18461:data<=16'd5618;
      18462:data<=16'd5043;
      18463:data<=16'd5172;
      18464:data<=16'd3266;
      18465:data<=16'd6922;
      18466:data<=16'd15054;
      18467:data<=16'd16195;
      18468:data<=16'd15405;
      18469:data<=16'd16783;
      18470:data<=16'd15587;
      18471:data<=16'd14778;
      18472:data<=16'd13894;
      18473:data<=16'd12163;
      18474:data<=16'd12916;
      18475:data<=16'd11934;
      18476:data<=16'd10669;
      18477:data<=16'd13120;
      18478:data<=16'd13267;
      18479:data<=16'd11591;
      18480:data<=16'd11333;
      18481:data<=16'd10254;
      18482:data<=16'd9906;
      18483:data<=16'd9947;
      18484:data<=16'd9521;
      18485:data<=16'd10178;
      18486:data<=16'd9357;
      18487:data<=16'd8652;
      18488:data<=16'd9658;
      18489:data<=16'd8050;
      18490:data<=16'd6472;
      18491:data<=16'd6760;
      18492:data<=16'd5477;
      18493:data<=16'd5773;
      18494:data<=16'd7594;
      18495:data<=16'd6578;
      18496:data<=16'd5664;
      18497:data<=16'd6390;
      18498:data<=16'd6222;
      18499:data<=16'd5673;
      18500:data<=16'd5321;
      18501:data<=16'd5165;
      18502:data<=16'd5739;
      18503:data<=16'd5941;
      18504:data<=16'd5054;
      18505:data<=16'd4531;
      18506:data<=16'd4875;
      18507:data<=16'd5092;
      18508:data<=16'd5315;
      18509:data<=16'd3786;
      18510:data<=-16'd2211;
      18511:data<=-16'd8247;
      18512:data<=-16'd9429;
      18513:data<=-16'd8624;
      18514:data<=-16'd8234;
      18515:data<=-16'd8425;
      18516:data<=-16'd9198;
      18517:data<=-16'd8416;
      18518:data<=-16'd7846;
      18519:data<=-16'd9776;
      18520:data<=-16'd10257;
      18521:data<=-16'd9770;
      18522:data<=-16'd11289;
      18523:data<=-16'd10760;
      18524:data<=-16'd8658;
      18525:data<=-16'd9550;
      18526:data<=-16'd10143;
      18527:data<=-16'd9929;
      18528:data<=-16'd13056;
      18529:data<=-16'd16193;
      18530:data<=-16'd17987;
      18531:data<=-16'd21910;
      18532:data<=-16'd24609;
      18533:data<=-16'd24125;
      18534:data<=-16'd23714;
      18535:data<=-16'd23531;
      18536:data<=-16'd23135;
      18537:data<=-16'd20157;
      18538:data<=-16'd14521;
      18539:data<=-16'd13564;
      18540:data<=-16'd15700;
      18541:data<=-16'd15197;
      18542:data<=-16'd15578;
      18543:data<=-16'd15729;
      18544:data<=-16'd14630;
      18545:data<=-16'd15767;
      18546:data<=-16'd14868;
      18547:data<=-16'd13339;
      18548:data<=-16'd13996;
      18549:data<=-16'd11474;
      18550:data<=-16'd14163;
      18551:data<=-16'd24800;
      18552:data<=-16'd27025;
      18553:data<=-16'd23482;
      18554:data<=-16'd24200;
      18555:data<=-16'd23639;
      18556:data<=-16'd21391;
      18557:data<=-16'd20098;
      18558:data<=-16'd18703;
      18559:data<=-16'd17699;
      18560:data<=-16'd16029;
      18561:data<=-16'd15847;
      18562:data<=-16'd16357;
      18563:data<=-16'd14108;
      18564:data<=-16'd14577;
      18565:data<=-16'd13124;
      18566:data<=-16'd2149;
      18567:data<=16'd5121;
      18568:data<=16'd4038;
      18569:data<=16'd4534;
      18570:data<=16'd5197;
      18571:data<=16'd4085;
      18572:data<=16'd3697;
      18573:data<=16'd3110;
      18574:data<=16'd2913;
      18575:data<=16'd2933;
      18576:data<=16'd2649;
      18577:data<=16'd2649;
      18578:data<=16'd1803;
      18579:data<=16'd1612;
      18580:data<=16'd2329;
      18581:data<=16'd1309;
      18582:data<=16'd234;
      18583:data<=16'd397;
      18584:data<=16'd928;
      18585:data<=16'd1906;
      18586:data<=16'd1838;
      18587:data<=16'd816;
      18588:data<=16'd775;
      18589:data<=16'd1186;
      18590:data<=16'd560;
      18591:data<=-16'd984;
      18592:data<=-16'd1619;
      18593:data<=-16'd1442;
      18594:data<=-16'd1210;
      18595:data<=-16'd217;
      18596:data<=-16'd422;
      18597:data<=16'd550;
      18598:data<=16'd6558;
      18599:data<=16'd9826;
      18600:data<=16'd7764;
      18601:data<=16'd7357;
      18602:data<=16'd7087;
      18603:data<=16'd5821;
      18604:data<=16'd5486;
      18605:data<=16'd4417;
      18606:data<=16'd4866;
      18607:data<=16'd6185;
      18608:data<=16'd5727;
      18609:data<=16'd6381;
      18610:data<=16'd6128;
      18611:data<=16'd4861;
      18612:data<=16'd5894;
      18613:data<=16'd5382;
      18614:data<=16'd4713;
      18615:data<=16'd3286;
      18616:data<=-16'd6507;
      18617:data<=-16'd15810;
      18618:data<=-16'd15985;
      18619:data<=-16'd14404;
      18620:data<=-16'd13088;
      18621:data<=-16'd12031;
      18622:data<=-16'd12716;
      18623:data<=-16'd11712;
      18624:data<=-16'd10636;
      18625:data<=-16'd10442;
      18626:data<=-16'd8637;
      18627:data<=-16'd8363;
      18628:data<=-16'd8956;
      18629:data<=-16'd7849;
      18630:data<=-16'd8017;
      18631:data<=-16'd8487;
      18632:data<=-16'd7544;
      18633:data<=-16'd7275;
      18634:data<=-16'd7479;
      18635:data<=-16'd7462;
      18636:data<=-16'd6913;
      18637:data<=-16'd5194;
      18638:data<=-16'd3712;
      18639:data<=-16'd4211;
      18640:data<=-16'd6034;
      18641:data<=-16'd6244;
      18642:data<=-16'd5121;
      18643:data<=-16'd5460;
      18644:data<=-16'd5074;
      18645:data<=-16'd3375;
      18646:data<=-16'd3758;
      18647:data<=-16'd4275;
      18648:data<=-16'd3243;
      18649:data<=-16'd2887;
      18650:data<=-16'd2851;
      18651:data<=-16'd2632;
      18652:data<=-16'd3074;
      18653:data<=-16'd3856;
      18654:data<=-16'd3641;
      18655:data<=-16'd2400;
      18656:data<=-16'd2535;
      18657:data<=-16'd3040;
      18658:data<=-16'd2059;
      18659:data<=-16'd1647;
      18660:data<=-16'd936;
      18661:data<=-16'd520;
      18662:data<=-16'd1366;
      18663:data<=16'd872;
      18664:data<=-16'd617;
      18665:data<=-16'd8619;
      18666:data<=-16'd5118;
      18667:data<=16'd7083;
      18668:data<=16'd8875;
      18669:data<=16'd6542;
      18670:data<=16'd7714;
      18671:data<=16'd7447;
      18672:data<=16'd7603;
      18673:data<=16'd8037;
      18674:data<=16'd6892;
      18675:data<=16'd7188;
      18676:data<=16'd7600;
      18677:data<=16'd6777;
      18678:data<=16'd5648;
      18679:data<=16'd4266;
      18680:data<=16'd4560;
      18681:data<=16'd5248;
      18682:data<=16'd4326;
      18683:data<=16'd4496;
      18684:data<=16'd5974;
      18685:data<=16'd6786;
      18686:data<=16'd6331;
      18687:data<=16'd4699;
      18688:data<=16'd3748;
      18689:data<=16'd3660;
      18690:data<=16'd2678;
      18691:data<=16'd1074;
      18692:data<=16'd347;
      18693:data<=16'd1010;
      18694:data<=16'd1459;
      18695:data<=16'd1651;
      18696:data<=16'd2823;
      18697:data<=16'd3049;
      18698:data<=16'd2775;
      18699:data<=16'd3353;
      18700:data<=16'd2810;
      18701:data<=16'd2440;
      18702:data<=16'd2335;
      18703:data<=16'd846;
      18704:data<=16'd732;
      18705:data<=16'd738;
      18706:data<=-16'd282;
      18707:data<=16'd855;
      18708:data<=16'd1692;
      18709:data<=16'd1503;
      18710:data<=16'd1967;
      18711:data<=16'd1315;
      18712:data<=16'd1632;
      18713:data<=16'd2249;
      18714:data<=16'd2082;
      18715:data<=16'd3401;
      18716:data<=-16'd2513;
      18717:data<=-16'd14671;
      18718:data<=-16'd17196;
      18719:data<=-16'd14481;
      18720:data<=-16'd14954;
      18721:data<=-16'd13949;
      18722:data<=-16'd13520;
      18723:data<=-16'd13493;
      18724:data<=-16'd10824;
      18725:data<=-16'd9784;
      18726:data<=-16'd9586;
      18727:data<=-16'd9403;
      18728:data<=-16'd10496;
      18729:data<=-16'd9897;
      18730:data<=-16'd9687;
      18731:data<=-16'd8437;
      18732:data<=-16'd1865;
      18733:data<=16'd2364;
      18734:data<=16'd1700;
      18735:data<=16'd1771;
      18736:data<=16'd1777;
      18737:data<=16'd2164;
      18738:data<=16'd3336;
      18739:data<=16'd2851;
      18740:data<=16'd2851;
      18741:data<=16'd4215;
      18742:data<=16'd5419;
      18743:data<=16'd6261;
      18744:data<=16'd5794;
      18745:data<=16'd5213;
      18746:data<=16'd5233;
      18747:data<=16'd4282;
      18748:data<=16'd3952;
      18749:data<=16'd5233;
      18750:data<=16'd5739;
      18751:data<=16'd5046;
      18752:data<=16'd5310;
      18753:data<=16'd6501;
      18754:data<=16'd6702;
      18755:data<=16'd7247;
      18756:data<=16'd8231;
      18757:data<=16'd7338;
      18758:data<=16'd7019;
      18759:data<=16'd7433;
      18760:data<=16'd6311;
      18761:data<=16'd6334;
      18762:data<=16'd6842;
      18763:data<=16'd6839;
      18764:data<=16'd7037;
      18765:data<=16'd5752;
      18766:data<=16'd11188;
      18767:data<=16'd24107;
      18768:data<=16'd27425;
      18769:data<=16'd23846;
      18770:data<=16'd24665;
      18771:data<=16'd23570;
      18772:data<=16'd21541;
      18773:data<=16'd22381;
      18774:data<=16'd21200;
      18775:data<=16'd20169;
      18776:data<=16'd19737;
      18777:data<=16'd18265;
      18778:data<=16'd19117;
      18779:data<=16'd19076;
      18780:data<=16'd17523;
      18781:data<=16'd18348;
      18782:data<=16'd17723;
      18783:data<=16'd15600;
      18784:data<=16'd15587;
      18785:data<=16'd15814;
      18786:data<=16'd15292;
      18787:data<=16'd13960;
      18788:data<=16'd12533;
      18789:data<=16'd12369;
      18790:data<=16'd12314;
      18791:data<=16'd12831;
      18792:data<=16'd13150;
      18793:data<=16'd11630;
      18794:data<=16'd11389;
      18795:data<=16'd12149;
      18796:data<=16'd11681;
      18797:data<=16'd11750;
      18798:data<=16'd9718;
      18799:data<=16'd3539;
      18800:data<=-16'd528;
      18801:data<=16'd79;
      18802:data<=16'd1115;
      18803:data<=16'd1833;
      18804:data<=16'd3137;
      18805:data<=16'd3124;
      18806:data<=16'd2858;
      18807:data<=16'd3454;
      18808:data<=16'd2578;
      18809:data<=16'd2156;
      18810:data<=16'd2596;
      18811:data<=16'd1133;
      18812:data<=16'd870;
      18813:data<=16'd811;
      18814:data<=16'd262;
      18815:data<=16'd3811;
      18816:data<=16'd898;
      18817:data<=-16'd11994;
      18818:data<=-16'd16433;
      18819:data<=-16'd13532;
      18820:data<=-16'd14531;
      18821:data<=-16'd13957;
      18822:data<=-16'd12369;
      18823:data<=-16'd12747;
      18824:data<=-16'd10862;
      18825:data<=-16'd9734;
      18826:data<=-16'd10440;
      18827:data<=-16'd9749;
      18828:data<=-16'd9553;
      18829:data<=-16'd8957;
      18830:data<=-16'd7163;
      18831:data<=-16'd7322;
      18832:data<=-16'd7832;
      18833:data<=-16'd6576;
      18834:data<=-16'd6053;
      18835:data<=-16'd6740;
      18836:data<=-16'd6363;
      18837:data<=-16'd5391;
      18838:data<=-16'd5363;
      18839:data<=-16'd5288;
      18840:data<=-16'd4226;
      18841:data<=-16'd2399;
      18842:data<=-16'd1022;
      18843:data<=-16'd981;
      18844:data<=-16'd299;
      18845:data<=16'd391;
      18846:data<=-16'd781;
      18847:data<=-16'd1028;
      18848:data<=-16'd238;
      18849:data<=16'd209;
      18850:data<=16'd919;
      18851:data<=16'd218;
      18852:data<=16'd429;
      18853:data<=16'd2798;
      18854:data<=16'd2616;
      18855:data<=16'd1991;
      18856:data<=16'd2541;
      18857:data<=16'd1615;
      18858:data<=16'd2000;
      18859:data<=16'd2587;
      18860:data<=16'd1353;
      18861:data<=16'd1477;
      18862:data<=16'd1983;
      18863:data<=16'd2343;
      18864:data<=16'd1706;
      18865:data<=16'd1789;
      18866:data<=16'd12836;
      18867:data<=16'd27419;
      18868:data<=16'd29329;
      18869:data<=16'd26837;
      18870:data<=16'd27539;
      18871:data<=16'd25949;
      18872:data<=16'd24080;
      18873:data<=16'd23123;
      18874:data<=16'd21303;
      18875:data<=16'd20912;
      18876:data<=16'd20785;
      18877:data<=16'd20034;
      18878:data<=16'd20659;
      18879:data<=16'd20930;
      18880:data<=16'd19352;
      18881:data<=16'd18111;
      18882:data<=16'd17887;
      18883:data<=16'd16832;
      18884:data<=16'd15531;
      18885:data<=16'd15101;
      18886:data<=16'd14377;
      18887:data<=16'd14152;
      18888:data<=16'd13615;
      18889:data<=16'd11038;
      18890:data<=16'd10725;
      18891:data<=16'd12493;
      18892:data<=16'd11638;
      18893:data<=16'd10598;
      18894:data<=16'd10455;
      18895:data<=16'd9433;
      18896:data<=16'd9030;
      18897:data<=16'd8490;
      18898:data<=16'd7218;
      18899:data<=16'd6570;
      18900:data<=16'd6363;
      18901:data<=16'd6522;
      18902:data<=16'd5937;
      18903:data<=16'd5542;
      18904:data<=16'd6828;
      18905:data<=16'd6169;
      18906:data<=16'd4698;
      18907:data<=16'd5347;
      18908:data<=16'd4360;
      18909:data<=16'd2963;
      18910:data<=16'd3159;
      18911:data<=16'd2071;
      18912:data<=16'd1738;
      18913:data<=16'd1941;
      18914:data<=16'd1583;
      18915:data<=16'd3802;
      18916:data<=16'd1309;
      18917:data<=-16'd9529;
      18918:data<=-16'd15805;
      18919:data<=-16'd15171;
      18920:data<=-16'd15273;
      18921:data<=-16'd14941;
      18922:data<=-16'd13473;
      18923:data<=-16'd13136;
      18924:data<=-16'd13027;
      18925:data<=-16'd12698;
      18926:data<=-16'd12419;
      18927:data<=-16'd12216;
      18928:data<=-16'd11602;
      18929:data<=-16'd10047;
      18930:data<=-16'd8698;
      18931:data<=-16'd8379;
      18932:data<=-16'd11197;
      18933:data<=-16'd17033;
      18934:data<=-16'd18900;
      18935:data<=-16'd16788;
      18936:data<=-16'd17290;
      18937:data<=-16'd18077;
      18938:data<=-16'd16917;
      18939:data<=-16'd16557;
      18940:data<=-16'd15637;
      18941:data<=-16'd14339;
      18942:data<=-16'd14586;
      18943:data<=-16'd14422;
      18944:data<=-16'd13426;
      18945:data<=-16'd12972;
      18946:data<=-16'd13215;
      18947:data<=-16'd13295;
      18948:data<=-16'd11885;
      18949:data<=-16'd10419;
      18950:data<=-16'd10592;
      18951:data<=-16'd10945;
      18952:data<=-16'd10484;
      18953:data<=-16'd9881;
      18954:data<=-16'd10342;
      18955:data<=-16'd11444;
      18956:data<=-16'd11309;
      18957:data<=-16'd10552;
      18958:data<=-16'd10103;
      18959:data<=-16'd9875;
      18960:data<=-16'd10009;
      18961:data<=-16'd9653;
      18962:data<=-16'd9545;
      18963:data<=-16'd9345;
      18964:data<=-16'd8483;
      18965:data<=-16'd10807;
      18966:data<=-16'd10759;
      18967:data<=-16'd752;
      18968:data<=16'd7385;
      18969:data<=16'd6727;
      18970:data<=16'd6554;
      18971:data<=16'd7395;
      18972:data<=16'd6429;
      18973:data<=16'd6222;
      18974:data<=16'd6100;
      18975:data<=16'd5827;
      18976:data<=16'd5724;
      18977:data<=16'd5080;
      18978:data<=16'd4614;
      18979:data<=16'd3239;
      18980:data<=16'd1659;
      18981:data<=16'd1982;
      18982:data<=16'd2314;
      18983:data<=16'd2087;
      18984:data<=16'd2153;
      18985:data<=16'd2255;
      18986:data<=16'd2400;
      18987:data<=16'd1556;
      18988:data<=16'd795;
      18989:data<=16'd1068;
      18990:data<=16'd159;
      18991:data<=-16'd1043;
      18992:data<=-16'd1560;
      18993:data<=-16'd2071;
      18994:data<=-16'd1977;
      18995:data<=-16'd2423;
      18996:data<=-16'd2137;
      18997:data<=-16'd1272;
      18998:data<=-16'd3362;
      18999:data<=-16'd1911;
      19000:data<=16'd4996;
      19001:data<=16'd6930;
      19002:data<=16'd5424;
      19003:data<=16'd5351;
      19004:data<=16'd3378;
      19005:data<=16'd1765;
      19006:data<=16'd1845;
      19007:data<=16'd1365;
      19008:data<=16'd1327;
      19009:data<=16'd1010;
      19010:data<=16'd940;
      19011:data<=16'd1416;
      19012:data<=16'd829;
      19013:data<=16'd1381;
      19014:data<=16'd1845;
      19015:data<=16'd1318;
      19016:data<=16'd743;
      19017:data<=-16'd6884;
      19018:data<=-16'd17479;
      19019:data<=-16'd19058;
      19020:data<=-16'd17553;
      19021:data<=-16'd17596;
      19022:data<=-16'd15719;
      19023:data<=-16'd15277;
      19024:data<=-16'd15346;
      19025:data<=-16'd14287;
      19026:data<=-16'd14565;
      19027:data<=-16'd13585;
      19028:data<=-16'd13312;
      19029:data<=-16'd15594;
      19030:data<=-16'd14792;
      19031:data<=-16'd12915;
      19032:data<=-16'd13352;
      19033:data<=-16'd12927;
      19034:data<=-16'd12040;
      19035:data<=-16'd11697;
      19036:data<=-16'd11110;
      19037:data<=-16'd10798;
      19038:data<=-16'd10557;
      19039:data<=-16'd10261;
      19040:data<=-16'd9999;
      19041:data<=-16'd10481;
      19042:data<=-16'd11312;
      19043:data<=-16'd10320;
      19044:data<=-16'd9447;
      19045:data<=-16'd9433;
      19046:data<=-16'd8413;
      19047:data<=-16'd9116;
      19048:data<=-16'd9994;
      19049:data<=-16'd7944;
      19050:data<=-16'd7371;
      19051:data<=-16'd8053;
      19052:data<=-16'd7194;
      19053:data<=-16'd7238;
      19054:data<=-16'd7985;
      19055:data<=-16'd7971;
      19056:data<=-16'd7389;
      19057:data<=-16'd6725;
      19058:data<=-16'd6410;
      19059:data<=-16'd5369;
      19060:data<=-16'd5389;
      19061:data<=-16'd5924;
      19062:data<=-16'd3997;
      19063:data<=-16'd4276;
      19064:data<=-16'd4808;
      19065:data<=-16'd3001;
      19066:data<=-16'd8194;
      19067:data<=-16'd10302;
      19068:data<=16'd1216;
      19069:data<=16'd6056;
      19070:data<=16'd1654;
      19071:data<=16'd2927;
      19072:data<=16'd3547;
      19073:data<=16'd2162;
      19074:data<=16'd4090;
      19075:data<=16'd3648;
      19076:data<=16'd2372;
      19077:data<=16'd3107;
      19078:data<=16'd2535;
      19079:data<=16'd1730;
      19080:data<=16'd763;
      19081:data<=16'd572;
      19082:data<=16'd2449;
      19083:data<=16'd2005;
      19084:data<=16'd123;
      19085:data<=16'd485;
      19086:data<=16'd1333;
      19087:data<=16'd1532;
      19088:data<=16'd1162;
      19089:data<=16'd1122;
      19090:data<=16'd1158;
      19091:data<=-16'd576;
      19092:data<=-16'd1124;
      19093:data<=16'd144;
      19094:data<=-16'd203;
      19095:data<=-16'd441;
      19096:data<=-16'd264;
      19097:data<=-16'd1289;
      19098:data<=-16'd1228;
      19099:data<=-16'd811;
      19100:data<=-16'd1858;
      19101:data<=-16'd2044;
      19102:data<=-16'd1113;
      19103:data<=-16'd1680;
      19104:data<=-16'd3240;
      19105:data<=-16'd3371;
      19106:data<=-16'd2943;
      19107:data<=-16'd2801;
      19108:data<=-16'd2282;
      19109:data<=-16'd2537;
      19110:data<=-16'd2137;
      19111:data<=-16'd823;
      19112:data<=-16'd1465;
      19113:data<=-16'd1316;
      19114:data<=-16'd811;
      19115:data<=-16'd1398;
      19116:data<=16'd860;
      19117:data<=-16'd3403;
      19118:data<=-16'd16804;
      19119:data<=-16'd20653;
      19120:data<=-16'd16816;
      19121:data<=-16'd17315;
      19122:data<=-16'd16530;
      19123:data<=-16'd15074;
      19124:data<=-16'd15371;
      19125:data<=-16'd13800;
      19126:data<=-16'd13556;
      19127:data<=-16'd13170;
      19128:data<=-16'd11652;
      19129:data<=-16'd13241;
      19130:data<=-16'd13082;
      19131:data<=-16'd11314;
      19132:data<=-16'd12096;
      19133:data<=-16'd8974;
      19134:data<=-16'd2497;
      19135:data<=-16'd2;
      19136:data<=-16'd232;
      19137:data<=-16'd162;
      19138:data<=16'd80;
      19139:data<=16'd115;
      19140:data<=16'd908;
      19141:data<=16'd2156;
      19142:data<=16'd1595;
      19143:data<=16'd1034;
      19144:data<=16'd1949;
      19145:data<=16'd2332;
      19146:data<=16'd2651;
      19147:data<=16'd3039;
      19148:data<=16'd2922;
      19149:data<=16'd3113;
      19150:data<=16'd3692;
      19151:data<=16'd4605;
      19152:data<=16'd4605;
      19153:data<=16'd4770;
      19154:data<=16'd7110;
      19155:data<=16'd7852;
      19156:data<=16'd6887;
      19157:data<=16'd7209;
      19158:data<=16'd6971;
      19159:data<=16'd6680;
      19160:data<=16'd6607;
      19161:data<=16'd6144;
      19162:data<=16'd6586;
      19163:data<=16'd6026;
      19164:data<=16'd6689;
      19165:data<=16'd8204;
      19166:data<=16'd6109;
      19167:data<=16'd11365;
      19168:data<=16'd24318;
      19169:data<=16'd27216;
      19170:data<=16'd24457;
      19171:data<=16'd25049;
      19172:data<=16'd23739;
      19173:data<=16'd22557;
      19174:data<=16'd22156;
      19175:data<=16'd20301;
      19176:data<=16'd20433;
      19177:data<=16'd20284;
      19178:data<=16'd18827;
      19179:data<=16'd19317;
      19180:data<=16'd19870;
      19181:data<=16'd19317;
      19182:data<=16'd18360;
      19183:data<=16'd17649;
      19184:data<=16'd17473;
      19185:data<=16'd16543;
      19186:data<=16'd15887;
      19187:data<=16'd15318;
      19188:data<=16'd14445;
      19189:data<=16'd15023;
      19190:data<=16'd14064;
      19191:data<=16'd12396;
      19192:data<=16'd14305;
      19193:data<=16'd15414;
      19194:data<=16'd14135;
      19195:data<=16'd13967;
      19196:data<=16'd13723;
      19197:data<=16'd12057;
      19198:data<=16'd10349;
      19199:data<=16'd10621;
      19200:data<=16'd9222;
      19201:data<=16'd3015;
      19202:data<=16'd437;
      19203:data<=16'd2090;
      19204:data<=16'd873;
      19205:data<=16'd1209;
      19206:data<=16'd2807;
      19207:data<=16'd1668;
      19208:data<=16'd2065;
      19209:data<=16'd2349;
      19210:data<=16'd1213;
      19211:data<=16'd1386;
      19212:data<=16'd1272;
      19213:data<=16'd2249;
      19214:data<=16'd2035;
      19215:data<=-16'd206;
      19216:data<=16'd2464;
      19217:data<=16'd960;
      19218:data<=-16'd10410;
      19219:data<=-16'd15339;
      19220:data<=-16'd13218;
      19221:data<=-16'd13772;
      19222:data<=-16'd13361;
      19223:data<=-16'd12320;
      19224:data<=-16'd12889;
      19225:data<=-16'd11893;
      19226:data<=-16'd10777;
      19227:data<=-16'd10777;
      19228:data<=-16'd9994;
      19229:data<=-16'd8317;
      19230:data<=-16'd6898;
      19231:data<=-16'd6576;
      19232:data<=-16'd6366;
      19233:data<=-16'd6531;
      19234:data<=-16'd7598;
      19235:data<=-16'd7218;
      19236:data<=-16'd6216;
      19237:data<=-16'd6161;
      19238:data<=-16'd5551;
      19239:data<=-16'd5219;
      19240:data<=-16'd5015;
      19241:data<=-16'd3383;
      19242:data<=-16'd2137;
      19243:data<=-16'd2012;
      19244:data<=-16'd2056;
      19245:data<=-16'd2065;
      19246:data<=-16'd1744;
      19247:data<=-16'd1312;
      19248:data<=-16'd851;
      19249:data<=-16'd987;
      19250:data<=-16'd1298;
      19251:data<=-16'd9;
      19252:data<=16'd505;
      19253:data<=-16'd94;
      19254:data<=16'd1750;
      19255:data<=16'd3366;
      19256:data<=16'd2799;
      19257:data<=16'd2746;
      19258:data<=16'd2573;
      19259:data<=16'd2150;
      19260:data<=16'd2287;
      19261:data<=16'd2229;
      19262:data<=16'd1864;
      19263:data<=16'd978;
      19264:data<=16'd2029;
      19265:data<=16'd3372;
      19266:data<=16'd1246;
      19267:data<=16'd7265;
      19268:data<=16'd23704;
      19269:data<=16'd30635;
      19270:data<=16'd27802;
      19271:data<=16'd27801;
      19272:data<=16'd26880;
      19273:data<=16'd24577;
      19274:data<=16'd24509;
      19275:data<=16'd23175;
      19276:data<=16'd21473;
      19277:data<=16'd20666;
      19278:data<=16'd19525;
      19279:data<=16'd19622;
      19280:data<=16'd19476;
      19281:data<=16'd18019;
      19282:data<=16'd17054;
      19283:data<=16'd16042;
      19284:data<=16'd15541;
      19285:data<=16'd15961;
      19286:data<=16'd15491;
      19287:data<=16'd14451;
      19288:data<=16'd13867;
      19289:data<=16'd13515;
      19290:data<=16'd12945;
      19291:data<=16'd12885;
      19292:data<=16'd14070;
      19293:data<=16'd14014;
      19294:data<=16'd12299;
      19295:data<=16'd11609;
      19296:data<=16'd11144;
      19297:data<=16'd10434;
      19298:data<=16'd10267;
      19299:data<=16'd9602;
      19300:data<=16'd9113;
      19301:data<=16'd8504;
      19302:data<=16'd6739;
      19303:data<=16'd6197;
      19304:data<=16'd6839;
      19305:data<=16'd6865;
      19306:data<=16'd6777;
      19307:data<=16'd6237;
      19308:data<=16'd5394;
      19309:data<=16'd4910;
      19310:data<=16'd4404;
      19311:data<=16'd4005;
      19312:data<=16'd3439;
      19313:data<=16'd3394;
      19314:data<=16'd3579;
      19315:data<=16'd2429;
      19316:data<=16'd2957;
      19317:data<=16'd2602;
      19318:data<=-16'd5876;
      19319:data<=-16'd14401;
      19320:data<=-16'd14716;
      19321:data<=-16'd13761;
      19322:data<=-16'd13913;
      19323:data<=-16'd12963;
      19324:data<=-16'd13355;
      19325:data<=-16'd13955;
      19326:data<=-16'd13035;
      19327:data<=-16'd12417;
      19328:data<=-16'd12372;
      19329:data<=-16'd11511;
      19330:data<=-16'd9447;
      19331:data<=-16'd8651;
      19332:data<=-16'd8790;
      19333:data<=-16'd7577;
      19334:data<=-16'd10108;
      19335:data<=-16'd16219;
      19336:data<=-16'd17646;
      19337:data<=-16'd16710;
      19338:data<=-16'd17070;
      19339:data<=-16'd16175;
      19340:data<=-16'd15743;
      19341:data<=-16'd15203;
      19342:data<=-16'd13620;
      19343:data<=-16'd14333;
      19344:data<=-16'd14753;
      19345:data<=-16'd13439;
      19346:data<=-16'd13315;
      19347:data<=-16'd13160;
      19348:data<=-16'd13315;
      19349:data<=-16'd13597;
      19350:data<=-16'd11776;
      19351:data<=-16'd11007;
      19352:data<=-16'd11732;
      19353:data<=-16'd10921;
      19354:data<=-16'd10534;
      19355:data<=-16'd11555;
      19356:data<=-16'd11775;
      19357:data<=-16'd10945;
      19358:data<=-16'd10903;
      19359:data<=-16'd11506;
      19360:data<=-16'd10511;
      19361:data<=-16'd9382;
      19362:data<=-16'd9291;
      19363:data<=-16'd9130;
      19364:data<=-16'd10047;
      19365:data<=-16'd9671;
      19366:data<=-16'd8601;
      19367:data<=-16'd10243;
      19368:data<=-16'd5186;
      19369:data<=16'd5959;
      19370:data<=16'd7835;
      19371:data<=16'd5366;
      19372:data<=16'd6651;
      19373:data<=16'd5665;
      19374:data<=16'd5001;
      19375:data<=16'd6445;
      19376:data<=16'd5125;
      19377:data<=16'd4407;
      19378:data<=16'd5316;
      19379:data<=16'd3912;
      19380:data<=16'd1757;
      19381:data<=16'd1336;
      19382:data<=16'd1689;
      19383:data<=16'd995;
      19384:data<=16'd419;
      19385:data<=16'd889;
      19386:data<=16'd663;
      19387:data<=16'd972;
      19388:data<=16'd1572;
      19389:data<=16'd848;
      19390:data<=16'd1295;
      19391:data<=16'd1321;
      19392:data<=-16'd400;
      19393:data<=-16'd904;
      19394:data<=-16'd1902;
      19395:data<=-16'd2472;
      19396:data<=-16'd1175;
      19397:data<=-16'd2121;
      19398:data<=-16'd2670;
      19399:data<=-16'd1527;
      19400:data<=-16'd2628;
      19401:data<=-16'd875;
      19402:data<=16'd4898;
      19403:data<=16'd6714;
      19404:data<=16'd4631;
      19405:data<=16'd3278;
      19406:data<=16'd2795;
      19407:data<=16'd1867;
      19408:data<=16'd1175;
      19409:data<=16'd1213;
      19410:data<=16'd764;
      19411:data<=16'd910;
      19412:data<=16'd1162;
      19413:data<=16'd373;
      19414:data<=16'd1666;
      19415:data<=16'd1945;
      19416:data<=-16'd41;
      19417:data<=16'd746;
      19418:data<=-16'd4802;
      19419:data<=-16'd17811;
      19420:data<=-16'd20776;
      19421:data<=-16'd17064;
      19422:data<=-16'd17687;
      19423:data<=-16'd17500;
      19424:data<=-16'd16404;
      19425:data<=-16'd15929;
      19426:data<=-16'd14640;
      19427:data<=-16'd15599;
      19428:data<=-16'd15528;
      19429:data<=-16'd13274;
      19430:data<=-16'd14004;
      19431:data<=-16'd14522;
      19432:data<=-16'd13265;
      19433:data<=-16'd13101;
      19434:data<=-16'd12249;
      19435:data<=-16'd11388;
      19436:data<=-16'd11405;
      19437:data<=-16'd10869;
      19438:data<=-16'd11109;
      19439:data<=-16'd11291;
      19440:data<=-16'd10288;
      19441:data<=-16'd10016;
      19442:data<=-16'd10443;
      19443:data<=-16'd10954;
      19444:data<=-16'd11303;
      19445:data<=-16'd10919;
      19446:data<=-16'd10364;
      19447:data<=-16'd9875;
      19448:data<=-16'd9636;
      19449:data<=-16'd9320;
      19450:data<=-16'd8311;
      19451:data<=-16'd8049;
      19452:data<=-16'd8150;
      19453:data<=-16'd6980;
      19454:data<=-16'd6405;
      19455:data<=-16'd7602;
      19456:data<=-16'd8382;
      19457:data<=-16'd7485;
      19458:data<=-16'd6946;
      19459:data<=-16'd7671;
      19460:data<=-16'd7109;
      19461:data<=-16'd5770;
      19462:data<=-16'd5382;
      19463:data<=-16'd5069;
      19464:data<=-16'd5673;
      19465:data<=-16'd5328;
      19466:data<=-16'd3570;
      19467:data<=-16'd5277;
      19468:data<=-16'd4387;
      19469:data<=16'd3083;
      19470:data<=16'd5212;
      19471:data<=16'd2833;
      19472:data<=16'd4519;
      19473:data<=16'd5115;
      19474:data<=16'd3762;
      19475:data<=16'd3823;
      19476:data<=16'd3218;
      19477:data<=16'd3653;
      19478:data<=16'd4657;
      19479:data<=16'd3277;
      19480:data<=16'd1798;
      19481:data<=16'd834;
      19482:data<=16'd475;
      19483:data<=16'd1366;
      19484:data<=16'd1392;
      19485:data<=16'd1143;
      19486:data<=16'd1472;
      19487:data<=16'd1595;
      19488:data<=16'd1945;
      19489:data<=16'd1468;
      19490:data<=16'd1412;
      19491:data<=16'd2810;
      19492:data<=16'd1535;
      19493:data<=-16'd867;
      19494:data<=-16'd405;
      19495:data<=-16'd23;
      19496:data<=-16'd133;
      19497:data<=16'd785;
      19498:data<=16'd234;
      19499:data<=-16'd575;
      19500:data<=16'd917;
      19501:data<=16'd1507;
      19502:data<=16'd346;
      19503:data<=16'd422;
      19504:data<=-16'd35;
      19505:data<=-16'd1859;
      19506:data<=-16'd1713;
      19507:data<=-16'd1210;
      19508:data<=-16'd1996;
      19509:data<=-16'd1707;
      19510:data<=-16'd1318;
      19511:data<=-16'd1462;
      19512:data<=-16'd1365;
      19513:data<=-16'd1149;
      19514:data<=16'd94;
      19515:data<=-16'd520;
      19516:data<=-16'd1736;
      19517:data<=16'd569;
      19518:data<=-16'd4270;
      19519:data<=-16'd17324;
      19520:data<=-16'd20973;
      19521:data<=-16'd17391;
      19522:data<=-16'd17602;
      19523:data<=-16'd17452;
      19524:data<=-16'd15985;
      19525:data<=-16'd15203;
      19526:data<=-16'd13718;
      19527:data<=-16'd13214;
      19528:data<=-16'd12824;
      19529:data<=-16'd11909;
      19530:data<=-16'd12957;
      19531:data<=-16'd13723;
      19532:data<=-16'd12099;
      19533:data<=-16'd11206;
      19534:data<=-16'd11740;
      19535:data<=-16'd8504;
      19536:data<=-16'd1821;
      19537:data<=16'd390;
      19538:data<=-16'd417;
      19539:data<=16'd614;
      19540:data<=16'd267;
      19541:data<=16'd156;
      19542:data<=16'd1685;
      19543:data<=16'd960;
      19544:data<=16'd857;
      19545:data<=16'd2149;
      19546:data<=16'd1880;
      19547:data<=16'd1759;
      19548:data<=16'd1433;
      19549:data<=16'd1688;
      19550:data<=16'd3334;
      19551:data<=16'd3101;
      19552:data<=16'd2867;
      19553:data<=16'd3571;
      19554:data<=16'd3422;
      19555:data<=16'd4425;
      19556:data<=16'd5092;
      19557:data<=16'd5236;
      19558:data<=16'd6705;
      19559:data<=16'd6737;
      19560:data<=16'd6434;
      19561:data<=16'd6543;
      19562:data<=16'd5762;
      19563:data<=16'd6138;
      19564:data<=16'd5829;
      19565:data<=16'd6184;
      19566:data<=16'd7859;
      19567:data<=16'd5835;
      19568:data<=16'd10129;
      19569:data<=16'd23282;
      19570:data<=16'd27395;
      19571:data<=16'd24745;
      19572:data<=16'd25146;
      19573:data<=16'd23927;
      19574:data<=16'd22569;
      19575:data<=16'd22172;
      19576:data<=16'd20481;
      19577:data<=16'd20287;
      19578:data<=16'd19729;
      19579:data<=16'd18882;
      19580:data<=16'd20071;
      19581:data<=16'd20216;
      19582:data<=16'd19930;
      19583:data<=16'd19713;
      19584:data<=16'd18272;
      19585:data<=16'd17629;
      19586:data<=16'd17115;
      19587:data<=16'd16424;
      19588:data<=16'd15890;
      19589:data<=16'd14757;
      19590:data<=16'd15013;
      19591:data<=16'd14971;
      19592:data<=16'd13973;
      19593:data<=16'd14736;
      19594:data<=16'd14366;
      19595:data<=16'd13591;
      19596:data<=16'd13944;
      19597:data<=16'd12530;
      19598:data<=16'd12495;
      19599:data<=16'd12604;
      19600:data<=16'd10378;
      19601:data<=16'd10687;
      19602:data<=16'd8313;
      19603:data<=16'd1709;
      19604:data<=16'd399;
      19605:data<=16'd1312;
      19606:data<=16'd1304;
      19607:data<=16'd2905;
      19608:data<=16'd2199;
      19609:data<=16'd843;
      19610:data<=16'd1623;
      19611:data<=16'd1789;
      19612:data<=16'd1811;
      19613:data<=16'd1427;
      19614:data<=16'd1545;
      19615:data<=16'd2315;
      19616:data<=16'd1078;
      19617:data<=16'd1835;
      19618:data<=16'd681;
      19619:data<=-16'd9348;
      19620:data<=-16'd15543;
      19621:data<=-16'd13408;
      19622:data<=-16'd13869;
      19623:data<=-16'd14505;
      19624:data<=-16'd12175;
      19625:data<=-16'd11606;
      19626:data<=-16'd11897;
      19627:data<=-16'd11556;
      19628:data<=-16'd10933;
      19629:data<=-16'd10047;
      19630:data<=-16'd9256;
      19631:data<=-16'd7897;
      19632:data<=-16'd7388;
      19633:data<=-16'd7562;
      19634:data<=-16'd6458;
      19635:data<=-16'd6152;
      19636:data<=-16'd6197;
      19637:data<=-16'd5565;
      19638:data<=-16'd6335;
      19639:data<=-16'd6219;
      19640:data<=-16'd5131;
      19641:data<=-16'd5354;
      19642:data<=-16'd3624;
      19643:data<=-16'd1064;
      19644:data<=-16'd1152;
      19645:data<=-16'd1456;
      19646:data<=-16'd1313;
      19647:data<=-16'd1319;
      19648:data<=-16'd1169;
      19649:data<=-16'd1463;
      19650:data<=-16'd1099;
      19651:data<=-16'd708;
      19652:data<=-16'd1039;
      19653:data<=-16'd432;
      19654:data<=16'd129;
      19655:data<=16'd817;
      19656:data<=16'd1855;
      19657:data<=16'd1333;
      19658:data<=16'd1723;
      19659:data<=16'd2963;
      19660:data<=16'd2684;
      19661:data<=16'd3153;
      19662:data<=16'd2892;
      19663:data<=16'd1577;
      19664:data<=16'd2405;
      19665:data<=16'd2842;
      19666:data<=16'd2786;
      19667:data<=16'd2792;
      19668:data<=16'd4411;
      19669:data<=16'd16228;
      19670:data<=16'd29731;
      19671:data<=16'd30365;
      19672:data<=16'd27795;
      19673:data<=16'd27869;
      19674:data<=16'd25713;
      19675:data<=16'd24967;
      19676:data<=16'd24222;
      19677:data<=16'd22045;
      19678:data<=16'd22516;
      19679:data<=16'd22250;
      19680:data<=16'd21347;
      19681:data<=16'd22319;
      19682:data<=16'd21892;
      19683:data<=16'd21153;
      19684:data<=16'd20263;
      19685:data<=16'd18036;
      19686:data<=16'd17625;
      19687:data<=16'd17608;
      19688:data<=16'd16553;
      19689:data<=16'd16217;
      19690:data<=16'd15355;
      19691:data<=16'd14004;
      19692:data<=16'd13194;
      19693:data<=16'd13447;
      19694:data<=16'd14193;
      19695:data<=16'd13112;
      19696:data<=16'd12486;
      19697:data<=16'd12516;
      19698:data<=16'd10511;
      19699:data<=16'd10205;
      19700:data<=16'd10205;
      19701:data<=16'd7744;
      19702:data<=16'd7990;
      19703:data<=16'd8338;
      19704:data<=16'd5973;
      19705:data<=16'd6369;
      19706:data<=16'd8087;
      19707:data<=16'd8217;
      19708:data<=16'd7527;
      19709:data<=16'd5504;
      19710:data<=16'd4328;
      19711:data<=16'd4573;
      19712:data<=16'd4443;
      19713:data<=16'd4094;
      19714:data<=16'd3415;
      19715:data<=16'd2952;
      19716:data<=16'd2258;
      19717:data<=16'd2455;
      19718:data<=16'd3604;
      19719:data<=-16'd2854;
      19720:data<=-16'd13338;
      19721:data<=-16'd14562;
      19722:data<=-16'd12663;
      19723:data<=-16'd14105;
      19724:data<=-16'd13732;
      19725:data<=-16'd13230;
      19726:data<=-16'd12904;
      19727:data<=-16'd11486;
      19728:data<=-16'd12140;
      19729:data<=-16'd12405;
      19730:data<=-16'd11276;
      19731:data<=-16'd10695;
      19732:data<=-16'd9680;
      19733:data<=-16'd10044;
      19734:data<=-16'd10102;
      19735:data<=-16'd8225;
      19736:data<=-16'd10845;
      19737:data<=-16'd16477;
      19738:data<=-16'd17866;
      19739:data<=-16'd16785;
      19740:data<=-16'd16509;
      19741:data<=-16'd16283;
      19742:data<=-16'd15396;
      19743:data<=-16'd14469;
      19744:data<=-16'd14013;
      19745:data<=-16'd13682;
      19746:data<=-16'd13981;
      19747:data<=-16'd14220;
      19748:data<=-16'd13617;
      19749:data<=-16'd13527;
      19750:data<=-16'd12850;
      19751:data<=-16'd11565;
      19752:data<=-16'd11872;
      19753:data<=-16'd11758;
      19754:data<=-16'd10727;
      19755:data<=-16'd10965;
      19756:data<=-16'd11869;
      19757:data<=-16'd12625;
      19758:data<=-16'd12207;
      19759:data<=-16'd10956;
      19760:data<=-16'd10525;
      19761:data<=-16'd9909;
      19762:data<=-16'd9514;
      19763:data<=-16'd9538;
      19764:data<=-16'd9003;
      19765:data<=-16'd9260;
      19766:data<=-16'd8536;
      19767:data<=-16'd8434;
      19768:data<=-16'd11297;
      19769:data<=-16'd6100;
      19770:data<=16'd6169;
      19771:data<=16'd8740;
      19772:data<=16'd5527;
      19773:data<=16'd6351;
      19774:data<=16'd6529;
      19775:data<=16'd6090;
      19776:data<=16'd6564;
      19777:data<=16'd5215;
      19778:data<=16'd4755;
      19779:data<=16'd5770;
      19780:data<=16'd4625;
      19781:data<=16'd2065;
      19782:data<=16'd846;
      19783:data<=16'd1568;
      19784:data<=16'd2256;
      19785:data<=16'd1463;
      19786:data<=16'd473;
      19787:data<=16'd406;
      19788:data<=16'd1054;
      19789:data<=16'd1168;
      19790:data<=16'd584;
      19791:data<=16'd723;
      19792:data<=16'd534;
      19793:data<=-16'd699;
      19794:data<=-16'd1397;
      19795:data<=-16'd2006;
      19796:data<=-16'd2544;
      19797:data<=-16'd2044;
      19798:data<=-16'd1657;
      19799:data<=-16'd1647;
      19800:data<=-16'd1418;
      19801:data<=-16'd1936;
      19802:data<=-16'd2535;
      19803:data<=16'd355;
      19804:data<=16'd5553;
      19805:data<=16'd6020;
      19806:data<=16'd2952;
      19807:data<=16'd2641;
      19808:data<=16'd2525;
      19809:data<=16'd1606;
      19810:data<=16'd2341;
      19811:data<=16'd1848;
      19812:data<=16'd1278;
      19813:data<=16'd1883;
      19814:data<=16'd1002;
      19815:data<=16'd1160;
      19816:data<=16'd1017;
      19817:data<=16'd20;
      19818:data<=16'd1824;
      19819:data<=-16'd3783;
      19820:data<=-16'd17133;
      19821:data<=-16'd20313;
      19822:data<=-16'd17036;
      19823:data<=-16'd17699;
      19824:data<=-16'd16959;
      19825:data<=-16'd15719;
      19826:data<=-16'd15778;
      19827:data<=-16'd14122;
      19828:data<=-16'd13277;
      19829:data<=-16'd12971;
      19830:data<=-16'd12974;
      19831:data<=-16'd14910;
      19832:data<=-16'd15064;
      19833:data<=-16'd14207;
      19834:data<=-16'd14293;
      19835:data<=-16'd12536;
      19836:data<=-16'd11615;
      19837:data<=-16'd12819;
      19838:data<=-16'd12084;
      19839:data<=-16'd10619;
      19840:data<=-16'd10568;
      19841:data<=-16'd10263;
      19842:data<=-16'd9658;
      19843:data<=-16'd10304;
      19844:data<=-16'd11242;
      19845:data<=-16'd10789;
      19846:data<=-16'd10351;
      19847:data<=-16'd10267;
      19848:data<=-16'd9544;
      19849:data<=-16'd9633;
      19850:data<=-16'd9397;
      19851:data<=-16'd7802;
      19852:data<=-16'd7459;
      19853:data<=-16'd7201;
      19854:data<=-16'd6076;
      19855:data<=-16'd6546;
      19856:data<=-16'd7818;
      19857:data<=-16'd8228;
      19858:data<=-16'd7627;
      19859:data<=-16'd6526;
      19860:data<=-16'd5503;
      19861:data<=-16'd4473;
      19862:data<=-16'd4990;
      19863:data<=-16'd5597;
      19864:data<=-16'd4294;
      19865:data<=-16'd4272;
      19866:data<=-16'd3539;
      19867:data<=-16'd2543;
      19868:data<=-16'd5833;
      19869:data<=-16'd2698;
      19870:data<=16'd7203;
      19871:data<=16'd6677;
      19872:data<=16'd2080;
      19873:data<=16'd3997;
      19874:data<=16'd4288;
      19875:data<=16'd3530;
      19876:data<=16'd4438;
      19877:data<=16'd3303;
      19878:data<=16'd3109;
      19879:data<=16'd3709;
      19880:data<=16'd2810;
      19881:data<=16'd2335;
      19882:data<=16'd1280;
      19883:data<=16'd896;
      19884:data<=16'd1926;
      19885:data<=16'd1157;
      19886:data<=16'd784;
      19887:data<=16'd1606;
      19888:data<=16'd1162;
      19889:data<=16'd1343;
      19890:data<=16'd1751;
      19891:data<=16'd1183;
      19892:data<=16'd1507;
      19893:data<=16'd1280;
      19894:data<=-16'd341;
      19895:data<=-16'd817;
      19896:data<=-16'd340;
      19897:data<=-16'd381;
      19898:data<=-16'd244;
      19899:data<=16'd625;
      19900:data<=16'd1108;
      19901:data<=16'd682;
      19902:data<=16'd170;
      19903:data<=16'd261;
      19904:data<=16'd828;
      19905:data<=-16'd8;
      19906:data<=-16'd2224;
      19907:data<=-16'd2409;
      19908:data<=-16'd1310;
      19909:data<=-16'd1613;
      19910:data<=-16'd2079;
      19911:data<=-16'd2070;
      19912:data<=-16'd1594;
      19913:data<=-16'd869;
      19914:data<=-16'd1090;
      19915:data<=-16'd1198;
      19916:data<=-16'd1189;
      19917:data<=-16'd506;
      19918:data<=16'd1224;
      19919:data<=-16'd4240;
      19920:data<=-16'd16495;
      19921:data<=-16'd21185;
      19922:data<=-16'd18565;
      19923:data<=-16'd17614;
      19924:data<=-16'd16668;
      19925:data<=-16'd15004;
      19926:data<=-16'd14719;
      19927:data<=-16'd14320;
      19928:data<=-16'd12794;
      19929:data<=-16'd10810;
      19930:data<=-16'd10869;
      19931:data<=-16'd12522;
      19932:data<=-16'd12113;
      19933:data<=-16'd11126;
      19934:data<=-16'd10957;
      19935:data<=-16'd10295;
      19936:data<=-16'd9451;
      19937:data<=-16'd5800;
      19938:data<=-16'd155;
      19939:data<=16'd1111;
      19940:data<=16'd0;
      19941:data<=16'd961;
      19942:data<=16'd1550;
      19943:data<=16'd1130;
      19944:data<=16'd1707;
      19945:data<=16'd2593;
      19946:data<=16'd2405;
      19947:data<=16'd2056;
      19948:data<=16'd2613;
      19949:data<=16'd2635;
      19950:data<=16'd2328;
      19951:data<=16'd3136;
      19952:data<=16'd3519;
      19953:data<=16'd3369;
      19954:data<=16'd3748;
      19955:data<=16'd4199;
      19956:data<=16'd5332;
      19957:data<=16'd6091;
      19958:data<=16'd5427;
      19959:data<=16'd5518;
      19960:data<=16'd6467;
      19961:data<=16'd7147;
      19962:data<=16'd7192;
      19963:data<=16'd6300;
      19964:data<=16'd5891;
      19965:data<=16'd6291;
      19966:data<=16'd7034;
      19967:data<=16'd6705;
      19968:data<=16'd4640;
      19969:data<=16'd9203;
      19970:data<=16'd21200;
      19971:data<=16'd26166;
      19972:data<=16'd24080;
      19973:data<=16'd24160;
      19974:data<=16'd23588;
      19975:data<=16'd21966;
      19976:data<=16'd21560;
      19977:data<=16'd20037;
      19978:data<=16'd18713;
      19979:data<=16'd18146;
      19980:data<=16'd17655;
      19981:data<=16'd18525;
      19982:data<=16'd18938;
      19983:data<=16'd18545;
      19984:data<=16'd18459;
      19985:data<=16'd17676;
      19986:data<=16'd16844;
      19987:data<=16'd15854;
      19988:data<=16'd14695;
      19989:data<=16'd14402;
      19990:data<=16'd13869;
      19991:data<=16'd13544;
      19992:data<=16'd13218;
      19993:data<=16'd12360;
      19994:data<=16'd13224;
      19995:data<=16'd13379;
      19996:data<=16'd11825;
      19997:data<=16'd11999;
      19998:data<=16'd11790;
      19999:data<=16'd11244;
      20000:data<=16'd11483;
      20001:data<=16'd9404;
      20002:data<=16'd8513;
      20003:data<=16'd8939;
      20004:data<=16'd4532;
      20005:data<=-16'd162;
      20006:data<=-16'd591;
      20007:data<=16'd187;
      20008:data<=16'd1233;
      20009:data<=16'd1530;
      20010:data<=16'd672;
      20011:data<=16'd96;
      20012:data<=16'd29;
      20013:data<=16'd625;
      20014:data<=16'd535;
      20015:data<=-16'd321;
      20016:data<=-16'd908;
      20017:data<=-16'd1334;
      20018:data<=16'd911;
      20019:data<=16'd873;
      20020:data<=-16'd8598;
      20021:data<=-16'd16421;
      20022:data<=-16'd15185;
      20023:data<=-16'd14125;
      20024:data<=-16'd14469;
      20025:data<=-16'd13500;
      20026:data<=-16'd13714;
      20027:data<=-16'd13147;
      20028:data<=-16'd11350;
      20029:data<=-16'd11100;
      20030:data<=-16'd11101;
      20031:data<=-16'd10053;
      20032:data<=-16'd8348;
      20033:data<=-16'd6993;
      20034:data<=-16'd7048;
      20035:data<=-16'd7207;
      20036:data<=-16'd6583;
      20037:data<=-16'd5874;
      20038:data<=-16'd5388;
      20039:data<=-16'd5215;
      20040:data<=-16'd4998;
      20041:data<=-16'd5024;
      20042:data<=-16'd5065;
      20043:data<=-16'd3339;
      20044:data<=-16'd1005;
      20045:data<=-16'd461;
      20046:data<=-16'd681;
      20047:data<=-16'd497;
      20048:data<=-16'd757;
      20049:data<=-16'd1730;
      20050:data<=-16'd1770;
      20051:data<=-16'd500;
      20052:data<=-16'd100;
      20053:data<=-16'd214;
      20054:data<=16'd133;
      20055:data<=-16'd26;
      20056:data<=16'd1243;
      20057:data<=16'd3365;
      20058:data<=16'd2693;
      20059:data<=16'd2129;
      20060:data<=16'd3057;
      20061:data<=16'd2611;
      20062:data<=16'd2751;
      20063:data<=16'd3348;
      20064:data<=16'd2528;
      20065:data<=16'd2340;
      20066:data<=16'd2258;
      20067:data<=16'd2293;
      20068:data<=16'd2889;
      20069:data<=16'd3812;
      20070:data<=16'd12345;
      20071:data<=16'd26116;
      20072:data<=16'd30095;
      20073:data<=16'd26946;
      20074:data<=16'd26606;
      20075:data<=16'd26242;
      20076:data<=16'd24856;
      20077:data<=16'd23807;
      20078:data<=16'd22121;
      20079:data<=16'd21109;
      20080:data<=16'd20427;
      20081:data<=16'd20398;
      20082:data<=16'd21352;
      20083:data<=16'd20404;
      20084:data<=16'd19238;
      20085:data<=16'd19291;
      20086:data<=16'd18039;
      20087:data<=16'd16848;
      20088:data<=16'd16070;
      20089:data<=16'd14358;
      20090:data<=16'd13788;
      20091:data<=16'd14063;
      20092:data<=16'd13186;
      20093:data<=16'd12141;
      20094:data<=16'd12413;
      20095:data<=16'd13182;
      20096:data<=16'd12411;
      20097:data<=16'd11130;
      20098:data<=16'd10965;
      20099:data<=16'd10749;
      20100:data<=16'd10251;
      20101:data<=16'd9168;
      20102:data<=16'd7732;
      20103:data<=16'd7483;
      20104:data<=16'd6595;
      20105:data<=16'd5093;
      20106:data<=16'd5797;
      20107:data<=16'd6922;
      20108:data<=16'd6670;
      20109:data<=16'd6035;
      20110:data<=16'd5579;
      20111:data<=16'd5002;
      20112:data<=16'd3917;
      20113:data<=16'd3959;
      20114:data<=16'd4097;
      20115:data<=16'd2779;
      20116:data<=16'd3213;
      20117:data<=16'd2942;
      20118:data<=16'd1886;
      20119:data<=16'd4827;
      20120:data<=16'd576;
      20121:data<=-16'd12345;
      20122:data<=-16'd15256;
      20123:data<=-16'd12079;
      20124:data<=-16'd13449;
      20125:data<=-16'd12872;
      20126:data<=-16'd12257;
      20127:data<=-16'd13215;
      20128:data<=-16'd10806;
      20129:data<=-16'd10208;
      20130:data<=-16'd11650;
      20131:data<=-16'd10285;
      20132:data<=-16'd8948;
      20133:data<=-16'd8056;
      20134:data<=-16'd7800;
      20135:data<=-16'd8859;
      20136:data<=-16'd7890;
      20137:data<=-16'd8182;
      20138:data<=-16'd12954;
      20139:data<=-16'd15875;
      20140:data<=-16'd15010;
      20141:data<=-16'd14762;
      20142:data<=-16'd15038;
      20143:data<=-16'd14037;
      20144:data<=-16'd13556;
      20145:data<=-16'd13837;
      20146:data<=-16'd12813;
      20147:data<=-16'd11950;
      20148:data<=-16'd12064;
      20149:data<=-16'd11659;
      20150:data<=-16'd11914;
      20151:data<=-16'd12098;
      20152:data<=-16'd10866;
      20153:data<=-16'd10448;
      20154:data<=-16'd10220;
      20155:data<=-16'd9285;
      20156:data<=-16'd9770;
      20157:data<=-16'd10939;
      20158:data<=-16'd10806;
      20159:data<=-16'd9972;
      20160:data<=-16'd10029;
      20161:data<=-16'd9762;
      20162:data<=-16'd8003;
      20163:data<=-16'd8026;
      20164:data<=-16'd8511;
      20165:data<=-16'd7286;
      20166:data<=-16'd8304;
      20167:data<=-16'd7993;
      20168:data<=-16'd6552;
      20169:data<=-16'd10431;
      20170:data<=-16'd6728;
      20171:data<=16'd7175;
      20172:data<=16'd10587;
      20173:data<=16'd6781;
      20174:data<=16'd7841;
      20175:data<=16'd7310;
      20176:data<=16'd5962;
      20177:data<=16'd7094;
      20178:data<=16'd6369;
      20179:data<=16'd5172;
      20180:data<=16'd4643;
      20181:data<=16'd3542;
      20182:data<=16'd2523;
      20183:data<=16'd1454;
      20184:data<=16'd1659;
      20185:data<=16'd2367;
      20186:data<=16'd1888;
      20187:data<=16'd1930;
      20188:data<=16'd1565;
      20189:data<=16'd607;
      20190:data<=16'd972;
      20191:data<=16'd970;
      20192:data<=16'd388;
      20193:data<=16'd30;
      20194:data<=-16'd1086;
      20195:data<=-16'd2067;
      20196:data<=-16'd2208;
      20197:data<=-16'd2008;
      20198:data<=-16'd1971;
      20199:data<=-16'd1985;
      20200:data<=-16'd1322;
      20201:data<=-16'd1193;
      20202:data<=-16'd1753;
      20203:data<=-16'd2182;
      20204:data<=-16'd1709;
      20205:data<=16'd2381;
      20206:data<=16'd5627;
      20207:data<=16'd3369;
      20208:data<=16'd2425;
      20209:data<=16'd3488;
      20210:data<=16'd2514;
      20211:data<=16'd2296;
      20212:data<=16'd1738;
      20213:data<=16'd722;
      20214:data<=16'd1219;
      20215:data<=16'd933;
      20216:data<=16'd1539;
      20217:data<=16'd1481;
      20218:data<=-16'd85;
      20219:data<=16'd1633;
      20220:data<=-16'd3325;
      20221:data<=-16'd16537;
      20222:data<=-16'd20113;
      20223:data<=-16'd17467;
      20224:data<=-16'd18002;
      20225:data<=-16'd16427;
      20226:data<=-16'd15390;
      20227:data<=-16'd15979;
      20228:data<=-16'd14525;
      20229:data<=-16'd14119;
      20230:data<=-16'd13693;
      20231:data<=-16'd13435;
      20232:data<=-16'd15153;
      20233:data<=-16'd14465;
      20234:data<=-16'd13380;
      20235:data<=-16'd14028;
      20236:data<=-16'd12939;
      20237:data<=-16'd12234;
      20238:data<=-16'd12237;
      20239:data<=-16'd10906;
      20240:data<=-16'd10258;
      20241:data<=-16'd10348;
      20242:data<=-16'd10228;
      20243:data<=-16'd9552;
      20244:data<=-16'd9354;
      20245:data<=-16'd11072;
      20246:data<=-16'd11088;
      20247:data<=-16'd9373;
      20248:data<=-16'd9608;
      20249:data<=-16'd9549;
      20250:data<=-16'd8921;
      20251:data<=-16'd9185;
      20252:data<=-16'd8537;
      20253:data<=-16'd7576;
      20254:data<=-16'd6755;
      20255:data<=-16'd6320;
      20256:data<=-16'd7295;
      20257:data<=-16'd7961;
      20258:data<=-16'd8047;
      20259:data<=-16'd7961;
      20260:data<=-16'd7511;
      20261:data<=-16'd7138;
      20262:data<=-16'd5583;
      20263:data<=-16'd4798;
      20264:data<=-16'd5357;
      20265:data<=-16'd4381;
      20266:data<=-16'd4790;
      20267:data<=-16'd4636;
      20268:data<=-16'd2722;
      20269:data<=-16'd5521;
      20270:data<=-16'd2874;
      20271:data<=16'd8343;
      20272:data<=16'd8699;
      20273:data<=16'd2930;
      20274:data<=16'd4246;
      20275:data<=16'd4205;
      20276:data<=16'd2660;
      20277:data<=16'd3491;
      20278:data<=16'd2896;
      20279:data<=16'd2964;
      20280:data<=16'd3107;
      20281:data<=16'd2014;
      20282:data<=16'd1971;
      20283:data<=16'd643;
      20284:data<=-16'd334;
      20285:data<=16'd848;
      20286:data<=16'd614;
      20287:data<=16'd235;
      20288:data<=16'd737;
      20289:data<=16'd1328;
      20290:data<=16'd2482;
      20291:data<=16'd2469;
      20292:data<=16'd2522;
      20293:data<=16'd3095;
      20294:data<=16'd1888;
      20295:data<=16'd1063;
      20296:data<=16'd795;
      20297:data<=16'd405;
      20298:data<=16'd1337;
      20299:data<=16'd1309;
      20300:data<=16'd919;
      20301:data<=16'd1726;
      20302:data<=16'd1419;
      20303:data<=16'd1143;
      20304:data<=16'd1418;
      20305:data<=16'd1213;
      20306:data<=16'd1095;
      20307:data<=-16'd50;
      20308:data<=-16'd705;
      20309:data<=-16'd133;
      20310:data<=-16'd566;
      20311:data<=-16'd472;
      20312:data<=-16'd240;
      20313:data<=-16'd760;
      20314:data<=-16'd749;
      20315:data<=-16'd1322;
      20316:data<=-16'd676;
      20317:data<=16'd50;
      20318:data<=-16'd1181;
      20319:data<=16'd149;
      20320:data<=-16'd3336;
      20321:data<=-16'd15600;
      20322:data<=-16'd20588;
      20323:data<=-16'd17949;
      20324:data<=-16'd17793;
      20325:data<=-16'd16757;
      20326:data<=-16'd15054;
      20327:data<=-16'd14411;
      20328:data<=-16'd13380;
      20329:data<=-16'd13515;
      20330:data<=-16'd12351;
      20331:data<=-16'd11330;
      20332:data<=-16'd13247;
      20333:data<=-16'd12759;
      20334:data<=-16'd11133;
      20335:data<=-16'd11245;
      20336:data<=-16'd10477;
      20337:data<=-16'd10360;
      20338:data<=-16'd8610;
      20339:data<=-16'd3312;
      20340:data<=-16'd801;
      20341:data<=-16'd1303;
      20342:data<=-16'd1149;
      20343:data<=-16'd735;
      20344:data<=-16'd281;
      20345:data<=-16'd109;
      20346:data<=16'd246;
      20347:data<=16'd649;
      20348:data<=16'd56;
      20349:data<=16'd194;
      20350:data<=16'd933;
      20351:data<=16'd1048;
      20352:data<=16'd1477;
      20353:data<=16'd1747;
      20354:data<=16'd1956;
      20355:data<=16'd2352;
      20356:data<=16'd2381;
      20357:data<=16'd3233;
      20358:data<=16'd4308;
      20359:data<=16'd4605;
      20360:data<=16'd4696;
      20361:data<=16'd4187;
      20362:data<=16'd4149;
      20363:data<=16'd4758;
      20364:data<=16'd5046;
      20365:data<=16'd5850;
      20366:data<=16'd5792;
      20367:data<=16'd5394;
      20368:data<=16'd5935;
      20369:data<=16'd5063;
      20370:data<=16'd8451;
      20371:data<=16'd19206;
      20372:data<=16'd25226;
      20373:data<=16'd23472;
      20374:data<=16'd22042;
      20375:data<=16'd21476;
      20376:data<=16'd20716;
      20377:data<=16'd20122;
      20378:data<=16'd19094;
      20379:data<=16'd18635;
      20380:data<=16'd17901;
      20381:data<=16'd17428;
      20382:data<=16'd18903;
      20383:data<=16'd19082;
      20384:data<=16'd17617;
      20385:data<=16'd17262;
      20386:data<=16'd16627;
      20387:data<=16'd15600;
      20388:data<=16'd15211;
      20389:data<=16'd14355;
      20390:data<=16'd13505;
      20391:data<=16'd13218;
      20392:data<=16'd12944;
      20393:data<=16'd12536;
      20394:data<=16'd12176;
      20395:data<=16'd12886;
      20396:data<=16'd13500;
      20397:data<=16'd12483;
      20398:data<=16'd12082;
      20399:data<=16'd12037;
      20400:data<=16'd10839;
      20401:data<=16'd10721;
      20402:data<=16'd10639;
      20403:data<=16'd9207;
      20404:data<=16'd9091;
      20405:data<=16'd7920;
      20406:data<=16'd3621;
      20407:data<=16'd2030;
      20408:data<=16'd3891;
      20409:data<=16'd3623;
      20410:data<=16'd2400;
      20411:data<=16'd3148;
      20412:data<=16'd3127;
      20413:data<=16'd2270;
      20414:data<=16'd2557;
      20415:data<=16'd1895;
      20416:data<=16'd1034;
      20417:data<=16'd1398;
      20418:data<=16'd710;
      20419:data<=16'd1580;
      20420:data<=16'd2205;
      20421:data<=-16'd5747;
      20422:data<=-16'd14548;
      20423:data<=-16'd14325;
      20424:data<=-16'd12860;
      20425:data<=-16'd13577;
      20426:data<=-16'd12401;
      20427:data<=-16'd11505;
      20428:data<=-16'd11576;
      20429:data<=-16'd11003;
      20430:data<=-16'd10313;
      20431:data<=-16'd9649;
      20432:data<=-16'd9151;
      20433:data<=-16'd7900;
      20434:data<=-16'd6379;
      20435:data<=-16'd6316;
      20436:data<=-16'd5899;
      20437:data<=-16'd5268;
      20438:data<=-16'd5695;
      20439:data<=-16'd5180;
      20440:data<=-16'd4410;
      20441:data<=-16'd4262;
      20442:data<=-16'd3877;
      20443:data<=-16'd4256;
      20444:data<=-16'd3941;
      20445:data<=-16'd1971;
      20446:data<=-16'd735;
      20447:data<=-16'd444;
      20448:data<=-16'd940;
      20449:data<=-16'd1551;
      20450:data<=-16'd820;
      20451:data<=-16'd502;
      20452:data<=-16'd1030;
      20453:data<=-16'd923;
      20454:data<=-16'd657;
      20455:data<=-16'd411;
      20456:data<=-16'd203;
      20457:data<=16'd302;
      20458:data<=16'd1260;
      20459:data<=16'd1633;
      20460:data<=16'd2165;
      20461:data<=16'd2466;
      20462:data<=16'd1686;
      20463:data<=16'd1801;
      20464:data<=16'd2090;
      20465:data<=16'd2182;
      20466:data<=16'd2931;
      20467:data<=16'd2159;
      20468:data<=16'd2093;
      20469:data<=16'd3210;
      20470:data<=16'd2711;
      20471:data<=16'd8549;
      20472:data<=16'd20980;
      20473:data<=16'd26398;
      20474:data<=16'd25461;
      20475:data<=16'd24861;
      20476:data<=16'd23044;
      20477:data<=16'd21729;
      20478:data<=16'd21933;
      20479:data<=16'd21217;
      20480:data<=16'd19984;
      20481:data<=16'd18691;
      20482:data<=16'd18418;
      20483:data<=16'd19127;
      20484:data<=16'd18604;
      20485:data<=16'd17740;
      20486:data<=16'd16967;
      20487:data<=16'd15690;
      20488:data<=16'd15126;
      20489:data<=16'd14390;
      20490:data<=16'd12950;
      20491:data<=16'd12041;
      20492:data<=16'd11400;
      20493:data<=16'd11013;
      20494:data<=16'd10880;
      20495:data<=16'd10836;
      20496:data<=16'd10878;
      20497:data<=16'd10176;
      20498:data<=16'd9615;
      20499:data<=16'd9682;
      20500:data<=16'd9115;
      20501:data<=16'd8511;
      20502:data<=16'd7884;
      20503:data<=16'd6953;
      20504:data<=16'd6643;
      20505:data<=16'd6068;
      20506:data<=16'd5295;
      20507:data<=16'd5650;
      20508:data<=16'd6639;
      20509:data<=16'd6896;
      20510:data<=16'd5702;
      20511:data<=16'd5204;
      20512:data<=16'd5562;
      20513:data<=16'd4099;
      20514:data<=16'd3230;
      20515:data<=16'd3339;
      20516:data<=16'd2725;
      20517:data<=16'd3788;
      20518:data<=16'd2758;
      20519:data<=16'd628;
      20520:data<=16'd3815;
      20521:data<=16'd312;
      20522:data<=-16'd12471;
      20523:data<=-16'd15995;
      20524:data<=-16'd12904;
      20525:data<=-16'd13661;
      20526:data<=-16'd13126;
      20527:data<=-16'd12298;
      20528:data<=-16'd13286;
      20529:data<=-16'd12173;
      20530:data<=-16'd11311;
      20531:data<=-16'd11752;
      20532:data<=-16'd10956;
      20533:data<=-16'd9380;
      20534:data<=-16'd7853;
      20535:data<=-16'd7755;
      20536:data<=-16'd8822;
      20537:data<=-16'd8355;
      20538:data<=-16'd7031;
      20539:data<=-16'd8156;
      20540:data<=-16'd11552;
      20541:data<=-16'd12938;
      20542:data<=-16'd12204;
      20543:data<=-16'd12610;
      20544:data<=-16'd12354;
      20545:data<=-16'd11145;
      20546:data<=-16'd11189;
      20547:data<=-16'd10842;
      20548:data<=-16'd10781;
      20549:data<=-16'd11371;
      20550:data<=-16'd10458;
      20551:data<=-16'd10044;
      20552:data<=-16'd9944;
      20553:data<=-16'd8636;
      20554:data<=-16'd8523;
      20555:data<=-16'd8875;
      20556:data<=-16'd8614;
      20557:data<=-16'd9101;
      20558:data<=-16'd9909;
      20559:data<=-16'd10273;
      20560:data<=-16'd9530;
      20561:data<=-16'd9303;
      20562:data<=-16'd9823;
      20563:data<=-16'd8093;
      20564:data<=-16'd7277;
      20565:data<=-16'd7774;
      20566:data<=-16'd6208;
      20567:data<=-16'd6889;
      20568:data<=-16'd7074;
      20569:data<=-16'd4880;
      20570:data<=-16'd7752;
      20571:data<=-16'd5062;
      20572:data<=16'd7844;
      20573:data<=16'd11709;
      20574:data<=16'd8332;
      20575:data<=16'd9295;
      20576:data<=16'd8584;
      20577:data<=16'd6778;
      20578:data<=16'd7407;
      20579:data<=16'd7124;
      20580:data<=16'd6940;
      20581:data<=16'd6563;
      20582:data<=16'd5090;
      20583:data<=16'd3896;
      20584:data<=16'd2431;
      20585:data<=16'd2441;
      20586:data<=16'd3178;
      20587:data<=16'd2114;
      20588:data<=16'd1895;
      20589:data<=16'd2109;
      20590:data<=16'd1318;
      20591:data<=16'd1312;
      20592:data<=16'd1084;
      20593:data<=16'd855;
      20594:data<=16'd1403;
      20595:data<=16'd499;
      20596:data<=-16'd1428;
      20597:data<=-16'd2305;
      20598:data<=-16'd1666;
      20599:data<=-16'd948;
      20600:data<=-16'd1225;
      20601:data<=-16'd1005;
      20602:data<=-16'd943;
      20603:data<=-16'd1419;
      20604:data<=-16'd1080;
      20605:data<=-16'd1419;
      20606:data<=-16'd115;
      20607:data<=16'd3973;
      20608:data<=16'd4704;
      20609:data<=16'd2786;
      20610:data<=16'd2290;
      20611:data<=16'd2490;
      20612:data<=16'd3218;
      20613:data<=16'd2787;
      20614:data<=16'd1765;
      20615:data<=16'd1997;
      20616:data<=16'd1410;
      20617:data<=16'd1771;
      20618:data<=16'd2046;
      20619:data<=16'd402;
      20620:data<=16'd1301;
      20621:data<=-16'd3207;
      20622:data<=-16'd15891;
      20623:data<=-16'd19948;
      20624:data<=-16'd16921;
      20625:data<=-16'd17101;
      20626:data<=-16'd15893;
      20627:data<=-16'd14684;
      20628:data<=-16'd15343;
      20629:data<=-16'd14413;
      20630:data<=-16'd14143;
      20631:data<=-16'd13474;
      20632:data<=-16'd12587;
      20633:data<=-16'd14069;
      20634:data<=-16'd13762;
      20635:data<=-16'd12627;
      20636:data<=-16'd12991;
      20637:data<=-16'd11808;
      20638:data<=-16'd10960;
      20639:data<=-16'd11101;
      20640:data<=-16'd10143;
      20641:data<=-16'd9303;
      20642:data<=-16'd8508;
      20643:data<=-16'd7990;
      20644:data<=-16'd7962;
      20645:data<=-16'd8066;
      20646:data<=-16'd9183;
      20647:data<=-16'd9150;
      20648:data<=-16'd8235;
      20649:data<=-16'd8731;
      20650:data<=-16'd8288;
      20651:data<=-16'd7767;
      20652:data<=-16'd8134;
      20653:data<=-16'd7087;
      20654:data<=-16'd6520;
      20655:data<=-16'd6583;
      20656:data<=-16'd6166;
      20657:data<=-16'd6968;
      20658:data<=-16'd7743;
      20659:data<=-16'd7650;
      20660:data<=-16'd7230;
      20661:data<=-16'd7039;
      20662:data<=-16'd7727;
      20663:data<=-16'd6534;
      20664:data<=-16'd5159;
      20665:data<=-16'd5890;
      20666:data<=-16'd4811;
      20667:data<=-16'd4578;
      20668:data<=-16'd5086;
      20669:data<=-16'd2869;
      20670:data<=-16'd4772;
      20671:data<=-16'd3777;
      20672:data<=16'd8472;
      20673:data<=16'd13217;
      20674:data<=16'd6740;
      20675:data<=16'd5098;
      20676:data<=16'd5806;
      20677:data<=16'd4723;
      20678:data<=16'd5250;
      20679:data<=16'd5027;
      20680:data<=16'd4244;
      20681:data<=16'd4394;
      20682:data<=16'd4087;
      20683:data<=16'd3092;
      20684:data<=16'd1610;
      20685:data<=16'd1609;
      20686:data<=16'd2504;
      20687:data<=16'd1600;
      20688:data<=16'd1321;
      20689:data<=16'd2203;
      20690:data<=16'd2065;
      20691:data<=16'd1783;
      20692:data<=16'd1266;
      20693:data<=16'd1104;
      20694:data<=16'd2049;
      20695:data<=16'd1495;
      20696:data<=-16'd127;
      20697:data<=-16'd417;
      20698:data<=-16'd147;
      20699:data<=16'd68;
      20700:data<=16'd376;
      20701:data<=16'd450;
      20702:data<=16'd243;
      20703:data<=16'd82;
      20704:data<=16'd64;
      20705:data<=-16'd188;
      20706:data<=16'd256;
      20707:data<=16'd1225;
      20708:data<=16'd440;
      20709:data<=-16'd890;
      20710:data<=-16'd898;
      20711:data<=-16'd622;
      20712:data<=-16'd203;
      20713:data<=-16'd83;
      20714:data<=-16'd344;
      20715:data<=-16'd328;
      20716:data<=-16'd1095;
      20717:data<=-16'd1219;
      20718:data<=-16'd325;
      20719:data<=-16'd496;
      20720:data<=16'd61;
      20721:data<=-16'd3042;
      20722:data<=-16'd13919;
      20723:data<=-16'd20280;
      20724:data<=-16'd17976;
      20725:data<=-16'd17135;
      20726:data<=-16'd16953;
      20727:data<=-16'd14971;
      20728:data<=-16'd14613;
      20729:data<=-16'd14349;
      20730:data<=-16'd13731;
      20731:data<=-16'd13159;
      20732:data<=-16'd11843;
      20733:data<=-16'd12114;
      20734:data<=-16'd12408;
      20735:data<=-16'd11359;
      20736:data<=-16'd11408;
      20737:data<=-16'd10316;
      20738:data<=-16'd8994;
      20739:data<=-16'd9864;
      20740:data<=-16'd7309;
      20741:data<=-16'd1956;
      20742:data<=-16'd358;
      20743:data<=-16'd779;
      20744:data<=-16'd408;
      20745:data<=-16'd64;
      20746:data<=16'd337;
      20747:data<=16'd785;
      20748:data<=16'd955;
      20749:data<=16'd795;
      20750:data<=16'd746;
      20751:data<=16'd1104;
      20752:data<=16'd1204;
      20753:data<=16'd1136;
      20754:data<=16'd1321;
      20755:data<=16'd1641;
      20756:data<=16'd1606;
      20757:data<=16'd1160;
      20758:data<=16'd2147;
      20759:data<=16'd3959;
      20760:data<=16'd3914;
      20761:data<=16'd3321;
      20762:data<=16'd3360;
      20763:data<=16'd3334;
      20764:data<=16'd3471;
      20765:data<=16'd3542;
      20766:data<=16'd4264;
      20767:data<=16'd4810;
      20768:data<=16'd4090;
      20769:data<=16'd4484;
      20770:data<=16'd4376;
      20771:data<=16'd5909;
      20772:data<=16'd15843;
      20773:data<=16'd24283;
      20774:data<=16'd22909;
      20775:data<=16'd21563;
      20776:data<=16'd21867;
      20777:data<=16'd20439;
      20778:data<=16'd20394;
      20779:data<=16'd19556;
      20780:data<=16'd18017;
      20781:data<=16'd18219;
      20782:data<=16'd17230;
      20783:data<=16'd16936;
      20784:data<=16'd18031;
      20785:data<=16'd17000;
      20786:data<=16'd16446;
      20787:data<=16'd16678;
      20788:data<=16'd15620;
      20789:data<=16'd15176;
      20790:data<=16'd14228;
      20791:data<=16'd12643;
      20792:data<=16'd12657;
      20793:data<=16'd12401;
      20794:data<=16'd11509;
      20795:data<=16'd11442;
      20796:data<=16'd11674;
      20797:data<=16'd11852;
      20798:data<=16'd11253;
      20799:data<=16'd10806;
      20800:data<=16'd11621;
      20801:data<=16'd11163;
      20802:data<=16'd9744;
      20803:data<=16'd9555;
      20804:data<=16'd8798;
      20805:data<=16'd8176;
      20806:data<=16'd9300;
      20807:data<=16'd7680;
      20808:data<=16'd3159;
      20809:data<=16'd2362;
      20810:data<=16'd3847;
      20811:data<=16'd3148;
      20812:data<=16'd3307;
      20813:data<=16'd3921;
      20814:data<=16'd2717;
      20815:data<=16'd2840;
      20816:data<=16'd2638;
      20817:data<=16'd1478;
      20818:data<=16'd2713;
      20819:data<=16'd2074;
      20820:data<=16'd1313;
      20821:data<=16'd3805;
      20822:data<=-16'd2055;
      20823:data<=-16'd13259;
      20824:data<=-16'd14556;
      20825:data<=-16'd12537;
      20826:data<=-16'd13388;
      20827:data<=-16'd11759;
      20828:data<=-16'd10974;
      20829:data<=-16'd11784;
      20830:data<=-16'd10599;
      20831:data<=-16'd10138;
      20832:data<=-16'd10334;
      20833:data<=-16'd9192;
      20834:data<=-16'd7511;
      20835:data<=-16'd6341;
      20836:data<=-16'd6743;
      20837:data<=-16'd6749;
      20838:data<=-16'd5859;
      20839:data<=-16'd6050;
      20840:data<=-16'd5178;
      20841:data<=-16'd3805;
      20842:data<=-16'd4376;
      20843:data<=-16'd4667;
      20844:data<=-16'd4681;
      20845:data<=-16'd4485;
      20846:data<=-16'd2408;
      20847:data<=-16'd931;
      20848:data<=-16'd842;
      20849:data<=-16'd652;
      20850:data<=-16'd1198;
      20851:data<=-16'd1660;
      20852:data<=-16'd1043;
      20853:data<=-16'd726;
      20854:data<=-16'd955;
      20855:data<=-16'd770;
      20856:data<=-16'd875;
      20857:data<=-16'd1751;
      20858:data<=-16'd682;
      20859:data<=16'd1530;
      20860:data<=16'd1055;
      20861:data<=16'd412;
      20862:data<=16'd849;
      20863:data<=16'd285;
      20864:data<=16'd625;
      20865:data<=16'd872;
      20866:data<=16'd375;
      20867:data<=16'd923;
      20868:data<=16'd135;
      20869:data<=16'd355;
      20870:data<=16'd1595;
      20871:data<=-16'd11;
      20872:data<=16'd5353;
      20873:data<=16'd17484;
      20874:data<=16'd21852;
      20875:data<=16'd22573;
      20876:data<=16'd24474;
      20877:data<=16'd22526;
      20878:data<=16'd21061;
      20879:data<=16'd20873;
      20880:data<=16'd19215;
      20881:data<=16'd18968;
      20882:data<=16'd18580;
      20883:data<=16'd18060;
      20884:data<=16'd18595;
      20885:data<=16'd17440;
      20886:data<=16'd16540;
      20887:data<=16'd16164;
      20888:data<=16'd14531;
      20889:data<=16'd13923;
      20890:data<=16'd13095;
      20891:data<=16'd11724;
      20892:data<=16'd11753;
      20893:data<=16'd11094;
      20894:data<=16'd10029;
      20895:data<=16'd9944;
      20896:data<=16'd10225;
      20897:data<=16'd10480;
      20898:data<=16'd9265;
      20899:data<=16'd8276;
      20900:data<=16'd8866;
      20901:data<=16'd8385;
      20902:data<=16'd7884;
      20903:data<=16'd7964;
      20904:data<=16'd7015;
      20905:data<=16'd6504;
      20906:data<=16'd6469;
      20907:data<=16'd6237;
      20908:data<=16'd6102;
      20909:data<=16'd5988;
      20910:data<=16'd6660;
      20911:data<=16'd6672;
      20912:data<=16'd5745;
      20913:data<=16'd5275;
      20914:data<=16'd4162;
      20915:data<=16'd4073;
      20916:data<=16'd4190;
      20917:data<=16'd2643;
      20918:data<=16'd3703;
      20919:data<=16'd3779;
      20920:data<=16'd1754;
      20921:data<=16'd4535;
      20922:data<=16'd1149;
      20923:data<=-16'd11771;
      20924:data<=-16'd15596;
      20925:data<=-16'd12590;
      20926:data<=-16'd13618;
      20927:data<=-16'd13361;
      20928:data<=-16'd12188;
      20929:data<=-16'd12656;
      20930:data<=-16'd11646;
      20931:data<=-16'd11060;
      20932:data<=-16'd11776;
      20933:data<=-16'd11291;
      20934:data<=-16'd9618;
      20935:data<=-16'd8707;
      20936:data<=-16'd9242;
      20937:data<=-16'd8900;
      20938:data<=-16'd8190;
      20939:data<=-16'd8261;
      20940:data<=-16'd7301;
      20941:data<=-16'd8551;
      20942:data<=-16'd12730;
      20943:data<=-16'd14114;
      20944:data<=-16'd13574;
      20945:data<=-16'd13273;
      20946:data<=-16'd12034;
      20947:data<=-16'd11274;
      20948:data<=-16'd11053;
      20949:data<=-16'd10954;
      20950:data<=-16'd11353;
      20951:data<=-16'd11094;
      20952:data<=-16'd11050;
      20953:data<=-16'd11173;
      20954:data<=-16'd10187;
      20955:data<=-16'd9612;
      20956:data<=-16'd9492;
      20957:data<=-16'd9271;
      20958:data<=-16'd9781;
      20959:data<=-16'd10707;
      20960:data<=-16'd11356;
      20961:data<=-16'd10774;
      20962:data<=-16'd10110;
      20963:data<=-16'd10448;
      20964:data<=-16'd9718;
      20965:data<=-16'd9420;
      20966:data<=-16'd9899;
      20967:data<=-16'd8705;
      20968:data<=-16'd8724;
      20969:data<=-16'd8536;
      20970:data<=-16'd7371;
      20971:data<=-16'd10131;
      20972:data<=-16'd6990;
      20973:data<=16'd5589;
      20974:data<=16'd9861;
      20975:data<=16'd6749;
      20976:data<=16'd7694;
      20977:data<=16'd7498;
      20978:data<=16'd5934;
      20979:data<=16'd6672;
      20980:data<=16'd6068;
      20981:data<=16'd5435;
      20982:data<=16'd5865;
      20983:data<=16'd4925;
      20984:data<=16'd3704;
      20985:data<=16'd2954;
      20986:data<=16'd2880;
      20987:data<=16'd2734;
      20988:data<=16'd1492;
      20989:data<=16'd1366;
      20990:data<=16'd1629;
      20991:data<=16'd872;
      20992:data<=16'd1105;
      20993:data<=16'd1204;
      20994:data<=16'd658;
      20995:data<=16'd766;
      20996:data<=-16'd199;
      20997:data<=-16'd1565;
      20998:data<=-16'd1477;
      20999:data<=-16'd987;
      21000:data<=-16'd801;
      21001:data<=-16'd1063;
      21002:data<=-16'd1011;
      21003:data<=-16'd550;
      21004:data<=-16'd808;
      21005:data<=-16'd732;
      21006:data<=-16'd861;
      21007:data<=-16'd1668;
      21008:data<=16'd67;
      21009:data<=16'd3008;
      21010:data<=16'd3627;
      21011:data<=16'd3275;
      21012:data<=16'd3089;
      21013:data<=16'd2687;
      21014:data<=16'd2353;
      21015:data<=16'd2534;
      21016:data<=16'd2728;
      21017:data<=16'd2135;
      21018:data<=16'd2164;
      21019:data<=16'd2231;
      21020:data<=16'd1677;
      21021:data<=16'd2560;
      21022:data<=-16'd1363;
      21023:data<=-16'd12091;
      21024:data<=-16'd16612;
      21025:data<=-16'd14522;
      21026:data<=-16'd14709;
      21027:data<=-16'd14178;
      21028:data<=-16'd12800;
      21029:data<=-16'd13244;
      21030:data<=-16'd12618;
      21031:data<=-16'd12195;
      21032:data<=-16'd12521;
      21033:data<=-16'd11952;
      21034:data<=-16'd12057;
      21035:data<=-16'd11885;
      21036:data<=-16'd11317;
      21037:data<=-16'd11323;
      21038:data<=-16'd10044;
      21039:data<=-16'd8945;
      21040:data<=-16'd8959;
      21041:data<=-16'd8153;
      21042:data<=-16'd7800;
      21043:data<=-16'd8269;
      21044:data<=-16'd7864;
      21045:data<=-16'd6673;
      21046:data<=-16'd6367;
      21047:data<=-16'd7918;
      21048:data<=-16'd8789;
      21049:data<=-16'd8062;
      21050:data<=-16'd7796;
      21051:data<=-16'd7451;
      21052:data<=-16'd7315;
      21053:data<=-16'd7420;
      21054:data<=-16'd6349;
      21055:data<=-16'd6179;
      21056:data<=-16'd6622;
      21057:data<=-16'd5853;
      21058:data<=-16'd5853;
      21059:data<=-16'd6284;
      21060:data<=-16'd6443;
      21061:data<=-16'd6833;
      21062:data<=-16'd6326;
      21063:data<=-16'd5946;
      21064:data<=-16'd5764;
      21065:data<=-16'd5121;
      21066:data<=-16'd5254;
      21067:data<=-16'd4801;
      21068:data<=-16'd4290;
      21069:data<=-16'd4297;
      21070:data<=-16'd3259;
      21071:data<=-16'd4739;
      21072:data<=-16'd4423;
      21073:data<=16'd5213;
      21074:data<=16'd12085;
      21075:data<=16'd8141;
      21076:data<=16'd4041;
      21077:data<=16'd3497;
      21078:data<=16'd3118;
      21079:data<=16'd3260;
      21080:data<=16'd3548;
      21081:data<=16'd3428;
      21082:data<=16'd3448;
      21083:data<=16'd3632;
      21084:data<=16'd2784;
      21085:data<=16'd960;
      21086:data<=16'd723;
      21087:data<=16'd1293;
      21088:data<=16'd1115;
      21089:data<=16'd1403;
      21090:data<=16'd1084;
      21091:data<=16'd532;
      21092:data<=16'd1183;
      21093:data<=16'd987;
      21094:data<=16'd813;
      21095:data<=16'd1406;
      21096:data<=16'd209;
      21097:data<=-16'd1124;
      21098:data<=-16'd711;
      21099:data<=-16'd162;
      21100:data<=16'd42;
      21101:data<=16'd315;
      21102:data<=16'd789;
      21103:data<=16'd725;
      21104:data<=16'd337;
      21105:data<=16'd945;
      21106:data<=16'd1063;
      21107:data<=16'd737;
      21108:data<=16'd1343;
      21109:data<=16'd602;
      21110:data<=-16'd647;
      21111:data<=-16'd168;
      21112:data<=-16'd77;
      21113:data<=-16'd171;
      21114:data<=16'd428;
      21115:data<=16'd337;
      21116:data<=16'd344;
      21117:data<=16'd664;
      21118:data<=16'd503;
      21119:data<=16'd127;
      21120:data<=16'd56;
      21121:data<=16'd1243;
      21122:data<=-16'd631;
      21123:data<=-16'd9459;
      21124:data<=-16'd16271;
      21125:data<=-16'd15338;
      21126:data<=-16'd13944;
      21127:data<=-16'd14004;
      21128:data<=-16'd12706;
      21129:data<=-16'd12217;
      21130:data<=-16'd12442;
      21131:data<=-16'd11626;
      21132:data<=-16'd10795;
      21133:data<=-16'd10126;
      21134:data<=-16'd10117;
      21135:data<=-16'd10953;
      21136:data<=-16'd10470;
      21137:data<=-16'd9245;
      21138:data<=-16'd8851;
      21139:data<=-16'd7874;
      21140:data<=-16'd7066;
      21141:data<=-16'd7277;
      21142:data<=-16'd4707;
      21143:data<=16'd68;
      21144:data<=16'd1262;
      21145:data<=16'd273;
      21146:data<=16'd1178;
      21147:data<=16'd1726;
      21148:data<=16'd1398;
      21149:data<=16'd2009;
      21150:data<=16'd1842;
      21151:data<=16'd1287;
      21152:data<=16'd1865;
      21153:data<=16'd2097;
      21154:data<=16'd2050;
      21155:data<=16'd2067;
      21156:data<=16'd1804;
      21157:data<=16'd1906;
      21158:data<=16'd1806;
      21159:data<=16'd2519;
      21160:data<=16'd4322;
      21161:data<=16'd4367;
      21162:data<=16'd3929;
      21163:data<=16'd4282;
      21164:data<=16'd4102;
      21165:data<=16'd4575;
      21166:data<=16'd4651;
      21167:data<=16'd4211;
      21168:data<=16'd4975;
      21169:data<=16'd4611;
      21170:data<=16'd4551;
      21171:data<=16'd5121;
      21172:data<=16'd4927;
      21173:data<=16'd11794;
      21174:data<=16'd21573;
      21175:data<=16'd21804;
      21176:data<=16'd19737;
      21177:data<=16'd20301;
      21178:data<=16'd18897;
      21179:data<=16'd19138;
      21180:data<=16'd19690;
      21181:data<=16'd17854;
      21182:data<=16'd17274;
      21183:data<=16'd16515;
      21184:data<=16'd16386;
      21185:data<=16'd17989;
      21186:data<=16'd17112;
      21187:data<=16'd15729;
      21188:data<=16'd15427;
      21189:data<=16'd14410;
      21190:data<=16'd14331;
      21191:data<=16'd14096;
      21192:data<=16'd13071;
      21193:data<=16'd13035;
      21194:data<=16'd12898;
      21195:data<=16'd12590;
      21196:data<=16'd12422;
      21197:data<=16'd12659;
      21198:data<=16'd13317;
      21199:data<=16'd12107;
      21200:data<=16'd10749;
      21201:data<=16'd11168;
      21202:data<=16'd11153;
      21203:data<=16'd10860;
      21204:data<=16'd10383;
      21205:data<=16'd9969;
      21206:data<=16'd10144;
      21207:data<=16'd9502;
      21208:data<=16'd9741;
      21209:data<=16'd8840;
      21210:data<=16'd4554;
      21211:data<=16'd3497;
      21212:data<=16'd4513;
      21213:data<=16'd3582;
      21214:data<=16'd4387;
      21215:data<=16'd4698;
      21216:data<=16'd4044;
      21217:data<=16'd4482;
      21218:data<=16'd3133;
      21219:data<=16'd3107;
      21220:data<=16'd3435;
      21221:data<=16'd2452;
      21222:data<=16'd5562;
      21223:data<=16'd2173;
      21224:data<=-16'd9867;
      21225:data<=-16'd11794;
      21226:data<=-16'd8784;
      21227:data<=-16'd11030;
      21228:data<=-16'd10187;
      21229:data<=-16'd8722;
      21230:data<=-16'd9988;
      21231:data<=-16'd9295;
      21232:data<=-16'd8840;
      21233:data<=-16'd8637;
      21234:data<=-16'd7225;
      21235:data<=-16'd6266;
      21236:data<=-16'd5410;
      21237:data<=-16'd5688;
      21238:data<=-16'd6041;
      21239:data<=-16'd5046;
      21240:data<=-16'd4883;
      21241:data<=-16'd4599;
      21242:data<=-16'd4211;
      21243:data<=-16'd4454;
      21244:data<=-16'd3698;
      21245:data<=-16'd3770;
      21246:data<=-16'd3800;
      21247:data<=-16'd1877;
      21248:data<=-16'd1391;
      21249:data<=-16'd1639;
      21250:data<=-16'd867;
      21251:data<=-16'd1001;
      21252:data<=-16'd1609;
      21253:data<=-16'd1757;
      21254:data<=-16'd1158;
      21255:data<=-16'd829;
      21256:data<=-16'd1542;
      21257:data<=-16'd1333;
      21258:data<=-16'd1377;
      21259:data<=-16'd1312;
      21260:data<=16'd763;
      21261:data<=16'd770;
      21262:data<=-16'd133;
      21263:data<=16'd573;
      21264:data<=-16'd558;
      21265:data<=-16'd917;
      21266:data<=16'd6;
      21267:data<=-16'd469;
      21268:data<=16'd250;
      21269:data<=-16'd205;
      21270:data<=-16'd855;
      21271:data<=16'd500;
      21272:data<=-16'd1104;
      21273:data<=16'd3498;
      21274:data<=16'd15700;
      21275:data<=16'd17236;
      21276:data<=16'd15261;
      21277:data<=16'd20764;
      21278:data<=16'd21423;
      21279:data<=16'd18632;
      21280:data<=16'd19300;
      21281:data<=16'd18509;
      21282:data<=16'd17214;
      21283:data<=16'd16545;
      21284:data<=16'd15790;
      21285:data<=16'd16407;
      21286:data<=16'd15908;
      21287:data<=16'd14854;
      21288:data<=16'd14463;
      21289:data<=16'd12991;
      21290:data<=16'd12275;
      21291:data<=16'd11662;
      21292:data<=16'd10050;
      21293:data<=16'd9797;
      21294:data<=16'd9893;
      21295:data<=16'd9536;
      21296:data<=16'd8895;
      21297:data<=16'd8264;
      21298:data<=16'd9658;
      21299:data<=16'd10245;
      21300:data<=16'd8423;
      21301:data<=16'd7794;
      21302:data<=16'd7582;
      21303:data<=16'd6839;
      21304:data<=16'd6522;
      21305:data<=16'd5921;
      21306:data<=16'd5965;
      21307:data<=16'd6070;
      21308:data<=16'd5319;
      21309:data<=16'd5539;
      21310:data<=16'd6162;
      21311:data<=16'd5964;
      21312:data<=16'd5224;
      21313:data<=16'd4869;
      21314:data<=16'd5187;
      21315:data<=16'd4464;
      21316:data<=16'd4137;
      21317:data<=16'd4313;
      21318:data<=16'd2740;
      21319:data<=16'd3239;
      21320:data<=16'd3952;
      21321:data<=16'd1912;
      21322:data<=16'd3442;
      21323:data<=16'd1494;
      21324:data<=-16'd9219;
      21325:data<=-16'd13235;
      21326:data<=-16'd10763;
      21327:data<=-16'd11852;
      21328:data<=-16'd11309;
      21329:data<=-16'd10093;
      21330:data<=-16'd11705;
      21331:data<=-16'd11169;
      21332:data<=-16'd10125;
      21333:data<=-16'd10725;
      21334:data<=-16'd10155;
      21335:data<=-16'd8675;
      21336:data<=-16'd7583;
      21337:data<=-16'd7677;
      21338:data<=-16'd7703;
      21339:data<=-16'd6801;
      21340:data<=-16'd7230;
      21341:data<=-16'd7116;
      21342:data<=-16'd5729;
      21343:data<=-16'd7826;
      21344:data<=-16'd11809;
      21345:data<=-16'd12833;
      21346:data<=-16'd12054;
      21347:data<=-16'd11837;
      21348:data<=-16'd11841;
      21349:data<=-16'd11254;
      21350:data<=-16'd10898;
      21351:data<=-16'd11060;
      21352:data<=-16'd10769;
      21353:data<=-16'd10615;
      21354:data<=-16'd10539;
      21355:data<=-16'd9800;
      21356:data<=-16'd9404;
      21357:data<=-16'd9549;
      21358:data<=-16'd9676;
      21359:data<=-16'd9703;
      21360:data<=-16'd10108;
      21361:data<=-16'd10798;
      21362:data<=-16'd9932;
      21363:data<=-16'd9159;
      21364:data<=-16'd10304;
      21365:data<=-16'd10352;
      21366:data<=-16'd10140;
      21367:data<=-16'd10387;
      21368:data<=-16'd8986;
      21369:data<=-16'd8915;
      21370:data<=-16'd8434;
      21371:data<=-16'd6414;
      21372:data<=-16'd8906;
      21373:data<=-16'd7450;
      21374:data<=16'd3178;
      21375:data<=16'd7300;
      21376:data<=16'd4438;
      21377:data<=16'd5034;
      21378:data<=16'd5106;
      21379:data<=16'd4088;
      21380:data<=16'd5122;
      21381:data<=16'd4957;
      21382:data<=16'd4176;
      21383:data<=16'd4306;
      21384:data<=16'd3964;
      21385:data<=16'd2889;
      21386:data<=16'd1345;
      21387:data<=16'd663;
      21388:data<=16'd526;
      21389:data<=16'd221;
      21390:data<=16'd913;
      21391:data<=16'd558;
      21392:data<=-16'd910;
      21393:data<=-16'd553;
      21394:data<=-16'd428;
      21395:data<=-16'd1057;
      21396:data<=-16'd429;
      21397:data<=-16'd578;
      21398:data<=-16'd1848;
      21399:data<=-16'd2272;
      21400:data<=-16'd1953;
      21401:data<=-16'd1428;
      21402:data<=-16'd1545;
      21403:data<=-16'd2243;
      21404:data<=-16'd2285;
      21405:data<=-16'd2285;
      21406:data<=-16'd2657;
      21407:data<=-16'd2002;
      21408:data<=-16'd1421;
      21409:data<=-16'd2749;
      21410:data<=-16'd2240;
      21411:data<=16'd1660;
      21412:data<=16'd3065;
      21413:data<=16'd1985;
      21414:data<=16'd2419;
      21415:data<=16'd2262;
      21416:data<=16'd1713;
      21417:data<=16'd2009;
      21418:data<=16'd1600;
      21419:data<=16'd1996;
      21420:data<=16'd1751;
      21421:data<=16'd490;
      21422:data<=16'd1512;
      21423:data<=-16'd2273;
      21424:data<=-16'd12571;
      21425:data<=-16'd17023;
      21426:data<=-16'd15544;
      21427:data<=-16'd15059;
      21428:data<=-16'd14316;
      21429:data<=-16'd13923;
      21430:data<=-16'd14504;
      21431:data<=-16'd13732;
      21432:data<=-16'd12352;
      21433:data<=-16'd11615;
      21434:data<=-16'd11775;
      21435:data<=-16'd12589;
      21436:data<=-16'd13112;
      21437:data<=-16'd12730;
      21438:data<=-16'd11212;
      21439:data<=-16'd10220;
      21440:data<=-16'd10457;
      21441:data<=-16'd10151;
      21442:data<=-16'd9476;
      21443:data<=-16'd8884;
      21444:data<=-16'd8411;
      21445:data<=-16'd8314;
      21446:data<=-16'd7770;
      21447:data<=-16'd8492;
      21448:data<=-16'd10460;
      21449:data<=-16'd10146;
      21450:data<=-16'd9262;
      21451:data<=-16'd9238;
      21452:data<=-16'd8169;
      21453:data<=-16'd7686;
      21454:data<=-16'd7823;
      21455:data<=-16'd7001;
      21456:data<=-16'd6545;
      21457:data<=-16'd6631;
      21458:data<=-16'd6807;
      21459:data<=-16'd6795;
      21460:data<=-16'd6595;
      21461:data<=-16'd6933;
      21462:data<=-16'd6504;
      21463:data<=-16'd5835;
      21464:data<=-16'd6096;
      21465:data<=-16'd5483;
      21466:data<=-16'd5278;
      21467:data<=-16'd5463;
      21468:data<=-16'd4275;
      21469:data<=-16'd4554;
      21470:data<=-16'd4400;
      21471:data<=-16'd2713;
      21472:data<=-16'd4525;
      21473:data<=-16'd3777;
      21474:data<=16'd4558;
      21475:data<=16'd11098;
      21476:data<=16'd12081;
      21477:data<=16'd9639;
      21478:data<=16'd4943;
      21479:data<=16'd3257;
      21480:data<=16'd4589;
      21481:data<=16'd4535;
      21482:data<=16'd4237;
      21483:data<=16'd4541;
      21484:data<=16'd4563;
      21485:data<=16'd4121;
      21486:data<=16'd2893;
      21487:data<=16'd2094;
      21488:data<=16'd1830;
      21489:data<=16'd1736;
      21490:data<=16'd2497;
      21491:data<=16'd2369;
      21492:data<=16'd1548;
      21493:data<=16'd1811;
      21494:data<=16'd1571;
      21495:data<=16'd1366;
      21496:data<=16'd2130;
      21497:data<=16'd1971;
      21498:data<=16'd1406;
      21499:data<=16'd901;
      21500:data<=16'd503;
      21501:data<=16'd1168;
      21502:data<=16'd1160;
      21503:data<=16'd975;
      21504:data<=16'd2026;
      21505:data<=16'd2002;
      21506:data<=16'd1674;
      21507:data<=16'd1786;
      21508:data<=16'd1254;
      21509:data<=16'd2003;
      21510:data<=16'd1921;
      21511:data<=-16'd271;
      21512:data<=-16'd238;
      21513:data<=16'd525;
      21514:data<=16'd470;
      21515:data<=16'd1348;
      21516:data<=16'd1122;
      21517:data<=16'd989;
      21518:data<=16'd1773;
      21519:data<=16'd1057;
      21520:data<=16'd1057;
      21521:data<=16'd1215;
      21522:data<=16'd520;
      21523:data<=-16'd149;
      21524:data<=-16'd6613;
      21525:data<=-16'd15371;
      21526:data<=-16'd16140;
      21527:data<=-16'd14058;
      21528:data<=-16'd13972;
      21529:data<=-16'd12924;
      21530:data<=-16'd12445;
      21531:data<=-16'd12575;
      21532:data<=-16'd12005;
      21533:data<=-16'd11038;
      21534:data<=-16'd9474;
      21535:data<=-16'd9620;
      21536:data<=-16'd10833;
      21537:data<=-16'd10386;
      21538:data<=-16'd9386;
      21539:data<=-16'd8182;
      21540:data<=-16'd7412;
      21541:data<=-16'd6936;
      21542:data<=-16'd5739;
      21543:data<=-16'd6021;
      21544:data<=-16'd4554;
      21545:data<=16'd687;
      21546:data<=16'd2375;
      21547:data<=16'd1089;
      21548:data<=16'd1698;
      21549:data<=16'd1956;
      21550:data<=16'd1594;
      21551:data<=16'd1709;
      21552:data<=16'd2258;
      21553:data<=16'd2951;
      21554:data<=16'd2387;
      21555:data<=16'd2387;
      21556:data<=16'd2783;
      21557:data<=16'd2114;
      21558:data<=16'd2943;
      21559:data<=16'd3263;
      21560:data<=16'd2758;
      21561:data<=16'd4667;
      21562:data<=16'd5160;
      21563:data<=16'd4538;
      21564:data<=16'd5436;
      21565:data<=16'd5153;
      21566:data<=16'd5615;
      21567:data<=16'd6032;
      21568:data<=16'd4719;
      21569:data<=16'd5559;
      21570:data<=16'd5568;
      21571:data<=16'd5057;
      21572:data<=16'd6617;
      21573:data<=16'd5752;
      21574:data<=16'd10290;
      21575:data<=16'd21567;
      21576:data<=16'd23840;
      21577:data<=16'd21440;
      21578:data<=16'd22375;
      21579:data<=16'd20619;
      21580:data<=16'd19634;
      21581:data<=16'd20632;
      21582:data<=16'd19287;
      21583:data<=16'd18700;
      21584:data<=16'd17935;
      21585:data<=16'd17001;
      21586:data<=16'd18459;
      21587:data<=16'd18419;
      21588:data<=16'd17199;
      21589:data<=16'd16590;
      21590:data<=16'd15302;
      21591:data<=16'd15098;
      21592:data<=16'd14830;
      21593:data<=16'd13465;
      21594:data<=16'd13233;
      21595:data<=16'd13342;
      21596:data<=16'd13391;
      21597:data<=16'd13188;
      21598:data<=16'd12927;
      21599:data<=16'd13866;
      21600:data<=16'd13684;
      21601:data<=16'd12654;
      21602:data<=16'd12443;
      21603:data<=16'd11634;
      21604:data<=16'd11523;
      21605:data<=16'd11107;
      21606:data<=16'd9928;
      21607:data<=16'd10974;
      21608:data<=16'd10525;
      21609:data<=16'd9191;
      21610:data<=16'd10880;
      21611:data<=16'd9388;
      21612:data<=16'd5043;
      21613:data<=16'd3797;
      21614:data<=16'd3870;
      21615:data<=16'd4168;
      21616:data<=16'd3933;
      21617:data<=16'd3301;
      21618:data<=16'd3639;
      21619:data<=16'd2934;
      21620:data<=16'd3025;
      21621:data<=16'd3013;
      21622:data<=16'd1400;
      21623:data<=16'd3956;
      21624:data<=16'd2132;
      21625:data<=-16'd9288;
      21626:data<=-16'd13080;
      21627:data<=-16'd10119;
      21628:data<=-16'd11409;
      21629:data<=-16'd10727;
      21630:data<=-16'd9106;
      21631:data<=-16'd10398;
      21632:data<=-16'd9911;
      21633:data<=-16'd9356;
      21634:data<=-16'd9544;
      21635:data<=-16'd8257;
      21636:data<=-16'd6912;
      21637:data<=-16'd5617;
      21638:data<=-16'd5139;
      21639:data<=-16'd5080;
      21640:data<=-16'd4331;
      21641:data<=-16'd4880;
      21642:data<=-16'd4952;
      21643:data<=-16'd3755;
      21644:data<=-16'd3929;
      21645:data<=-16'd3859;
      21646:data<=-16'd3477;
      21647:data<=-16'd3718;
      21648:data<=-16'd2478;
      21649:data<=-16'd917;
      21650:data<=-16'd811;
      21651:data<=-16'd1356;
      21652:data<=-16'd1594;
      21653:data<=-16'd1263;
      21654:data<=-16'd1527;
      21655:data<=-16'd1762;
      21656:data<=-16'd1328;
      21657:data<=-16'd1524;
      21658:data<=-16'd1510;
      21659:data<=-16'd1418;
      21660:data<=-16'd1243;
      21661:data<=16'd391;
      21662:data<=16'd1014;
      21663:data<=16'd705;
      21664:data<=16'd1102;
      21665:data<=16'd196;
      21666:data<=-16'd294;
      21667:data<=16'd187;
      21668:data<=-16'd238;
      21669:data<=16'd167;
      21670:data<=16'd103;
      21671:data<=16'd56;
      21672:data<=16'd1301;
      21673:data<=16'd403;
      21674:data<=16'd4410;
      21675:data<=16'd15370;
      21676:data<=16'd18061;
      21677:data<=16'd14798;
      21678:data<=16'd17653;
      21679:data<=16'd20618;
      21680:data<=16'd19845;
      21681:data<=16'd19610;
      21682:data<=16'd19423;
      21683:data<=16'd18342;
      21684:data<=16'd16833;
      21685:data<=16'd16427;
      21686:data<=16'd17306;
      21687:data<=16'd16678;
      21688:data<=16'd15247;
      21689:data<=16'd14404;
      21690:data<=16'd13438;
      21691:data<=16'd13083;
      21692:data<=16'd12747;
      21693:data<=16'd11852;
      21694:data<=16'd11223;
      21695:data<=16'd10443;
      21696:data<=16'd9682;
      21697:data<=16'd8969;
      21698:data<=16'd8942;
      21699:data<=16'd10273;
      21700:data<=16'd10311;
      21701:data<=16'd9432;
      21702:data<=16'd9562;
      21703:data<=16'd8540;
      21704:data<=16'd7289;
      21705:data<=16'd7374;
      21706:data<=16'd7068;
      21707:data<=16'd6722;
      21708:data<=16'd5937;
      21709:data<=16'd4751;
      21710:data<=16'd5468;
      21711:data<=16'd6454;
      21712:data<=16'd5912;
      21713:data<=16'd5089;
      21714:data<=16'd4687;
      21715:data<=16'd4599;
      21716:data<=16'd4112;
      21717:data<=16'd3952;
      21718:data<=16'd3817;
      21719:data<=16'd2481;
      21720:data<=16'd2599;
      21721:data<=16'd2359;
      21722:data<=16'd315;
      21723:data<=16'd1980;
      21724:data<=16'd453;
      21725:data<=-16'd9653;
      21726:data<=-16'd14195;
      21727:data<=-16'd11920;
      21728:data<=-16'd12800;
      21729:data<=-16'd12977;
      21730:data<=-16'd11784;
      21731:data<=-16'd12833;
      21732:data<=-16'd12569;
      21733:data<=-16'd11703;
      21734:data<=-16'd12078;
      21735:data<=-16'd11350;
      21736:data<=-16'd10295;
      21737:data<=-16'd9708;
      21738:data<=-16'd8919;
      21739:data<=-16'd8713;
      21740:data<=-16'd8963;
      21741:data<=-16'd9031;
      21742:data<=-16'd8893;
      21743:data<=-16'd8213;
      21744:data<=-16'd7708;
      21745:data<=-16'd9837;
      21746:data<=-16'd13659;
      21747:data<=-16'd14653;
      21748:data<=-16'd13693;
      21749:data<=-16'd13825;
      21750:data<=-16'd13577;
      21751:data<=-16'd13312;
      21752:data<=-16'd13529;
      21753:data<=-16'd12562;
      21754:data<=-16'd12093;
      21755:data<=-16'd12304;
      21756:data<=-16'd11734;
      21757:data<=-16'd11617;
      21758:data<=-16'd11288;
      21759:data<=-16'd10593;
      21760:data<=-16'd11030;
      21761:data<=-16'd11878;
      21762:data<=-16'd12654;
      21763:data<=-16'd12343;
      21764:data<=-16'd11062;
      21765:data<=-16'd11113;
      21766:data<=-16'd11382;
      21767:data<=-16'd11048;
      21768:data<=-16'd10699;
      21769:data<=-16'd10035;
      21770:data<=-16'd10437;
      21771:data<=-16'd9850;
      21772:data<=-16'd8410;
      21773:data<=-16'd10507;
      21774:data<=-16'd8637;
      21775:data<=16'd849;
      21776:data<=16'd5488;
      21777:data<=16'd4061;
      21778:data<=16'd3861;
      21779:data<=16'd3533;
      21780:data<=16'd3075;
      21781:data<=16'd3518;
      21782:data<=16'd3336;
      21783:data<=16'd3093;
      21784:data<=16'd2635;
      21785:data<=16'd1967;
      21786:data<=16'd1403;
      21787:data<=16'd249;
      21788:data<=-16'd165;
      21789:data<=16'd3;
      21790:data<=-16'd350;
      21791:data<=-16'd197;
      21792:data<=-16'd221;
      21793:data<=-16'd537;
      21794:data<=-16'd282;
      21795:data<=-16'd607;
      21796:data<=-16'd931;
      21797:data<=-16'd526;
      21798:data<=-16'd738;
      21799:data<=-16'd1830;
      21800:data<=-16'd2825;
      21801:data<=-16'd2634;
      21802:data<=-16'd2381;
      21803:data<=-16'd3206;
      21804:data<=-16'd3287;
      21805:data<=-16'd2966;
      21806:data<=-16'd2851;
      21807:data<=-16'd2127;
      21808:data<=-16'd2466;
      21809:data<=-16'd2729;
      21810:data<=-16'd2244;
      21811:data<=-16'd3486;
      21812:data<=-16'd2403;
      21813:data<=16'd1744;
      21814:data<=16'd2423;
      21815:data<=16'd1245;
      21816:data<=16'd1559;
      21817:data<=16'd1905;
      21818:data<=16'd2165;
      21819:data<=16'd1412;
      21820:data<=16'd588;
      21821:data<=16'd1246;
      21822:data<=16'd1528;
      21823:data<=16'd1522;
      21824:data<=-16'd1980;
      21825:data<=-16'd11157;
      21826:data<=-16'd16736;
      21827:data<=-16'd15941;
      21828:data<=-16'd15488;
      21829:data<=-16'd15050;
      21830:data<=-16'd13943;
      21831:data<=-16'd14014;
      21832:data<=-16'd13634;
      21833:data<=-16'd12747;
      21834:data<=-16'd12229;
      21835:data<=-16'd11837;
      21836:data<=-16'd12314;
      21837:data<=-16'd13013;
      21838:data<=-16'd12659;
      21839:data<=-16'd11761;
      21840:data<=-16'd11197;
      21841:data<=-16'd10719;
      21842:data<=-16'd9953;
      21843:data<=-16'd9608;
      21844:data<=-16'd9263;
      21845:data<=-16'd8434;
      21846:data<=-16'd8014;
      21847:data<=-16'd7517;
      21848:data<=-16'd7918;
      21849:data<=-16'd9800;
      21850:data<=-16'd9712;
      21851:data<=-16'd8490;
      21852:data<=-16'd8587;
      21853:data<=-16'd7843;
      21854:data<=-16'd6858;
      21855:data<=-16'd6798;
      21856:data<=-16'd6443;
      21857:data<=-16'd6484;
      21858:data<=-16'd6288;
      21859:data<=-16'd5538;
      21860:data<=-16'd5503;
      21861:data<=-16'd5606;
      21862:data<=-16'd6598;
      21863:data<=-16'd7518;
      21864:data<=-16'd6167;
      21865:data<=-16'd5295;
      21866:data<=-16'd5363;
      21867:data<=-16'd4814;
      21868:data<=-16'd4657;
      21869:data<=-16'd3850;
      21870:data<=-16'd3577;
      21871:data<=-16'd4326;
      21872:data<=-16'd2843;
      21873:data<=-16'd3157;
      21874:data<=-16'd4579;
      21875:data<=16'd2159;
      21876:data<=16'd10687;
      21877:data<=16'd11568;
      21878:data<=16'd10246;
      21879:data<=16'd8375;
      21880:data<=16'd4573;
      21881:data<=16'd3601;
      21882:data<=16'd4581;
      21883:data<=16'd4299;
      21884:data<=16'd4438;
      21885:data<=16'd4561;
      21886:data<=16'd3573;
      21887:data<=16'd2452;
      21888:data<=16'd1539;
      21889:data<=16'd1579;
      21890:data<=16'd2203;
      21891:data<=16'd2043;
      21892:data<=16'd1851;
      21893:data<=16'd2015;
      21894:data<=16'd1895;
      21895:data<=16'd1926;
      21896:data<=16'd2526;
      21897:data<=16'd3247;
      21898:data<=16'd2845;
      21899:data<=16'd1403;
      21900:data<=16'd669;
      21901:data<=16'd655;
      21902:data<=16'd823;
      21903:data<=16'd1213;
      21904:data<=16'd1096;
      21905:data<=16'd939;
      21906:data<=16'd1380;
      21907:data<=16'd1747;
      21908:data<=16'd1891;
      21909:data<=16'd1980;
      21910:data<=16'd2249;
      21911:data<=16'd1744;
      21912:data<=16'd85;
      21913:data<=-16'd80;
      21914:data<=16'd682;
      21915:data<=16'd420;
      21916:data<=16'd952;
      21917:data<=16'd1600;
      21918:data<=16'd1310;
      21919:data<=16'd1207;
      21920:data<=16'd1011;
      21921:data<=16'd1788;
      21922:data<=16'd2265;
      21923:data<=16'd1436;
      21924:data<=16'd1438;
      21925:data<=-16'd3880;
      21926:data<=-16'd13910;
      21927:data<=-16'd15835;
      21928:data<=-16'd13157;
      21929:data<=-16'd13515;
      21930:data<=-16'd12634;
      21931:data<=-16'd11814;
      21932:data<=-16'd11991;
      21933:data<=-16'd10690;
      21934:data<=-16'd10025;
      21935:data<=-16'd8980;
      21936:data<=-16'd8531;
      21937:data<=-16'd10228;
      21938:data<=-16'd9409;
      21939:data<=-16'd7897;
      21940:data<=-16'd8269;
      21941:data<=-16'd7356;
      21942:data<=-16'd6454;
      21943:data<=-16'd6217;
      21944:data<=-16'd5871;
      21945:data<=-16'd5480;
      21946:data<=-16'd2097;
      21947:data<=16'd1870;
      21948:data<=16'd2399;
      21949:data<=16'd2273;
      21950:data<=16'd2510;
      21951:data<=16'd2504;
      21952:data<=16'd3153;
      21953:data<=16'd3742;
      21954:data<=16'd3944;
      21955:data<=16'd4167;
      21956:data<=16'd4249;
      21957:data<=16'd3802;
      21958:data<=16'd3612;
      21959:data<=16'd4275;
      21960:data<=16'd4105;
      21961:data<=16'd4739;
      21962:data<=16'd6805;
      21963:data<=16'd6308;
      21964:data<=16'd5703;
      21965:data<=16'd6737;
      21966:data<=16'd6178;
      21967:data<=16'd6100;
      21968:data<=16'd6253;
      21969:data<=16'd5929;
      21970:data<=16'd6930;
      21971:data<=16'd5909;
      21972:data<=16'd5664;
      21973:data<=16'd7304;
      21974:data<=16'd5903;
      21975:data<=16'd11201;
      21976:data<=16'd22773;
      21977:data<=16'd24589;
      21978:data<=16'd21966;
      21979:data<=16'd22371;
      21980:data<=16'd21346;
      21981:data<=16'd20979;
      21982:data<=16'd20535;
      21983:data<=16'd19191;
      21984:data<=16'd19544;
      21985:data<=16'd18177;
      21986:data<=16'd17279;
      21987:data<=16'd19074;
      21988:data<=16'd18594;
      21989:data<=16'd17424;
      21990:data<=16'd17165;
      21991:data<=16'd16363;
      21992:data<=16'd16184;
      21993:data<=16'd15414;
      21994:data<=16'd14549;
      21995:data<=16'd14351;
      21996:data<=16'd13265;
      21997:data<=16'd13054;
      21998:data<=16'd13271;
      21999:data<=16'd13262;
      22000:data<=16'd14246;
      22001:data<=16'd13459;
      22002:data<=16'd12113;
      22003:data<=16'd12340;
      22004:data<=16'd11439;
      22005:data<=16'd10775;
      22006:data<=16'd10712;
      22007:data<=16'd9800;
      22008:data<=16'd10008;
      22009:data<=16'd9659;
      22010:data<=16'd8375;
      22011:data<=16'd9072;
      22012:data<=16'd9529;
      22013:data<=16'd7250;
      22014:data<=16'd3576;
      22015:data<=16'd1952;
      22016:data<=16'd2937;
      22017:data<=16'd2836;
      22018:data<=16'd2684;
      22019:data<=16'd2934;
      22020:data<=16'd1607;
      22021:data<=16'd2168;
      22022:data<=16'd2382;
      22023:data<=16'd1021;
      22024:data<=16'd3691;
      22025:data<=16'd1151;
      22026:data<=-16'd10178;
      22027:data<=-16'd14054;
      22028:data<=-16'd11209;
      22029:data<=-16'd11435;
      22030:data<=-16'd11171;
      22031:data<=-16'd10369;
      22032:data<=-16'd10624;
      22033:data<=-16'd9897;
      22034:data<=-16'd9950;
      22035:data<=-16'd9881;
      22036:data<=-16'd8404;
      22037:data<=-16'd7511;
      22038:data<=-16'd6573;
      22039:data<=-16'd5962;
      22040:data<=-16'd6164;
      22041:data<=-16'd5583;
      22042:data<=-16'd5200;
      22043:data<=-16'd5160;
      22044:data<=-16'd4772;
      22045:data<=-16'd5060;
      22046:data<=-16'd4899;
      22047:data<=-16'd4279;
      22048:data<=-16'd4602;
      22049:data<=-16'd3689;
      22050:data<=-16'd1601;
      22051:data<=-16'd1228;
      22052:data<=-16'd1309;
      22053:data<=-16'd763;
      22054:data<=-16'd1108;
      22055:data<=-16'd1269;
      22056:data<=-16'd740;
      22057:data<=-16'd1074;
      22058:data<=-16'd1099;
      22059:data<=-16'd775;
      22060:data<=-16'd1439;
      22061:data<=-16'd637;
      22062:data<=16'd1260;
      22063:data<=16'd1064;
      22064:data<=16'd629;
      22065:data<=16'd1011;
      22066:data<=16'd952;
      22067:data<=16'd975;
      22068:data<=16'd393;
      22069:data<=16'd126;
      22070:data<=16'd926;
      22071:data<=16'd352;
      22072:data<=16'd423;
      22073:data<=16'd1033;
      22074:data<=-16'd303;
      22075:data<=16'd4637;
      22076:data<=16'd15925;
      22077:data<=16'd19273;
      22078:data<=16'd15879;
      22079:data<=16'd16365;
      22080:data<=16'd19516;
      22081:data<=16'd21217;
      22082:data<=16'd20663;
      22083:data<=16'd19259;
      22084:data<=16'd18812;
      22085:data<=16'd17713;
      22086:data<=16'd16948;
      22087:data<=16'd18266;
      22088:data<=16'd18175;
      22089:data<=16'd16706;
      22090:data<=16'd16384;
      22091:data<=16'd15687;
      22092:data<=16'd14577;
      22093:data<=16'd14023;
      22094:data<=16'd13362;
      22095:data<=16'd12821;
      22096:data<=16'd12246;
      22097:data<=16'd11392;
      22098:data<=16'd10696;
      22099:data<=16'd10446;
      22100:data<=16'd11162;
      22101:data<=16'd11539;
      22102:data<=16'd10339;
      22103:data<=16'd9374;
      22104:data<=16'd9282;
      22105:data<=16'd8815;
      22106:data<=16'd7891;
      22107:data<=16'd7163;
      22108:data<=16'd6904;
      22109:data<=16'd6369;
      22110:data<=16'd5597;
      22111:data<=16'd5679;
      22112:data<=16'd6178;
      22113:data<=16'd6473;
      22114:data<=16'd6440;
      22115:data<=16'd5780;
      22116:data<=16'd5028;
      22117:data<=16'd4613;
      22118:data<=16'd4469;
      22119:data<=16'd3644;
      22120:data<=16'd2288;
      22121:data<=16'd2535;
      22122:data<=16'd2087;
      22123:data<=16'd722;
      22124:data<=16'd2945;
      22125:data<=16'd1234;
      22126:data<=-16'd8981;
      22127:data<=-16'd14108;
      22128:data<=-16'd12226;
      22129:data<=-16'd12575;
      22130:data<=-16'd12787;
      22131:data<=-16'd11941;
      22132:data<=-16'd12480;
      22133:data<=-16'd12034;
      22134:data<=-16'd11800;
      22135:data<=-16'd12363;
      22136:data<=-16'd11582;
      22137:data<=-16'd10693;
      22138:data<=-16'd9643;
      22139:data<=-16'd8349;
      22140:data<=-16'd8624;
      22141:data<=-16'd9236;
      22142:data<=-16'd8760;
      22143:data<=-16'd8392;
      22144:data<=-16'd8781;
      22145:data<=-16'd8633;
      22146:data<=-16'd8907;
      22147:data<=-16'd12228;
      22148:data<=-16'd14857;
      22149:data<=-16'd13879;
      22150:data<=-16'd13582;
      22151:data<=-16'd13885;
      22152:data<=-16'd12859;
      22153:data<=-16'd12674;
      22154:data<=-16'd12780;
      22155:data<=-16'd12515;
      22156:data<=-16'd12521;
      22157:data<=-16'd12137;
      22158:data<=-16'd12011;
      22159:data<=-16'd11735;
      22160:data<=-16'd11086;
      22161:data<=-16'd11212;
      22162:data<=-16'd11426;
      22163:data<=-16'd12220;
      22164:data<=-16'd13015;
      22165:data<=-16'd12207;
      22166:data<=-16'd11641;
      22167:data<=-16'd11235;
      22168:data<=-16'd10930;
      22169:data<=-16'd11423;
      22170:data<=-16'd10505;
      22171:data<=-16'd10243;
      22172:data<=-16'd10549;
      22173:data<=-16'd8927;
      22174:data<=-16'd10558;
      22175:data<=-16'd10508;
      22176:data<=-16'd1074;
      22177:data<=16'd5426;
      22178:data<=16'd4067;
      22179:data<=16'd4047;
      22180:data<=16'd4479;
      22181:data<=16'd3629;
      22182:data<=16'd3604;
      22183:data<=16'd3210;
      22184:data<=16'd3143;
      22185:data<=16'd3424;
      22186:data<=16'd2914;
      22187:data<=16'd2240;
      22188:data<=16'd914;
      22189:data<=-16'd127;
      22190:data<=-16'd23;
      22191:data<=-16'd59;
      22192:data<=-16'd190;
      22193:data<=-16'd669;
      22194:data<=-16'd1187;
      22195:data<=-16'd795;
      22196:data<=-16'd789;
      22197:data<=-16'd1052;
      22198:data<=-16'd1090;
      22199:data<=-16'd2032;
      22200:data<=-16'd3099;
      22201:data<=-16'd3624;
      22202:data<=-16'd3974;
      22203:data<=-16'd4021;
      22204:data<=-16'd3871;
      22205:data<=-16'd3312;
      22206:data<=-16'd3093;
      22207:data<=-16'd3541;
      22208:data<=-16'd3430;
      22209:data<=-16'd3480;
      22210:data<=-16'd3351;
      22211:data<=-16'd2810;
      22212:data<=-16'd4499;
      22213:data<=-16'd5077;
      22214:data<=-16'd1124;
      22215:data<=16'd1489;
      22216:data<=16'd911;
      22217:data<=16'd869;
      22218:data<=16'd823;
      22219:data<=16'd359;
      22220:data<=16'd270;
      22221:data<=16'd475;
      22222:data<=16'd983;
      22223:data<=16'd614;
      22224:data<=16'd317;
      22225:data<=-16'd1189;
      22226:data<=-16'd9119;
      22227:data<=-16'd17164;
      22228:data<=-16'd17145;
      22229:data<=-16'd15676;
      22230:data<=-16'd15854;
      22231:data<=-16'd14487;
      22232:data<=-16'd14404;
      22233:data<=-16'd14659;
      22234:data<=-16'd13132;
      22235:data<=-16'd12703;
      22236:data<=-16'd12342;
      22237:data<=-16'd12116;
      22238:data<=-16'd13435;
      22239:data<=-16'd12974;
      22240:data<=-16'd11618;
      22241:data<=-16'd11543;
      22242:data<=-16'd10759;
      22243:data<=-16'd10119;
      22244:data<=-16'd9940;
      22245:data<=-16'd9273;
      22246:data<=-16'd9374;
      22247:data<=-16'd8862;
      22248:data<=-16'd7420;
      22249:data<=-16'd7941;
      22250:data<=-16'd9467;
      22251:data<=-16'd9538;
      22252:data<=-16'd8669;
      22253:data<=-16'd8067;
      22254:data<=-16'd7711;
      22255:data<=-16'd7447;
      22256:data<=-16'd7462;
      22257:data<=-16'd6855;
      22258:data<=-16'd5877;
      22259:data<=-16'd5741;
      22260:data<=-16'd5357;
      22261:data<=-16'd4751;
      22262:data<=-16'd5095;
      22263:data<=-16'd6028;
      22264:data<=-16'd6789;
      22265:data<=-16'd6059;
      22266:data<=-16'd5134;
      22267:data<=-16'd5506;
      22268:data<=-16'd4919;
      22269:data<=-16'd4138;
      22270:data<=-16'd3988;
      22271:data<=-16'd3580;
      22272:data<=-16'd4282;
      22273:data<=-16'd3312;
      22274:data<=-16'd2511;
      22275:data<=-16'd5298;
      22276:data<=-16'd344;
      22277:data<=16'd10590;
      22278:data<=16'd12286;
      22279:data<=16'd10925;
      22280:data<=16'd11160;
      22281:data<=16'd6793;
      22282:data<=16'd4173;
      22283:data<=16'd4910;
      22284:data<=16'd4106;
      22285:data<=16'd4625;
      22286:data<=16'd5236;
      22287:data<=16'd4094;
      22288:data<=16'd3128;
      22289:data<=16'd1936;
      22290:data<=16'd1886;
      22291:data<=16'd2394;
      22292:data<=16'd1888;
      22293:data<=16'd2293;
      22294:data<=16'd2479;
      22295:data<=16'd2091;
      22296:data<=16'd2476;
      22297:data<=16'd2369;
      22298:data<=16'd2584;
      22299:data<=16'd2719;
      22300:data<=16'd1360;
      22301:data<=16'd617;
      22302:data<=16'd387;
      22303:data<=16'd44;
      22304:data<=16'd469;
      22305:data<=16'd763;
      22306:data<=16'd922;
      22307:data<=16'd911;
      22308:data<=16'd549;
      22309:data<=16'd760;
      22310:data<=16'd1422;
      22311:data<=16'd2196;
      22312:data<=16'd1151;
      22313:data<=-16'd1263;
      22314:data<=-16'd942;
      22315:data<=-16'd183;
      22316:data<=-16'd804;
      22317:data<=16'd62;
      22318:data<=16'd321;
      22319:data<=-16'd12;
      22320:data<=16'd617;
      22321:data<=16'd526;
      22322:data<=16'd1613;
      22323:data<=16'd1989;
      22324:data<=16'd678;
      22325:data<=16'd1624;
      22326:data<=-16'd3237;
      22327:data<=-16'd14384;
      22328:data<=-16'd17027;
      22329:data<=-16'd14487;
      22330:data<=-16'd14901;
      22331:data<=-16'd13885;
      22332:data<=-16'd12803;
      22333:data<=-16'd12748;
      22334:data<=-16'd11132;
      22335:data<=-16'd10125;
      22336:data<=-16'd9476;
      22337:data<=-16'd9439;
      22338:data<=-16'd10836;
      22339:data<=-16'd10352;
      22340:data<=-16'd9141;
      22341:data<=-16'd8809;
      22342:data<=-16'd7768;
      22343:data<=-16'd7262;
      22344:data<=-16'd6552;
      22345:data<=-16'd5520;
      22346:data<=-16'd6100;
      22347:data<=-16'd4317;
      22348:data<=16'd588;
      22349:data<=16'd2776;
      22350:data<=16'd2362;
      22351:data<=16'd2661;
      22352:data<=16'd3128;
      22353:data<=16'd3334;
      22354:data<=16'd4090;
      22355:data<=16'd4546;
      22356:data<=16'd4185;
      22357:data<=16'd4370;
      22358:data<=16'd4918;
      22359:data<=16'd5095;
      22360:data<=16'd5053;
      22361:data<=16'd4435;
      22362:data<=16'd5162;
      22363:data<=16'd7218;
      22364:data<=16'd7078;
      22365:data<=16'd6570;
      22366:data<=16'd7163;
      22367:data<=16'd6830;
      22368:data<=16'd7071;
      22369:data<=16'd7191;
      22370:data<=16'd6722;
      22371:data<=16'd7474;
      22372:data<=16'd6866;
      22373:data<=16'd7036;
      22374:data<=16'd8664;
      22375:data<=16'd7212;
      22376:data<=16'd11761;
      22377:data<=16'd23341;
      22378:data<=16'd26159;
      22379:data<=16'd23705;
      22380:data<=16'd24260;
      22381:data<=16'd22801;
      22382:data<=16'd21763;
      22383:data<=16'd22195;
      22384:data<=16'd20407;
      22385:data<=16'd19691;
      22386:data<=16'd19432;
      22387:data<=16'd18795;
      22388:data<=16'd20039;
      22389:data<=16'd19506;
      22390:data<=16'd17628;
      22391:data<=16'd17778;
      22392:data<=16'd17676;
      22393:data<=16'd16745;
      22394:data<=16'd15643;
      22395:data<=16'd14827;
      22396:data<=16'd15192;
      22397:data<=16'd14686;
      22398:data<=16'd13421;
      22399:data<=16'd13251;
      22400:data<=16'd13438;
      22401:data<=16'd13944;
      22402:data<=16'd14063;
      22403:data<=16'd13150;
      22404:data<=16'd12684;
      22405:data<=16'd12498;
      22406:data<=16'd12046;
      22407:data<=16'd11304;
      22408:data<=16'd10275;
      22409:data<=16'd10173;
      22410:data<=16'd10214;
      22411:data<=16'd9172;
      22412:data<=16'd8752;
      22413:data<=16'd9380;
      22414:data<=16'd8542;
      22415:data<=16'd5688;
      22416:data<=16'd4361;
      22417:data<=16'd4808;
      22418:data<=16'd3794;
      22419:data<=16'd3280;
      22420:data<=16'd3644;
      22421:data<=16'd2676;
      22422:data<=16'd3001;
      22423:data<=16'd2611;
      22424:data<=16'd1063;
      22425:data<=16'd3412;
      22426:data<=16'd1005;
      22427:data<=-16'd9579;
      22428:data<=-16'd13700;
      22429:data<=-16'd11600;
      22430:data<=-16'd11881;
      22431:data<=-16'd11570;
      22432:data<=-16'd10927;
      22433:data<=-16'd11141;
      22434:data<=-16'd9824;
      22435:data<=-16'd9254;
      22436:data<=-16'd9538;
      22437:data<=-16'd8636;
      22438:data<=-16'd7412;
      22439:data<=-16'd6072;
      22440:data<=-16'd5676;
      22441:data<=-16'd6440;
      22442:data<=-16'd6579;
      22443:data<=-16'd6378;
      22444:data<=-16'd5739;
      22445:data<=-16'd4931;
      22446:data<=-16'd5380;
      22447:data<=-16'd5642;
      22448:data<=-16'd5207;
      22449:data<=-16'd5210;
      22450:data<=-16'd4093;
      22451:data<=-16'd1958;
      22452:data<=-16'd1613;
      22453:data<=-16'd2240;
      22454:data<=-16'd1712;
      22455:data<=-16'd1536;
      22456:data<=-16'd1977;
      22457:data<=-16'd1528;
      22458:data<=-16'd1735;
      22459:data<=-16'd2238;
      22460:data<=-16'd1559;
      22461:data<=-16'd1879;
      22462:data<=-16'd1519;
      22463:data<=16'd1052;
      22464:data<=16'd1515;
      22465:data<=16'd693;
      22466:data<=16'd881;
      22467:data<=16'd500;
      22468:data<=16'd920;
      22469:data<=16'd1489;
      22470:data<=16'd928;
      22471:data<=16'd1122;
      22472:data<=16'd669;
      22473:data<=16'd634;
      22474:data<=16'd1648;
      22475:data<=16'd513;
      22476:data<=16'd4109;
      22477:data<=16'd14267;
      22478:data<=16'd18475;
      22479:data<=16'd16677;
      22480:data<=16'd16342;
      22481:data<=16'd17035;
      22482:data<=16'd18692;
      22483:data<=16'd19220;
      22484:data<=16'd17344;
      22485:data<=16'd16722;
      22486:data<=16'd16178;
      22487:data<=16'd15509;
      22488:data<=16'd16838;
      22489:data<=16'd16739;
      22490:data<=16'd15270;
      22491:data<=16'd15186;
      22492:data<=16'd14938;
      22493:data<=16'd14319;
      22494:data<=16'd13415;
      22495:data<=16'd11969;
      22496:data<=16'd11462;
      22497:data<=16'd10978;
      22498:data<=16'd9834;
      22499:data<=16'd9274;
      22500:data<=16'd9072;
      22501:data<=16'd9221;
      22502:data<=16'd9529;
      22503:data<=16'd9218;
      22504:data<=16'd8552;
      22505:data<=16'd7561;
      22506:data<=16'd6731;
      22507:data<=16'd6628;
      22508:data<=16'd6563;
      22509:data<=16'd6244;
      22510:data<=16'd5523;
      22511:data<=16'd4593;
      22512:data<=16'd4135;
      22513:data<=16'd4087;
      22514:data<=16'd4454;
      22515:data<=16'd4657;
      22516:data<=16'd4300;
      22517:data<=16'd3993;
      22518:data<=16'd3109;
      22519:data<=16'd2020;
      22520:data<=16'd1445;
      22521:data<=16'd813;
      22522:data<=16'd1316;
      22523:data<=16'd1290;
      22524:data<=-16'd303;
      22525:data<=16'd1128;
      22526:data<=16'd560;
      22527:data<=-16'd8216;
      22528:data<=-16'd14518;
      22529:data<=-16'd13696;
      22530:data<=-16'd13747;
      22531:data<=-16'd14280;
      22532:data<=-16'd13176;
      22533:data<=-16'd12877;
      22534:data<=-16'd12601;
      22535:data<=-16'd12081;
      22536:data<=-16'd12028;
      22537:data<=-16'd11634;
      22538:data<=-16'd11006;
      22539:data<=-16'd10031;
      22540:data<=-16'd9103;
      22541:data<=-16'd9136;
      22542:data<=-16'd9420;
      22543:data<=-16'd9468;
      22544:data<=-16'd9063;
      22545:data<=-16'd8390;
      22546:data<=-16'd8354;
      22547:data<=-16'd8552;
      22548:data<=-16'd9429;
      22549:data<=-16'd11553;
      22550:data<=-16'd12584;
      22551:data<=-16'd11903;
      22552:data<=-16'd11580;
      22553:data<=-16'd11594;
      22554:data<=-16'd11038;
      22555:data<=-16'd10727;
      22556:data<=-16'd11082;
      22557:data<=-16'd11077;
      22558:data<=-16'd10883;
      22559:data<=-16'd10931;
      22560:data<=-16'd10270;
      22561:data<=-16'd9843;
      22562:data<=-16'd10392;
      22563:data<=-16'd10352;
      22564:data<=-16'd10357;
      22565:data<=-16'd10611;
      22566:data<=-16'd9920;
      22567:data<=-16'd9565;
      22568:data<=-16'd9354;
      22569:data<=-16'd8516;
      22570:data<=-16'd8076;
      22571:data<=-16'd7573;
      22572:data<=-16'd7759;
      22573:data<=-16'd8234;
      22574:data<=-16'd7442;
      22575:data<=-16'd8874;
      22576:data<=-16'd9204;
      22577:data<=-16'd1234;
      22578:data<=16'd6696;
      22579:data<=16'd7062;
      22580:data<=16'd5796;
      22581:data<=16'd5386;
      22582:data<=16'd4860;
      22583:data<=16'd4819;
      22584:data<=16'd4141;
      22585:data<=16'd3568;
      22586:data<=16'd3839;
      22587:data<=16'd3694;
      22588:data<=16'd2934;
      22589:data<=16'd1350;
      22590:data<=16'd312;
      22591:data<=16'd913;
      22592:data<=16'd1014;
      22593:data<=16'd590;
      22594:data<=16'd613;
      22595:data<=16'd519;
      22596:data<=16'd629;
      22597:data<=16'd367;
      22598:data<=-16'd20;
      22599:data<=16'd341;
      22600:data<=-16'd667;
      22601:data<=-16'd2431;
      22602:data<=-16'd2552;
      22603:data<=-16'd2626;
      22604:data<=-16'd3098;
      22605:data<=-16'd2989;
      22606:data<=-16'd3022;
      22607:data<=-16'd3019;
      22608:data<=-16'd2739;
      22609:data<=-16'd2573;
      22610:data<=-16'd2673;
      22611:data<=-16'd2804;
      22612:data<=-16'd2409;
      22613:data<=-16'd3366;
      22614:data<=-16'd5651;
      22615:data<=-16'd4757;
      22616:data<=-16'd1845;
      22617:data<=-16'd1136;
      22618:data<=-16'd1300;
      22619:data<=-16'd1474;
      22620:data<=-16'd2020;
      22621:data<=-16'd1861;
      22622:data<=-16'd1368;
      22623:data<=-16'd896;
      22624:data<=-16'd943;
      22625:data<=-16'd1313;
      22626:data<=-16'd2002;
      22627:data<=-16'd7943;
      22628:data<=-16'd17101;
      22629:data<=-16'd19603;
      22630:data<=-16'd17928;
      22631:data<=-16'd17828;
      22632:data<=-16'd16407;
      22633:data<=-16'd14983;
      22634:data<=-16'd15205;
      22635:data<=-16'd14481;
      22636:data<=-16'd13935;
      22637:data<=-16'd13653;
      22638:data<=-16'd13282;
      22639:data<=-16'd14324;
      22640:data<=-16'd14264;
      22641:data<=-16'd12857;
      22642:data<=-16'd12631;
      22643:data<=-16'd12246;
      22644:data<=-16'd11703;
      22645:data<=-16'd11515;
      22646:data<=-16'd10745;
      22647:data<=-16'd10514;
      22648:data<=-16'd10194;
      22649:data<=-16'd9045;
      22650:data<=-16'd9130;
      22651:data<=-16'd10079;
      22652:data<=-16'd10299;
      22653:data<=-16'd9730;
      22654:data<=-16'd8859;
      22655:data<=-16'd8379;
      22656:data<=-16'd7978;
      22657:data<=-16'd7676;
      22658:data<=-16'd7668;
      22659:data<=-16'd7125;
      22660:data<=-16'd6428;
      22661:data<=-16'd5752;
      22662:data<=-16'd5163;
      22663:data<=-16'd5755;
      22664:data<=-16'd6449;
      22665:data<=-16'd6187;
      22666:data<=-16'd5785;
      22667:data<=-16'd5368;
      22668:data<=-16'd4896;
      22669:data<=-16'd4350;
      22670:data<=-16'd3795;
      22671:data<=-16'd3092;
      22672:data<=-16'd2725;
      22673:data<=-16'd3748;
      22674:data<=-16'd3190;
      22675:data<=-16'd2155;
      22676:data<=-16'd4643;
      22677:data<=-16'd917;
      22678:data<=16'd10431;
      22679:data<=16'd13276;
      22680:data<=16'd10646;
      22681:data<=16'd12151;
      22682:data<=16'd10598;
      22683:data<=16'd6851;
      22684:data<=16'd6338;
      22685:data<=16'd5749;
      22686:data<=16'd5698;
      22687:data<=16'd5955;
      22688:data<=16'd4234;
      22689:data<=16'd3278;
      22690:data<=16'd3110;
      22691:data<=16'd2646;
      22692:data<=16'd3001;
      22693:data<=16'd3427;
      22694:data<=16'd3479;
      22695:data<=16'd3269;
      22696:data<=16'd3190;
      22697:data<=16'd3630;
      22698:data<=16'd3689;
      22699:data<=16'd3671;
      22700:data<=16'd3368;
      22701:data<=16'd2088;
      22702:data<=16'd1145;
      22703:data<=16'd881;
      22704:data<=16'd1084;
      22705:data<=16'd1199;
      22706:data<=16'd776;
      22707:data<=16'd1325;
      22708:data<=16'd1976;
      22709:data<=16'd1847;
      22710:data<=16'd2003;
      22711:data<=16'd1515;
      22712:data<=16'd1600;
      22713:data<=16'd2032;
      22714:data<=16'd194;
      22715:data<=-16'd734;
      22716:data<=-16'd412;
      22717:data<=-16'd1177;
      22718:data<=-16'd685;
      22719:data<=-16'd265;
      22720:data<=-16'd749;
      22721:data<=-16'd446;
      22722:data<=-16'd651;
      22723:data<=16'd94;
      22724:data<=16'd472;
      22725:data<=-16'd365;
      22726:data<=16'd1152;
      22727:data<=-16'd3383;
      22728:data<=-16'd14941;
      22729:data<=-16'd17983;
      22730:data<=-16'd15399;
      22731:data<=-16'd15796;
      22732:data<=-16'd14505;
      22733:data<=-16'd13113;
      22734:data<=-16'd13013;
      22735:data<=-16'd11414;
      22736:data<=-16'd10836;
      22737:data<=-16'd10322;
      22738:data<=-16'd9621;
      22739:data<=-16'd11010;
      22740:data<=-16'd10874;
      22741:data<=-16'd9336;
      22742:data<=-16'd9404;
      22743:data<=-16'd9004;
      22744:data<=-16'd8075;
      22745:data<=-16'd7806;
      22746:data<=-16'd7107;
      22747:data<=-16'd6557;
      22748:data<=-16'd6634;
      22749:data<=-16'd4899;
      22750:data<=-16'd884;
      22751:data<=16'd1333;
      22752:data<=16'd907;
      22753:data<=16'd958;
      22754:data<=16'd1148;
      22755:data<=16'd1268;
      22756:data<=16'd2246;
      22757:data<=16'd2388;
      22758:data<=16'd1800;
      22759:data<=16'd1836;
      22760:data<=16'd2673;
      22761:data<=16'd3617;
      22762:data<=16'd3231;
      22763:data<=16'd3726;
      22764:data<=16'd5630;
      22765:data<=16'd5573;
      22766:data<=16'd5705;
      22767:data<=16'd6575;
      22768:data<=16'd5742;
      22769:data<=16'd6096;
      22770:data<=16'd6816;
      22771:data<=16'd6194;
      22772:data<=16'd6816;
      22773:data<=16'd6942;
      22774:data<=16'd6754;
      22775:data<=16'd6946;
      22776:data<=16'd6200;
      22777:data<=16'd11973;
      22778:data<=16'd22789;
      22779:data<=16'd25364;
      22780:data<=16'd22952;
      22781:data<=16'd23102;
      22782:data<=16'd22592;
      22783:data<=16'd21828;
      22784:data<=16'd21610;
      22785:data<=16'd20172;
      22786:data<=16'd19188;
      22787:data<=16'd18800;
      22788:data<=16'd18842;
      22789:data<=16'd19951;
      22790:data<=16'd19886;
      22791:data<=16'd18389;
      22792:data<=16'd17643;
      22793:data<=16'd17566;
      22794:data<=16'd17114;
      22795:data<=16'd16392;
      22796:data<=16'd15820;
      22797:data<=16'd15323;
      22798:data<=16'd15076;
      22799:data<=16'd14512;
      22800:data<=16'd13338;
      22801:data<=16'd13737;
      22802:data<=16'd14722;
      22803:data<=16'd13670;
      22804:data<=16'd12915;
      22805:data<=16'd12871;
      22806:data<=16'd12057;
      22807:data<=16'd12090;
      22808:data<=16'd11981;
      22809:data<=16'd11028;
      22810:data<=16'd10866;
      22811:data<=16'd10358;
      22812:data<=16'd9796;
      22813:data<=16'd10022;
      22814:data<=16'd10342;
      22815:data<=16'd11048;
      22816:data<=16'd9429;
      22817:data<=16'd5695;
      22818:data<=16'd4701;
      22819:data<=16'd4808;
      22820:data<=16'd4225;
      22821:data<=16'd3976;
      22822:data<=16'd3030;
      22823:data<=16'd3372;
      22824:data<=16'd3507;
      22825:data<=16'd1892;
      22826:data<=16'd3720;
      22827:data<=16'd2076;
      22828:data<=-16'd8276;
      22829:data<=-16'd13051;
      22830:data<=-16'd10772;
      22831:data<=-16'd11227;
      22832:data<=-16'd11091;
      22833:data<=-16'd9803;
      22834:data<=-16'd10147;
      22835:data<=-16'd8933;
      22836:data<=-16'd7900;
      22837:data<=-16'd8493;
      22838:data<=-16'd7636;
      22839:data<=-16'd6115;
      22840:data<=-16'd5219;
      22841:data<=-16'd4654;
      22842:data<=-16'd4476;
      22843:data<=-16'd4475;
      22844:data<=-16'd4708;
      22845:data<=-16'd4485;
      22846:data<=-16'd4077;
      22847:data<=-16'd4206;
      22848:data<=-16'd3654;
      22849:data<=-16'd3247;
      22850:data<=-16'd3648;
      22851:data<=-16'd2667;
      22852:data<=-16'd807;
      22853:data<=-16'd83;
      22854:data<=-16'd414;
      22855:data<=-16'd701;
      22856:data<=-16'd356;
      22857:data<=-16'd252;
      22858:data<=-16'd447;
      22859:data<=-16'd277;
      22860:data<=16'd108;
      22861:data<=16'd447;
      22862:data<=-16'd378;
      22863:data<=-16'd879;
      22864:data<=16'd933;
      22865:data<=16'd1818;
      22866:data<=16'd1548;
      22867:data<=16'd2303;
      22868:data<=16'd2155;
      22869:data<=16'd1794;
      22870:data<=16'd1771;
      22871:data<=16'd1283;
      22872:data<=16'd2138;
      22873:data<=16'd2106;
      22874:data<=16'd1336;
      22875:data<=16'd2278;
      22876:data<=16'd1460;
      22877:data<=16'd4473;
      22878:data<=16'd14974;
      22879:data<=16'd19626;
      22880:data<=16'd17608;
      22881:data<=16'd17634;
      22882:data<=16'd16788;
      22883:data<=16'd16422;
      22884:data<=16'd18798;
      22885:data<=16'd18854;
      22886:data<=16'd17829;
      22887:data<=16'd17503;
      22888:data<=16'd16504;
      22889:data<=16'd16865;
      22890:data<=16'd17708;
      22891:data<=16'd16815;
      22892:data<=16'd15452;
      22893:data<=16'd14481;
      22894:data<=16'd13764;
      22895:data<=16'd12974;
      22896:data<=16'd12584;
      22897:data<=16'd12686;
      22898:data<=16'd11776;
      22899:data<=16'd10411;
      22900:data<=16'd9664;
      22901:data<=16'd9477;
      22902:data<=16'd10017;
      22903:data<=16'd9875;
      22904:data<=16'd9071;
      22905:data<=16'd8962;
      22906:data<=16'd8331;
      22907:data<=16'd7329;
      22908:data<=16'd6877;
      22909:data<=16'd6317;
      22910:data<=16'd6206;
      22911:data<=16'd6161;
      22912:data<=16'd5133;
      22913:data<=16'd4132;
      22914:data<=16'd4422;
      22915:data<=16'd5753;
      22916:data<=16'd5767;
      22917:data<=16'd4467;
      22918:data<=16'd4238;
      22919:data<=16'd3803;
      22920:data<=16'd3057;
      22921:data<=16'd3002;
      22922:data<=16'd1879;
      22923:data<=16'd1683;
      22924:data<=16'd2140;
      22925:data<=16'd188;
      22926:data<=16'd461;
      22927:data<=16'd679;
      22928:data<=-16'd6851;
      22929:data<=-16'd13888;
      22930:data<=-16'd13793;
      22931:data<=-16'd13382;
      22932:data<=-16'd13975;
      22933:data<=-16'd13251;
      22934:data<=-16'd12754;
      22935:data<=-16'd12492;
      22936:data<=-16'd12182;
      22937:data<=-16'd12120;
      22938:data<=-16'd11776;
      22939:data<=-16'd10963;
      22940:data<=-16'd9823;
      22941:data<=-16'd9253;
      22942:data<=-16'd9075;
      22943:data<=-16'd8305;
      22944:data<=-16'd8072;
      22945:data<=-16'd8329;
      22946:data<=-16'd8194;
      22947:data<=-16'd8557;
      22948:data<=-16'd8343;
      22949:data<=-16'd7459;
      22950:data<=-16'd8987;
      22951:data<=-16'd11579;
      22952:data<=-16'd11963;
      22953:data<=-16'd11523;
      22954:data<=-16'd11571;
      22955:data<=-16'd11485;
      22956:data<=-16'd11441;
      22957:data<=-16'd11177;
      22958:data<=-16'd10564;
      22959:data<=-16'd10348;
      22960:data<=-16'd10267;
      22961:data<=-16'd9984;
      22962:data<=-16'd9687;
      22963:data<=-16'd9417;
      22964:data<=-16'd10078;
      22965:data<=-16'd11348;
      22966:data<=-16'd11147;
      22967:data<=-16'd10276;
      22968:data<=-16'd10176;
      22969:data<=-16'd9665;
      22970:data<=-16'd9450;
      22971:data<=-16'd9702;
      22972:data<=-16'd8281;
      22973:data<=-16'd7887;
      22974:data<=-16'd9350;
      22975:data<=-16'd7900;
      22976:data<=-16'd7097;
      22977:data<=-16'd8990;
      22978:data<=-16'd3642;
      22979:data<=16'd5987;
      22980:data<=16'd7327;
      22981:data<=16'd5201;
      22982:data<=16'd6120;
      22983:data<=16'd5651;
      22984:data<=16'd4487;
      22985:data<=16'd4728;
      22986:data<=16'd4093;
      22987:data<=16'd3706;
      22988:data<=16'd4135;
      22989:data<=16'd3092;
      22990:data<=16'd1339;
      22991:data<=16'd845;
      22992:data<=16'd981;
      22993:data<=16'd517;
      22994:data<=16'd256;
      22995:data<=16'd629;
      22996:data<=16'd657;
      22997:data<=16'd754;
      22998:data<=16'd626;
      22999:data<=-16'd221;
      23000:data<=-16'd237;
      23001:data<=-16'd332;
      23002:data<=-16'd1630;
      23003:data<=-16'd2494;
      23004:data<=-16'd2867;
      23005:data<=-16'd2748;
      23006:data<=-16'd2273;
      23007:data<=-16'd2739;
      23008:data<=-16'd2877;
      23009:data<=-16'd2496;
      23010:data<=-16'd2911;
      23011:data<=-16'd3060;
      23012:data<=-16'd2893;
      23013:data<=-16'd2958;
      23014:data<=-16'd3457;
      23015:data<=-16'd4940;
      23016:data<=-16'd5482;
      23017:data<=-16'd3829;
      23018:data<=-16'd1368;
      23019:data<=16'd11;
      23020:data<=-16'd591;
      23021:data<=-16'd752;
      23022:data<=-16'd523;
      23023:data<=-16'd1401;
      23024:data<=-16'd792;
      23025:data<=-16'd829;
      23026:data<=-16'd2299;
      23027:data<=-16'd1977;
      23028:data<=-16'd7357;
      23029:data<=-16'd17793;
      23030:data<=-16'd19879;
      23031:data<=-16'd17311;
      23032:data<=-16'd17688;
      23033:data<=-16'd17256;
      23034:data<=-16'd16255;
      23035:data<=-16'd15549;
      23036:data<=-16'd14747;
      23037:data<=-16'd14960;
      23038:data<=-16'd14113;
      23039:data<=-16'd13775;
      23040:data<=-16'd15235;
      23041:data<=-16'd14883;
      23042:data<=-16'd14064;
      23043:data<=-16'd13794;
      23044:data<=-16'd12648;
      23045:data<=-16'd12425;
      23046:data<=-16'd12461;
      23047:data<=-16'd11925;
      23048:data<=-16'd11832;
      23049:data<=-16'd10868;
      23050:data<=-16'd9380;
      23051:data<=-16'd9098;
      23052:data<=-16'd10229;
      23053:data<=-16'd11415;
      23054:data<=-16'd10702;
      23055:data<=-16'd9556;
      23056:data<=-16'd9150;
      23057:data<=-16'd8624;
      23058:data<=-16'd8705;
      23059:data<=-16'd8243;
      23060:data<=-16'd7265;
      23061:data<=-16'd7709;
      23062:data<=-16'd7403;
      23063:data<=-16'd6228;
      23064:data<=-16'd6532;
      23065:data<=-16'd7620;
      23066:data<=-16'd8258;
      23067:data<=-16'd7292;
      23068:data<=-16'd6438;
      23069:data<=-16'd6965;
      23070:data<=-16'd6191;
      23071:data<=-16'd5686;
      23072:data<=-16'd5651;
      23073:data<=-16'd4150;
      23074:data<=-16'd4514;
      23075:data<=-16'd4158;
      23076:data<=-16'd2472;
      23077:data<=-16'd4555;
      23078:data<=-16'd1240;
      23079:data<=16'd9403;
      23080:data<=16'd12760;
      23081:data<=16'd10516;
      23082:data<=16'd10739;
      23083:data<=16'd10878;
      23084:data<=16'd9609;
      23085:data<=16'd6707;
      23086:data<=16'd4494;
      23087:data<=16'd5427;
      23088:data<=16'd5539;
      23089:data<=16'd4369;
      23090:data<=16'd3386;
      23091:data<=16'd2215;
      23092:data<=16'd2855;
      23093:data<=16'd3237;
      23094:data<=16'd2126;
      23095:data<=16'd2754;
      23096:data<=16'd3307;
      23097:data<=16'd2928;
      23098:data<=16'd3172;
      23099:data<=16'd2497;
      23100:data<=16'd2155;
      23101:data<=16'd2887;
      23102:data<=16'd2150;
      23103:data<=16'd652;
      23104:data<=16'd106;
      23105:data<=16'd365;
      23106:data<=16'd585;
      23107:data<=16'd506;
      23108:data<=16'd816;
      23109:data<=16'd1061;
      23110:data<=16'd1196;
      23111:data<=16'd1149;
      23112:data<=16'd661;
      23113:data<=16'd1510;
      23114:data<=16'd1782;
      23115:data<=-16'd422;
      23116:data<=-16'd1098;
      23117:data<=-16'd447;
      23118:data<=-16'd620;
      23119:data<=-16'd340;
      23120:data<=-16'd353;
      23121:data<=-16'd68;
      23122:data<=16'd358;
      23123:data<=-16'd596;
      23124:data<=-16'd202;
      23125:data<=16'd83;
      23126:data<=-16'd557;
      23127:data<=16'd402;
      23128:data<=-16'd4872;
      23129:data<=-16'd15740;
      23130:data<=-16'd18553;
      23131:data<=-16'd16043;
      23132:data<=-16'd15844;
      23133:data<=-16'd15432;
      23134:data<=-16'd14800;
      23135:data<=-16'd13847;
      23136:data<=-16'd12461;
      23137:data<=-16'd12372;
      23138:data<=-16'd11523;
      23139:data<=-16'd11089;
      23140:data<=-16'd12337;
      23141:data<=-16'd11928;
      23142:data<=-16'd11032;
      23143:data<=-16'd10580;
      23144:data<=-16'd9400;
      23145:data<=-16'd9180;
      23146:data<=-16'd9042;
      23147:data<=-16'd8316;
      23148:data<=-16'd7864;
      23149:data<=-16'd6749;
      23150:data<=-16'd6056;
      23151:data<=-16'd4696;
      23152:data<=-16'd1471;
      23153:data<=-16'd403;
      23154:data<=-16'd443;
      23155:data<=16'd948;
      23156:data<=16'd948;
      23157:data<=16'd508;
      23158:data<=16'd1127;
      23159:data<=16'd1139;
      23160:data<=16'd1260;
      23161:data<=16'd1847;
      23162:data<=16'd2191;
      23163:data<=16'd2406;
      23164:data<=16'd2990;
      23165:data<=16'd4614;
      23166:data<=16'd5439;
      23167:data<=16'd4786;
      23168:data<=16'd4927;
      23169:data<=16'd5503;
      23170:data<=16'd5642;
      23171:data<=16'd5524;
      23172:data<=16'd5480;
      23173:data<=16'd6161;
      23174:data<=16'd6270;
      23175:data<=16'd6496;
      23176:data<=16'd6824;
      23177:data<=16'd5641;
      23178:data<=16'd10557;
      23179:data<=16'd21814;
      23180:data<=16'd25401;
      23181:data<=16'd22660;
      23182:data<=16'd22297;
      23183:data<=16'd21842;
      23184:data<=16'd21413;
      23185:data<=16'd21241;
      23186:data<=16'd19785;
      23187:data<=16'd19792;
      23188:data<=16'd19417;
      23189:data<=16'd18322;
      23190:data<=16'd19517;
      23191:data<=16'd19488;
      23192:data<=16'd18207;
      23193:data<=16'd18221;
      23194:data<=16'd17327;
      23195:data<=16'd16519;
      23196:data<=16'd16512;
      23197:data<=16'd15943;
      23198:data<=16'd15731;
      23199:data<=16'd15053;
      23200:data<=16'd13893;
      23201:data<=16'd13430;
      23202:data<=16'd13405;
      23203:data<=16'd14249;
      23204:data<=16'd14140;
      23205:data<=16'd12684;
      23206:data<=16'd12549;
      23207:data<=16'd12516;
      23208:data<=16'd12151;
      23209:data<=16'd12105;
      23210:data<=16'd11147;
      23211:data<=16'd10819;
      23212:data<=16'd10705;
      23213:data<=16'd9617;
      23214:data<=16'd9832;
      23215:data<=16'd10282;
      23216:data<=16'd10480;
      23217:data<=16'd11107;
      23218:data<=16'd8969;
      23219:data<=16'd5429;
      23220:data<=16'd4264;
      23221:data<=16'd4422;
      23222:data<=16'd4290;
      23223:data<=16'd3664;
      23224:data<=16'd3659;
      23225:data<=16'd3479;
      23226:data<=16'd2851;
      23227:data<=16'd4736;
      23228:data<=16'd3057;
      23229:data<=-16'd6367;
      23230:data<=-16'd11911;
      23231:data<=-16'd10719;
      23232:data<=-16'd10451;
      23233:data<=-16'd10499;
      23234:data<=-16'd10161;
      23235:data<=-16'd10132;
      23236:data<=-16'd9188;
      23237:data<=-16'd8913;
      23238:data<=-16'd8733;
      23239:data<=-16'd7559;
      23240:data<=-16'd6485;
      23241:data<=-16'd5156;
      23242:data<=-16'd4778;
      23243:data<=-16'd5083;
      23244:data<=-16'd4269;
      23245:data<=-16'd4196;
      23246:data<=-16'd4573;
      23247:data<=-16'd4276;
      23248:data<=-16'd4431;
      23249:data<=-16'd3797;
      23250:data<=-16'd2830;
      23251:data<=-16'd2951;
      23252:data<=-16'd2147;
      23253:data<=-16'd391;
      23254:data<=16'd453;
      23255:data<=16'd246;
      23256:data<=16'd12;
      23257:data<=16'd255;
      23258:data<=-16'd297;
      23259:data<=-16'd1007;
      23260:data<=-16'd476;
      23261:data<=16'd36;
      23262:data<=16'd423;
      23263:data<=16'd482;
      23264:data<=16'd89;
      23265:data<=16'd1292;
      23266:data<=16'd2570;
      23267:data<=16'd2294;
      23268:data<=16'd2406;
      23269:data<=16'd2682;
      23270:data<=16'd2769;
      23271:data<=16'd2576;
      23272:data<=16'd1727;
      23273:data<=16'd2093;
      23274:data<=16'd2463;
      23275:data<=16'd1903;
      23276:data<=16'd2353;
      23277:data<=16'd2021;
      23278:data<=16'd4347;
      23279:data<=16'd13552;
      23280:data<=16'd19649;
      23281:data<=16'd18328;
      23282:data<=16'd17872;
      23283:data<=16'd18017;
      23284:data<=16'd16477;
      23285:data<=16'd17302;
      23286:data<=16'd19264;
      23287:data<=16'd18929;
      23288:data<=16'd17773;
      23289:data<=16'd17267;
      23290:data<=16'd17294;
      23291:data<=16'd17493;
      23292:data<=16'd16822;
      23293:data<=16'd15470;
      23294:data<=16'd14906;
      23295:data<=16'd14654;
      23296:data<=16'd13659;
      23297:data<=16'd12736;
      23298:data<=16'd12187;
      23299:data<=16'd11721;
      23300:data<=16'd11104;
      23301:data<=16'd9599;
      23302:data<=16'd9071;
      23303:data<=16'd10816;
      23304:data<=16'd11371;
      23305:data<=16'd9840;
      23306:data<=16'd9010;
      23307:data<=16'd8898;
      23308:data<=16'd8411;
      23309:data<=16'd7670;
      23310:data<=16'd7130;
      23311:data<=16'd6792;
      23312:data<=16'd6075;
      23313:data<=16'd5506;
      23314:data<=16'd5083;
      23315:data<=16'd4642;
      23316:data<=16'd5611;
      23317:data<=16'd6203;
      23318:data<=16'd4927;
      23319:data<=16'd4438;
      23320:data<=16'd3987;
      23321:data<=16'd3107;
      23322:data<=16'd3703;
      23323:data<=16'd3063;
      23324:data<=16'd1624;
      23325:data<=16'd1797;
      23326:data<=16'd978;
      23327:data<=16'd1694;
      23328:data<=16'd3156;
      23329:data<=-16'd3698;
      23330:data<=-16'd12839;
      23331:data<=-16'd13723;
      23332:data<=-16'd12434;
      23333:data<=-16'd13110;
      23334:data<=-16'd12627;
      23335:data<=-16'd12361;
      23336:data<=-16'd12542;
      23337:data<=-16'd11829;
      23338:data<=-16'd11479;
      23339:data<=-16'd11358;
      23340:data<=-16'd10419;
      23341:data<=-16'd8874;
      23342:data<=-16'd7935;
      23343:data<=-16'd8329;
      23344:data<=-16'd8551;
      23345:data<=-16'd8017;
      23346:data<=-16'd7809;
      23347:data<=-16'd7615;
      23348:data<=-16'd7289;
      23349:data<=-16'd7498;
      23350:data<=-16'd7556;
      23351:data<=-16'd7083;
      23352:data<=-16'd8102;
      23353:data<=-16'd10806;
      23354:data<=-16'd11486;
      23355:data<=-16'd10097;
      23356:data<=-16'd9991;
      23357:data<=-16'd10332;
      23358:data<=-16'd10107;
      23359:data<=-16'd9982;
      23360:data<=-16'd9112;
      23361:data<=-16'd8671;
      23362:data<=-16'd9059;
      23363:data<=-16'd8404;
      23364:data<=-16'd8150;
      23365:data<=-16'd8942;
      23366:data<=-16'd9371;
      23367:data<=-16'd9588;
      23368:data<=-16'd9206;
      23369:data<=-16'd8845;
      23370:data<=-16'd8874;
      23371:data<=-16'd8513;
      23372:data<=-16'd8940;
      23373:data<=-16'd8577;
      23374:data<=-16'd7253;
      23375:data<=-16'd7990;
      23376:data<=-16'd7445;
      23377:data<=-16'd7150;
      23378:data<=-16'd10169;
      23379:data<=-16'd5250;
      23380:data<=16'd6003;
      23381:data<=16'd8009;
      23382:data<=16'd5574;
      23383:data<=16'd6617;
      23384:data<=16'd6505;
      23385:data<=16'd6026;
      23386:data<=16'd6206;
      23387:data<=16'd4974;
      23388:data<=16'd4349;
      23389:data<=16'd4074;
      23390:data<=16'd2880;
      23391:data<=16'd1765;
      23392:data<=16'd1130;
      23393:data<=16'd1219;
      23394:data<=16'd1095;
      23395:data<=16'd849;
      23396:data<=16'd1033;
      23397:data<=-16'd61;
      23398:data<=-16'd828;
      23399:data<=-16'd21;
      23400:data<=-16'd205;
      23401:data<=-16'd531;
      23402:data<=-16'd588;
      23403:data<=-16'd1933;
      23404:data<=-16'd2804;
      23405:data<=-16'd2784;
      23406:data<=-16'd3203;
      23407:data<=-16'd3544;
      23408:data<=-16'd3165;
      23409:data<=-16'd2455;
      23410:data<=-16'd2757;
      23411:data<=-16'd3474;
      23412:data<=-16'd3466;
      23413:data<=-16'd3472;
      23414:data<=-16'd2830;
      23415:data<=-16'd2925;
      23416:data<=-16'd5104;
      23417:data<=-16'd5814;
      23418:data<=-16'd5209;
      23419:data<=-16'd4053;
      23420:data<=-16'd1146;
      23421:data<=-16'd381;
      23422:data<=-16'd1130;
      23423:data<=-16'd619;
      23424:data<=-16'd1466;
      23425:data<=-16'd1850;
      23426:data<=-16'd1895;
      23427:data<=-16'd2804;
      23428:data<=-16'd1721;
      23429:data<=-16'd6690;
      23430:data<=-16'd18063;
      23431:data<=-16'd20703;
      23432:data<=-16'd17887;
      23433:data<=-16'd18073;
      23434:data<=-16'd17059;
      23435:data<=-16'd16486;
      23436:data<=-16'd16962;
      23437:data<=-16'd15561;
      23438:data<=-16'd14994;
      23439:data<=-16'd14697;
      23440:data<=-16'd14363;
      23441:data<=-16'd15256;
      23442:data<=-16'd14774;
      23443:data<=-16'd13975;
      23444:data<=-16'd13951;
      23445:data<=-16'd13241;
      23446:data<=-16'd12599;
      23447:data<=-16'd11350;
      23448:data<=-16'd10478;
      23449:data<=-16'd11300;
      23450:data<=-16'd11162;
      23451:data<=-16'd10176;
      23452:data<=-16'd9609;
      23453:data<=-16'd10013;
      23454:data<=-16'd11644;
      23455:data<=-16'd11239;
      23456:data<=-16'd9529;
      23457:data<=-16'd9482;
      23458:data<=-16'd9303;
      23459:data<=-16'd8962;
      23460:data<=-16'd8434;
      23461:data<=-16'd7254;
      23462:data<=-16'd7457;
      23463:data<=-16'd7304;
      23464:data<=-16'd6049;
      23465:data<=-16'd6173;
      23466:data<=-16'd6990;
      23467:data<=-16'd7621;
      23468:data<=-16'd7165;
      23469:data<=-16'd6291;
      23470:data<=-16'd6551;
      23471:data<=-16'd5460;
      23472:data<=-16'd4543;
      23473:data<=-16'd5321;
      23474:data<=-16'd4602;
      23475:data<=-16'd4444;
      23476:data<=-16'd3635;
      23477:data<=-16'd1723;
      23478:data<=-16'd4428;
      23479:data<=-16'd2130;
      23480:data<=16'd8947;
      23481:data<=16'd12378;
      23482:data<=16'd9969;
      23483:data<=16'd11009;
      23484:data<=16'd10731;
      23485:data<=16'd10219;
      23486:data<=16'd9661;
      23487:data<=16'd5897;
      23488:data<=16'd4579;
      23489:data<=16'd5570;
      23490:data<=16'd4400;
      23491:data<=16'd2958;
      23492:data<=16'd2159;
      23493:data<=16'd2361;
      23494:data<=16'd3042;
      23495:data<=16'd2538;
      23496:data<=16'd2514;
      23497:data<=16'd2775;
      23498:data<=16'd2425;
      23499:data<=16'd2728;
      23500:data<=16'd2496;
      23501:data<=16'd1868;
      23502:data<=16'd2250;
      23503:data<=16'd1727;
      23504:data<=16'd194;
      23505:data<=-16'd126;
      23506:data<=16'd165;
      23507:data<=-16'd270;
      23508:data<=-16'd265;
      23509:data<=16'd384;
      23510:data<=16'd162;
      23511:data<=16'd120;
      23512:data<=16'd599;
      23513:data<=16'd464;
      23514:data<=16'd1134;
      23515:data<=16'd1087;
      23516:data<=-16'd1127;
      23517:data<=-16'd1598;
      23518:data<=-16'd643;
      23519:data<=-16'd663;
      23520:data<=-16'd708;
      23521:data<=-16'd948;
      23522:data<=-16'd652;
      23523:data<=-16'd396;
      23524:data<=-16'd998;
      23525:data<=-16'd62;
      23526:data<=-16'd411;
      23527:data<=-16'd1638;
      23528:data<=16'd35;
      23529:data<=-16'd4723;
      23530:data<=-16'd15705;
      23531:data<=-16'd18445;
      23532:data<=-16'd16301;
      23533:data<=-16'd16545;
      23534:data<=-16'd15661;
      23535:data<=-16'd15089;
      23536:data<=-16'd15001;
      23537:data<=-16'd13389;
      23538:data<=-16'd12645;
      23539:data<=-16'd11782;
      23540:data<=-16'd11045;
      23541:data<=-16'd11866;
      23542:data<=-16'd11297;
      23543:data<=-16'd10443;
      23544:data<=-16'd10769;
      23545:data<=-16'd10067;
      23546:data<=-16'd9313;
      23547:data<=-16'd8718;
      23548:data<=-16'd7677;
      23549:data<=-16'd7412;
      23550:data<=-16'd6689;
      23551:data<=-16'd5686;
      23552:data<=-16'd5309;
      23553:data<=-16'd2972;
      23554:data<=16'd253;
      23555:data<=16'd1195;
      23556:data<=16'd1415;
      23557:data<=16'd1903;
      23558:data<=16'd1424;
      23559:data<=16'd1202;
      23560:data<=16'd2149;
      23561:data<=16'd2555;
      23562:data<=16'd2394;
      23563:data<=16'd2467;
      23564:data<=16'd2194;
      23565:data<=16'd2990;
      23566:data<=16'd5103;
      23567:data<=16'd5671;
      23568:data<=16'd5344;
      23569:data<=16'd5607;
      23570:data<=16'd5806;
      23571:data<=16'd6410;
      23572:data<=16'd6537;
      23573:data<=16'd6228;
      23574:data<=16'd6746;
      23575:data<=16'd6443;
      23576:data<=16'd6687;
      23577:data<=16'd7459;
      23578:data<=16'd6216;
      23579:data<=16'd10508;
      23580:data<=16'd21033;
      23581:data<=16'd24891;
      23582:data<=16'd23244;
      23583:data<=16'd23282;
      23584:data<=16'd22441;
      23585:data<=16'd21614;
      23586:data<=16'd21620;
      23587:data<=16'd20239;
      23588:data<=16'd19341;
      23589:data<=16'd18375;
      23590:data<=16'd17403;
      23591:data<=16'd18726;
      23592:data<=16'd19109;
      23593:data<=16'd17916;
      23594:data<=16'd17908;
      23595:data<=16'd17760;
      23596:data<=16'd17124;
      23597:data<=16'd16496;
      23598:data<=16'd15476;
      23599:data<=16'd14854;
      23600:data<=16'd14084;
      23601:data<=16'd13103;
      23602:data<=16'd12713;
      23603:data<=16'd12646;
      23604:data<=16'd13370;
      23605:data<=16'd13591;
      23606:data<=16'd12328;
      23607:data<=16'd11972;
      23608:data<=16'd12292;
      23609:data<=16'd11925;
      23610:data<=16'd11670;
      23611:data<=16'd11163;
      23612:data<=16'd10396;
      23613:data<=16'd9844;
      23614:data<=16'd9113;
      23615:data<=16'd8975;
      23616:data<=16'd9811;
      23617:data<=16'd10473;
      23618:data<=16'd10326;
      23619:data<=16'd9730;
      23620:data<=16'd8067;
      23621:data<=16'd4907;
      23622:data<=16'd3686;
      23623:data<=16'd4807;
      23624:data<=16'd4285;
      23625:data<=16'd3987;
      23626:data<=16'd4475;
      23627:data<=16'd3371;
      23628:data<=16'd4399;
      23629:data<=16'd3809;
      23630:data<=-16'd4451;
      23631:data<=-16'd10611;
      23632:data<=-16'd10264;
      23633:data<=-16'd10539;
      23634:data<=-16'd11042;
      23635:data<=-16'd10290;
      23636:data<=-16'd9718;
      23637:data<=-16'd8669;
      23638:data<=-16'd7979;
      23639:data<=-16'd7498;
      23640:data<=-16'd6790;
      23641:data<=-16'd6349;
      23642:data<=-16'd4831;
      23643:data<=-16'd4002;
      23644:data<=-16'd4695;
      23645:data<=-16'd3908;
      23646:data<=-16'd3330;
      23647:data<=-16'd3965;
      23648:data<=-16'd3489;
      23649:data<=-16'd3054;
      23650:data<=-16'd2673;
      23651:data<=-16'd1680;
      23652:data<=-16'd1670;
      23653:data<=-16'd1300;
      23654:data<=16'd487;
      23655:data<=16'd1713;
      23656:data<=16'd1780;
      23657:data<=16'd1310;
      23658:data<=16'd723;
      23659:data<=16'd408;
      23660:data<=16'd911;
      23661:data<=16'd1530;
      23662:data<=16'd864;
      23663:data<=16'd793;
      23664:data<=16'd1686;
      23665:data<=16'd860;
      23666:data<=16'd687;
      23667:data<=16'd2717;
      23668:data<=16'd3380;
      23669:data<=16'd2843;
      23670:data<=16'd2672;
      23671:data<=16'd2481;
      23672:data<=16'd2661;
      23673:data<=16'd2522;
      23674:data<=16'd2158;
      23675:data<=16'd2284;
      23676:data<=16'd2174;
      23677:data<=16'd2250;
      23678:data<=16'd1874;
      23679:data<=16'd3227;
      23680:data<=16'd11314;
      23681:data<=16'd19435;
      23682:data<=16'd19594;
      23683:data<=16'd17734;
      23684:data<=16'd17541;
      23685:data<=16'd16595;
      23686:data<=16'd16434;
      23687:data<=16'd17632;
      23688:data<=16'd18616;
      23689:data<=16'd17998;
      23690:data<=16'd15869;
      23691:data<=16'd15779;
      23692:data<=16'd17150;
      23693:data<=16'd16625;
      23694:data<=16'd15646;
      23695:data<=16'd14574;
      23696:data<=16'd13394;
      23697:data<=16'd13637;
      23698:data<=16'd13062;
      23699:data<=16'd11556;
      23700:data<=16'd11309;
      23701:data<=16'd10571;
      23702:data<=16'd9206;
      23703:data<=16'd8795;
      23704:data<=16'd9112;
      23705:data<=16'd9693;
      23706:data<=16'd9145;
      23707:data<=16'd8067;
      23708:data<=16'd7840;
      23709:data<=16'd6865;
      23710:data<=16'd6034;
      23711:data<=16'd6495;
      23712:data<=16'd6106;
      23713:data<=16'd5479;
      23714:data<=16'd5409;
      23715:data<=16'd4634;
      23716:data<=16'd4399;
      23717:data<=16'd5607;
      23718:data<=16'd6229;
      23719:data<=16'd5127;
      23720:data<=16'd4037;
      23721:data<=16'd3788;
      23722:data<=16'd3121;
      23723:data<=16'd2698;
      23724:data<=16'd2594;
      23725:data<=16'd2290;
      23726:data<=16'd2837;
      23727:data<=16'd1804;
      23728:data<=16'd873;
      23729:data<=16'd3526;
      23730:data<=-16'd158;
      23731:data<=-16'd10960;
      23732:data<=-16'd14214;
      23733:data<=-16'd11914;
      23734:data<=-16'd11684;
      23735:data<=-16'd10448;
      23736:data<=-16'd9755;
      23737:data<=-16'd10386;
      23738:data<=-16'd9420;
      23739:data<=-16'd8851;
      23740:data<=-16'd8854;
      23741:data<=-16'd8234;
      23742:data<=-16'd7200;
      23743:data<=-16'd5946;
      23744:data<=-16'd6273;
      23745:data<=-16'd6696;
      23746:data<=-16'd5927;
      23747:data<=-16'd6343;
      23748:data<=-16'd6660;
      23749:data<=-16'd6176;
      23750:data<=-16'd6058;
      23751:data<=-16'd5432;
      23752:data<=-16'd5213;
      23753:data<=-16'd5718;
      23754:data<=-16'd6990;
      23755:data<=-16'd8950;
      23756:data<=-16'd8578;
      23757:data<=-16'd7777;
      23758:data<=-16'd8533;
      23759:data<=-16'd7897;
      23760:data<=-16'd7861;
      23761:data<=-16'd8715;
      23762:data<=-16'd8019;
      23763:data<=-16'd8234;
      23764:data<=-16'd8176;
      23765:data<=-16'd6975;
      23766:data<=-16'd7835;
      23767:data<=-16'd9022;
      23768:data<=-16'd9203;
      23769:data<=-16'd9250;
      23770:data<=-16'd9036;
      23771:data<=-16'd9185;
      23772:data<=-16'd8702;
      23773:data<=-16'd8493;
      23774:data<=-16'd9115;
      23775:data<=-16'd8429;
      23776:data<=-16'd8260;
      23777:data<=-16'd7524;
      23778:data<=-16'd6721;
      23779:data<=-16'd9987;
      23780:data<=-16'd7309;
      23781:data<=16'd2966;
      23782:data<=16'd5288;
      23783:data<=16'd3242;
      23784:data<=16'd4720;
      23785:data<=16'd3865;
      23786:data<=16'd2975;
      23787:data<=16'd3845;
      23788:data<=16'd2626;
      23789:data<=16'd2087;
      23790:data<=16'd2247;
      23791:data<=16'd1040;
      23792:data<=-16'd156;
      23793:data<=-16'd1049;
      23794:data<=-16'd760;
      23795:data<=-16'd349;
      23796:data<=-16'd1316;
      23797:data<=-16'd1644;
      23798:data<=-16'd1565;
      23799:data<=-16'd1853;
      23800:data<=-16'd1915;
      23801:data<=-16'd2000;
      23802:data<=-16'd1792;
      23803:data<=-16'd2751;
      23804:data<=-16'd4775;
      23805:data<=-16'd5134;
      23806:data<=-16'd5116;
      23807:data<=-16'd5395;
      23808:data<=-16'd4821;
      23809:data<=-16'd4679;
      23810:data<=-16'd4748;
      23811:data<=-16'd4498;
      23812:data<=-16'd4473;
      23813:data<=-16'd4473;
      23814:data<=-16'd4487;
      23815:data<=-16'd3940;
      23816:data<=-16'd4296;
      23817:data<=-16'd6182;
      23818:data<=-16'd6347;
      23819:data<=-16'd5868;
      23820:data<=-16'd5567;
      23821:data<=-16'd3196;
      23822:data<=-16'd1724;
      23823:data<=-16'd1713;
      23824:data<=-16'd1262;
      23825:data<=-16'd1730;
      23826:data<=-16'd1528;
      23827:data<=-16'd1525;
      23828:data<=-16'd2523;
      23829:data<=-16'd1626;
      23830:data<=-16'd5632;
      23831:data<=-16'd15159;
      23832:data<=-16'd17555;
      23833:data<=-16'd15086;
      23834:data<=-16'd15352;
      23835:data<=-16'd15077;
      23836:data<=-16'd14483;
      23837:data<=-16'd14581;
      23838:data<=-16'd13722;
      23839:data<=-16'd13101;
      23840:data<=-16'd12098;
      23841:data<=-16'd11491;
      23842:data<=-16'd12941;
      23843:data<=-16'd13406;
      23844:data<=-16'd12562;
      23845:data<=-16'd12049;
      23846:data<=-16'd10997;
      23847:data<=-16'd10395;
      23848:data<=-16'd10489;
      23849:data<=-16'd9609;
      23850:data<=-16'd8762;
      23851:data<=-16'd9001;
      23852:data<=-16'd8669;
      23853:data<=-16'd7409;
      23854:data<=-16'd7594;
      23855:data<=-16'd8853;
      23856:data<=-16'd8705;
      23857:data<=-16'd8357;
      23858:data<=-16'd8549;
      23859:data<=-16'd8000;
      23860:data<=-16'd7837;
      23861:data<=-16'd7862;
      23862:data<=-16'd6840;
      23863:data<=-16'd6232;
      23864:data<=-16'd6216;
      23865:data<=-16'd5896;
      23866:data<=-16'd6068;
      23867:data<=-16'd7156;
      23868:data<=-16'd7856;
      23869:data<=-16'd7087;
      23870:data<=-16'd6460;
      23871:data<=-16'd6220;
      23872:data<=-16'd4963;
      23873:data<=-16'd4993;
      23874:data<=-16'd5629;
      23875:data<=-16'd4394;
      23876:data<=-16'd4437;
      23877:data<=-16'd4331;
      23878:data<=-16'd3162;
      23879:data<=-16'd5439;
      23880:data<=-16'd3485;
      23881:data<=16'd5832;
      23882:data<=16'd8969;
      23883:data<=16'd7156;
      23884:data<=16'd8514;
      23885:data<=16'd8094;
      23886:data<=16'd6933;
      23887:data<=16'd7368;
      23888:data<=16'd4634;
      23889:data<=16'd2088;
      23890:data<=16'd2444;
      23891:data<=16'd1666;
      23892:data<=16'd538;
      23893:data<=16'd293;
      23894:data<=16'd277;
      23895:data<=16'd743;
      23896:data<=16'd543;
      23897:data<=16'd268;
      23898:data<=16'd525;
      23899:data<=16'd177;
      23900:data<=16'd86;
      23901:data<=16'd73;
      23902:data<=16'd30;
      23903:data<=16'd879;
      23904:data<=16'd147;
      23905:data<=-16'd1820;
      23906:data<=-16'd1745;
      23907:data<=-16'd1245;
      23908:data<=-16'd1368;
      23909:data<=-16'd875;
      23910:data<=-16'd647;
      23911:data<=-16'd388;
      23912:data<=16'd244;
      23913:data<=-16'd55;
      23914:data<=-16'd246;
      23915:data<=16'd379;
      23916:data<=-16'd6;
      23917:data<=-16'd1113;
      23918:data<=-16'd1389;
      23919:data<=-16'd1359;
      23920:data<=-16'd1310;
      23921:data<=-16'd1124;
      23922:data<=-16'd1287;
      23923:data<=-16'd829;
      23924:data<=16'd61;
      23925:data<=-16'd126;
      23926:data<=-16'd288;
      23927:data<=-16'd563;
      23928:data<=-16'd702;
      23929:data<=16'd629;
      23930:data<=-16'd2972;
      23931:data<=-16'd12317;
      23932:data<=-16'd15685;
      23933:data<=-16'd13336;
      23934:data<=-16'd13051;
      23935:data<=-16'd12610;
      23936:data<=-16'd11547;
      23937:data<=-16'd11476;
      23938:data<=-16'd10734;
      23939:data<=-16'd10470;
      23940:data<=-16'd10082;
      23941:data<=-16'd8801;
      23942:data<=-16'd9033;
      23943:data<=-16'd9454;
      23944:data<=-16'd9201;
      23945:data<=-16'd8922;
      23946:data<=-16'd7488;
      23947:data<=-16'd6678;
      23948:data<=-16'd6686;
      23949:data<=-16'd5735;
      23950:data<=-16'd5382;
      23951:data<=-16'd5093;
      23952:data<=-16'd4441;
      23953:data<=-16'd4676;
      23954:data<=-16'd3424;
      23955:data<=-16'd610;
      23956:data<=16'd1092;
      23957:data<=16'd1730;
      23958:data<=16'd1547;
      23959:data<=16'd1330;
      23960:data<=16'd1662;
      23961:data<=16'd1607;
      23962:data<=16'd1706;
      23963:data<=16'd2187;
      23964:data<=16'd2381;
      23965:data<=16'd2408;
      23966:data<=16'd2729;
      23967:data<=16'd3956;
      23968:data<=16'd4993;
      23969:data<=16'd5225;
      23970:data<=16'd5639;
      23971:data<=16'd5450;
      23972:data<=16'd5134;
      23973:data<=16'd5224;
      23974:data<=16'd4608;
      23975:data<=16'd4899;
      23976:data<=16'd5633;
      23977:data<=16'd5460;
      23978:data<=16'd5717;
      23979:data<=16'd5148;
      23980:data<=16'd7512;
      23981:data<=16'd16073;
      23982:data<=16'd20971;
      23983:data<=16'd19930;
      23984:data<=16'd20033;
      23985:data<=16'd19361;
      23986:data<=16'd17798;
      23987:data<=16'd17958;
      23988:data<=16'd17390;
      23989:data<=16'd16760;
      23990:data<=16'd16296;
      23991:data<=16'd15032;
      23992:data<=16'd15490;
      23993:data<=16'd16384;
      23994:data<=16'd15973;
      23995:data<=16'd15779;
      23996:data<=16'd15159;
      23997:data<=16'd14393;
      23998:data<=16'd14287;
      23999:data<=16'd13665;
      24000:data<=16'd12745;
      24001:data<=16'd12276;
      24002:data<=16'd12216;
      24003:data<=16'd11817;
      24004:data<=16'd11291;
      24005:data<=16'd12146;
      24006:data<=16'd12557;
      24007:data<=16'd11449;
      24008:data<=16'd11247;
      24009:data<=16'd11157;
      24010:data<=16'd10558;
      24011:data<=16'd10742;
      24012:data<=16'd10340;
      24013:data<=16'd9597;
      24014:data<=16'd9570;
      24015:data<=16'd8781;
      24016:data<=16'd7962;
      24017:data<=16'd8896;
      24018:data<=16'd10143;
      24019:data<=16'd9796;
      24020:data<=16'd8943;
      24021:data<=16'd8257;
      24022:data<=16'd5977;
      24023:data<=16'd4129;
      24024:data<=16'd4676;
      24025:data<=16'd4360;
      24026:data<=16'd3858;
      24027:data<=16'd4003;
      24028:data<=16'd2464;
      24029:data<=16'd3410;
      24030:data<=16'd5078;
      24031:data<=-16'd1151;
      24032:data<=-16'd8382;
      24033:data<=-16'd8464;
      24034:data<=-16'd7608;
      24035:data<=-16'd8085;
      24036:data<=-16'd7257;
      24037:data<=-16'd6736;
      24038:data<=-16'd6783;
      24039:data<=-16'd6407;
      24040:data<=-16'd6008;
      24041:data<=-16'd5635;
      24042:data<=-16'd4842;
      24043:data<=-16'd3404;
      24044:data<=-16'd2584;
      24045:data<=-16'd2811;
      24046:data<=-16'd2667;
      24047:data<=-16'd2467;
      24048:data<=-16'd2525;
      24049:data<=-16'd2341;
      24050:data<=-16'd2212;
      24051:data<=-16'd1516;
      24052:data<=-16'd1080;
      24053:data<=-16'd1886;
      24054:data<=-16'd1236;
      24055:data<=16'd795;
      24056:data<=16'd1501;
      24057:data<=16'd1685;
      24058:data<=16'd1633;
      24059:data<=16'd820;
      24060:data<=16'd690;
      24061:data<=16'd1233;
      24062:data<=16'd1219;
      24063:data<=16'd807;
      24064:data<=16'd925;
      24065:data<=16'd1300;
      24066:data<=16'd1078;
      24067:data<=16'd1527;
      24068:data<=16'd2461;
      24069:data<=16'd2361;
      24070:data<=16'd2878;
      24071:data<=16'd3295;
      24072:data<=16'd2187;
      24073:data<=16'd2111;
      24074:data<=16'd2105;
      24075:data<=16'd1509;
      24076:data<=16'd2322;
      24077:data<=16'd2224;
      24078:data<=16'd1818;
      24079:data<=16'd2323;
      24080:data<=16'd2244;
      24081:data<=16'd7427;
      24082:data<=16'd16281;
      24083:data<=16'd17546;
      24084:data<=16'd14995;
      24085:data<=16'd15473;
      24086:data<=16'd15159;
      24087:data<=16'd13896;
      24088:data<=16'd14122;
      24089:data<=16'd15546;
      24090:data<=16'd16551;
      24091:data<=16'd15549;
      24092:data<=16'd15164;
      24093:data<=16'd15763;
      24094:data<=16'd14945;
      24095:data<=16'd14571;
      24096:data<=16'd13963;
      24097:data<=16'd12299;
      24098:data<=16'd12437;
      24099:data<=16'd12340;
      24100:data<=16'd10634;
      24101:data<=16'd10022;
      24102:data<=16'd9953;
      24103:data<=16'd9464;
      24104:data<=16'd9110;
      24105:data<=16'd9312;
      24106:data<=16'd9690;
      24107:data<=16'd9047;
      24108:data<=16'd8663;
      24109:data<=16'd8854;
      24110:data<=16'd8035;
      24111:data<=16'd7383;
      24112:data<=16'd6717;
      24113:data<=16'd5659;
      24114:data<=16'd5691;
      24115:data<=16'd5319;
      24116:data<=16'd4610;
      24117:data<=16'd5353;
      24118:data<=16'd6249;
      24119:data<=16'd6335;
      24120:data<=16'd5303;
      24121:data<=16'd4258;
      24122:data<=16'd4422;
      24123:data<=16'd4020;
      24124:data<=16'd3576;
      24125:data<=16'd3257;
      24126:data<=16'd2319;
      24127:data<=16'd3055;
      24128:data<=16'd2657;
      24129:data<=16'd1421;
      24130:data<=16'd4108;
      24131:data<=16'd1445;
      24132:data<=-16'd8580;
      24133:data<=-16'd11546;
      24134:data<=-16'd9458;
      24135:data<=-16'd10386;
      24136:data<=-16'd10378;
      24137:data<=-16'd9703;
      24138:data<=-16'd9940;
      24139:data<=-16'd9226;
      24140:data<=-16'd9145;
      24141:data<=-16'd9227;
      24142:data<=-16'd7946;
      24143:data<=-16'd6570;
      24144:data<=-16'd5873;
      24145:data<=-16'd6231;
      24146:data<=-16'd6623;
      24147:data<=-16'd6100;
      24148:data<=-16'd5703;
      24149:data<=-16'd5651;
      24150:data<=-16'd5833;
      24151:data<=-16'd5826;
      24152:data<=-16'd5642;
      24153:data<=-16'd5999;
      24154:data<=-16'd5736;
      24155:data<=-16'd6149;
      24156:data<=-16'd8572;
      24157:data<=-16'd9277;
      24158:data<=-16'd8545;
      24159:data<=-16'd8989;
      24160:data<=-16'd8971;
      24161:data<=-16'd8668;
      24162:data<=-16'd8495;
      24163:data<=-16'd7915;
      24164:data<=-16'd8170;
      24165:data<=-16'd8099;
      24166:data<=-16'd7412;
      24167:data<=-16'd8225;
      24168:data<=-16'd9797;
      24169:data<=-16'd10426;
      24170:data<=-16'd9414;
      24171:data<=-16'd8461;
      24172:data<=-16'd8951;
      24173:data<=-16'd8702;
      24174:data<=-16'd8616;
      24175:data<=-16'd8978;
      24176:data<=-16'd7797;
      24177:data<=-16'd7987;
      24178:data<=-16'd7909;
      24179:data<=-16'd6673;
      24180:data<=-16'd9465;
      24181:data<=-16'd7477;
      24182:data<=16'd2778;
      24183:data<=16'd5535;
      24184:data<=16'd2429;
      24185:data<=16'd3636;
      24186:data<=16'd3792;
      24187:data<=16'd2491;
      24188:data<=16'd3113;
      24189:data<=16'd2902;
      24190:data<=16'd2561;
      24191:data<=16'd2648;
      24192:data<=16'd1607;
      24193:data<=-16'd187;
      24194:data<=-16'd1439;
      24195:data<=-16'd708;
      24196:data<=-16'd203;
      24197:data<=-16'd1201;
      24198:data<=-16'd1356;
      24199:data<=-16'd1536;
      24200:data<=-16'd1392;
      24201:data<=-16'd394;
      24202:data<=-16'd1263;
      24203:data<=-16'd1723;
      24204:data<=-16'd652;
      24205:data<=-16'd1459;
      24206:data<=-16'd2857;
      24207:data<=-16'd3554;
      24208:data<=-16'd4222;
      24209:data<=-16'd4030;
      24210:data<=-16'd3580;
      24211:data<=-16'd3519;
      24212:data<=-16'd3821;
      24213:data<=-16'd3838;
      24214:data<=-16'd3213;
      24215:data<=-16'd3486;
      24216:data<=-16'd3259;
      24217:data<=-16'd2496;
      24218:data<=-16'd4059;
      24219:data<=-16'd5013;
      24220:data<=-16'd4761;
      24221:data<=-16'd5755;
      24222:data<=-16'd4601;
      24223:data<=-16'd1713;
      24224:data<=-16'd526;
      24225:data<=-16'd405;
      24226:data<=-16'd863;
      24227:data<=-16'd693;
      24228:data<=-16'd784;
      24229:data<=-16'd1313;
      24230:data<=-16'd106;
      24231:data<=-16'd4356;
      24232:data<=-16'd14492;
      24233:data<=-16'd17388;
      24234:data<=-16'd14963;
      24235:data<=-16'd14973;
      24236:data<=-16'd14251;
      24237:data<=-16'd13353;
      24238:data<=-16'd13464;
      24239:data<=-16'd12737;
      24240:data<=-16'd12525;
      24241:data<=-16'd12055;
      24242:data<=-16'd11389;
      24243:data<=-16'd12151;
      24244:data<=-16'd12323;
      24245:data<=-16'd11899;
      24246:data<=-16'd11756;
      24247:data<=-16'd10837;
      24248:data<=-16'd9881;
      24249:data<=-16'd9500;
      24250:data<=-16'd9312;
      24251:data<=-16'd9009;
      24252:data<=-16'd8722;
      24253:data<=-16'd8514;
      24254:data<=-16'd7410;
      24255:data<=-16'd7423;
      24256:data<=-16'd9347;
      24257:data<=-16'd9191;
      24258:data<=-16'd8234;
      24259:data<=-16'd8671;
      24260:data<=-16'd7887;
      24261:data<=-16'd7083;
      24262:data<=-16'd6949;
      24263:data<=-16'd5930;
      24264:data<=-16'd5880;
      24265:data<=-16'd6106;
      24266:data<=-16'd5518;
      24267:data<=-16'd6088;
      24268:data<=-16'd7022;
      24269:data<=-16'd7194;
      24270:data<=-16'd6733;
      24271:data<=-16'd5783;
      24272:data<=-16'd5353;
      24273:data<=-16'd5078;
      24274:data<=-16'd5030;
      24275:data<=-16'd5013;
      24276:data<=-16'd4112;
      24277:data<=-16'd4294;
      24278:data<=-16'd3987;
      24279:data<=-16'd2547;
      24280:data<=-16'd4631;
      24281:data<=-16'd3398;
      24282:data<=16'd5876;
      24283:data<=16'd10147;
      24284:data<=16'd8012;
      24285:data<=16'd8736;
      24286:data<=16'd8900;
      24287:data<=16'd7512;
      24288:data<=16'd8366;
      24289:data<=16'd7529;
      24290:data<=16'd4631;
      24291:data<=16'd3667;
      24292:data<=16'd3444;
      24293:data<=16'd2346;
      24294:data<=16'd1347;
      24295:data<=16'd1387;
      24296:data<=16'd1858;
      24297:data<=16'd1718;
      24298:data<=16'd1779;
      24299:data<=16'd2002;
      24300:data<=16'd1680;
      24301:data<=16'd1997;
      24302:data<=16'd2584;
      24303:data<=16'd2334;
      24304:data<=16'd2161;
      24305:data<=16'd1845;
      24306:data<=16'd754;
      24307:data<=16'd152;
      24308:data<=16'd438;
      24309:data<=16'd528;
      24310:data<=16'd262;
      24311:data<=16'd234;
      24312:data<=16'd276;
      24313:data<=16'd388;
      24314:data<=16'd876;
      24315:data<=16'd1095;
      24316:data<=16'd1080;
      24317:data<=16'd1095;
      24318:data<=16'd308;
      24319:data<=-16'd382;
      24320:data<=-16'd221;
      24321:data<=-16'd440;
      24322:data<=-16'd496;
      24323:data<=-16'd50;
      24324:data<=-16'd50;
      24325:data<=16'd306;
      24326:data<=16'd1099;
      24327:data<=16'd1269;
      24328:data<=16'd719;
      24329:data<=16'd513;
      24330:data<=16'd1363;
      24331:data<=-16'd1504;
      24332:data<=-16'd10091;
      24333:data<=-16'd14982;
      24334:data<=-16'd13332;
      24335:data<=-16'd12592;
      24336:data<=-16'd12681;
      24337:data<=-16'd11467;
      24338:data<=-16'd11104;
      24339:data<=-16'd10568;
      24340:data<=-16'd9476;
      24341:data<=-16'd9253;
      24342:data<=-16'd9256;
      24343:data<=-16'd9438;
      24344:data<=-16'd9498;
      24345:data<=-16'd9224;
      24346:data<=-16'd9238;
      24347:data<=-16'd8452;
      24348:data<=-16'd7363;
      24349:data<=-16'd7063;
      24350:data<=-16'd6335;
      24351:data<=-16'd6100;
      24352:data<=-16'd6488;
      24353:data<=-16'd5272;
      24354:data<=-16'd4326;
      24355:data<=-16'd4777;
      24356:data<=-16'd3328;
      24357:data<=-16'd420;
      24358:data<=16'd678;
      24359:data<=16'd584;
      24360:data<=16'd928;
      24361:data<=16'd1169;
      24362:data<=16'd1421;
      24363:data<=16'd2003;
      24364:data<=16'd1947;
      24365:data<=16'd1820;
      24366:data<=16'd2173;
      24367:data<=16'd2173;
      24368:data<=16'd3069;
      24369:data<=16'd4758;
      24370:data<=16'd4971;
      24371:data<=16'd4901;
      24372:data<=16'd5388;
      24373:data<=16'd5204;
      24374:data<=16'd4977;
      24375:data<=16'd4855;
      24376:data<=16'd4773;
      24377:data<=16'd4916;
      24378:data<=16'd4637;
      24379:data<=16'd4692;
      24380:data<=16'd4778;
      24381:data<=16'd6519;
      24382:data<=16'd13838;
      24383:data<=16'd20401;
      24384:data<=16'd19930;
      24385:data<=16'd18738;
      24386:data<=16'd18958;
      24387:data<=16'd17981;
      24388:data<=16'd17596;
      24389:data<=16'd16804;
      24390:data<=16'd15688;
      24391:data<=16'd16158;
      24392:data<=16'd15734;
      24393:data<=16'd15245;
      24394:data<=16'd16137;
      24395:data<=16'd15810;
      24396:data<=16'd15362;
      24397:data<=16'd15417;
      24398:data<=16'd14236;
      24399:data<=16'd13330;
      24400:data<=16'd12969;
      24401:data<=16'd12360;
      24402:data<=16'd12340;
      24403:data<=16'd12034;
      24404:data<=16'd10975;
      24405:data<=16'd10816;
      24406:data<=16'd11928;
      24407:data<=16'd12317;
      24408:data<=16'd11282;
      24409:data<=16'd10887;
      24410:data<=16'd10857;
      24411:data<=16'd9962;
      24412:data<=16'd9596;
      24413:data<=16'd9153;
      24414:data<=16'd8196;
      24415:data<=16'd8164;
      24416:data<=16'd7702;
      24417:data<=16'd6852;
      24418:data<=16'd7588;
      24419:data<=16'd8819;
      24420:data<=16'd8947;
      24421:data<=16'd8064;
      24422:data<=16'd7515;
      24423:data<=16'd6851;
      24424:data<=16'd4852;
      24425:data<=16'd4325;
      24426:data<=16'd4958;
      24427:data<=16'd4088;
      24428:data<=16'd3803;
      24429:data<=16'd3298;
      24430:data<=16'd3362;
      24431:data<=16'd5824;
      24432:data<=16'd1591;
      24433:data<=-16'd7950;
      24434:data<=-16'd9529;
      24435:data<=-16'd7642;
      24436:data<=-16'd8900;
      24437:data<=-16'd8508;
      24438:data<=-16'd7680;
      24439:data<=-16'd7694;
      24440:data<=-16'd6555;
      24441:data<=-16'd6531;
      24442:data<=-16'd7169;
      24443:data<=-16'd6416;
      24444:data<=-16'd4915;
      24445:data<=-16'd3654;
      24446:data<=-16'd3918;
      24447:data<=-16'd4463;
      24448:data<=-16'd3924;
      24449:data<=-16'd3485;
      24450:data<=-16'd3113;
      24451:data<=-16'd3248;
      24452:data<=-16'd3673;
      24453:data<=-16'd3054;
      24454:data<=-16'd2919;
      24455:data<=-16'd2924;
      24456:data<=-16'd1588;
      24457:data<=-16'd597;
      24458:data<=-16'd187;
      24459:data<=16'd6;
      24460:data<=-16'd129;
      24461:data<=16'd70;
      24462:data<=-16'd167;
      24463:data<=-16'd102;
      24464:data<=16'd887;
      24465:data<=16'd766;
      24466:data<=16'd140;
      24467:data<=16'd58;
      24468:data<=16'd466;
      24469:data<=16'd1779;
      24470:data<=16'd2362;
      24471:data<=16'd2224;
      24472:data<=16'd2215;
      24473:data<=16'd1582;
      24474:data<=16'd1720;
      24475:data<=16'd1800;
      24476:data<=16'd1140;
      24477:data<=16'd1809;
      24478:data<=16'd1554;
      24479:data<=16'd1221;
      24480:data<=16'd2049;
      24481:data<=16'd825;
      24482:data<=16'd5004;
      24483:data<=16'd15365;
      24484:data<=16'd17506;
      24485:data<=16'd14383;
      24486:data<=16'd14662;
      24487:data<=16'd14102;
      24488:data<=16'd13411;
      24489:data<=16'd13365;
      24490:data<=16'd12331;
      24491:data<=16'd13156;
      24492:data<=16'd13520;
      24493:data<=16'd12897;
      24494:data<=16'd13961;
      24495:data<=16'd13637;
      24496:data<=16'd12836;
      24497:data<=16'd12880;
      24498:data<=16'd11415;
      24499:data<=16'd10724;
      24500:data<=16'd10680;
      24501:data<=16'd9691;
      24502:data<=16'd9491;
      24503:data<=16'd8981;
      24504:data<=16'd8131;
      24505:data<=16'd8011;
      24506:data<=16'd8044;
      24507:data<=16'd8695;
      24508:data<=16'd8472;
      24509:data<=16'd7383;
      24510:data<=16'd7028;
      24511:data<=16'd6431;
      24512:data<=16'd6639;
      24513:data<=16'd6492;
      24514:data<=16'd4672;
      24515:data<=16'd4722;
      24516:data<=16'd4657;
      24517:data<=16'd3377;
      24518:data<=16'd4481;
      24519:data<=16'd5297;
      24520:data<=16'd4948;
      24521:data<=16'd4839;
      24522:data<=16'd3812;
      24523:data<=16'd3876;
      24524:data<=16'd3956;
      24525:data<=16'd2983;
      24526:data<=16'd3203;
      24527:data<=16'd2528;
      24528:data<=16'd2023;
      24529:data<=16'd2041;
      24530:data<=16'd916;
      24531:data<=16'd3096;
      24532:data<=16'd1571;
      24533:data<=-16'd8522;
      24534:data<=-16'd11920;
      24535:data<=-16'd8901;
      24536:data<=-16'd9917;
      24537:data<=-16'd10135;
      24538:data<=-16'd9571;
      24539:data<=-16'd10357;
      24540:data<=-16'd9135;
      24541:data<=-16'd8974;
      24542:data<=-16'd9873;
      24543:data<=-16'd8680;
      24544:data<=-16'd7083;
      24545:data<=-16'd5968;
      24546:data<=-16'd6214;
      24547:data<=-16'd6912;
      24548:data<=-16'd6338;
      24549:data<=-16'd6216;
      24550:data<=-16'd5976;
      24551:data<=-16'd5647;
      24552:data<=-16'd6455;
      24553:data<=-16'd6226;
      24554:data<=-16'd5532;
      24555:data<=-16'd5529;
      24556:data<=-16'd5339;
      24557:data<=-16'd5921;
      24558:data<=-16'd6815;
      24559:data<=-16'd7356;
      24560:data<=-16'd7382;
      24561:data<=-16'd6525;
      24562:data<=-16'd6755;
      24563:data<=-16'd6957;
      24564:data<=-16'd6011;
      24565:data<=-16'd6347;
      24566:data<=-16'd6202;
      24567:data<=-16'd5400;
      24568:data<=-16'd6534;
      24569:data<=-16'd7676;
      24570:data<=-16'd8164;
      24571:data<=-16'd8214;
      24572:data<=-16'd7667;
      24573:data<=-16'd7699;
      24574:data<=-16'd6996;
      24575:data<=-16'd6766;
      24576:data<=-16'd7627;
      24577:data<=-16'd6833;
      24578:data<=-16'd7087;
      24579:data<=-16'd7048;
      24580:data<=-16'd5187;
      24581:data<=-16'd7524;
      24582:data<=-16'd6167;
      24583:data<=16'd3748;
      24584:data<=16'd6899;
      24585:data<=16'd3876;
      24586:data<=16'd4872;
      24587:data<=16'd5157;
      24588:data<=16'd4299;
      24589:data<=16'd4878;
      24590:data<=16'd3952;
      24591:data<=16'd3463;
      24592:data<=16'd3896;
      24593:data<=16'd2773;
      24594:data<=16'd1451;
      24595:data<=16'd617;
      24596:data<=16'd376;
      24597:data<=16'd663;
      24598:data<=16'd514;
      24599:data<=16'd394;
      24600:data<=-16'd130;
      24601:data<=-16'd611;
      24602:data<=16'd441;
      24603:data<=16'd849;
      24604:data<=-16'd70;
      24605:data<=-16'd109;
      24606:data<=-16'd532;
      24607:data<=-16'd2500;
      24608:data<=-16'd3427;
      24609:data<=-16'd2767;
      24610:data<=-16'd2874;
      24611:data<=-16'd3189;
      24612:data<=-16'd2657;
      24613:data<=-16'd3058;
      24614:data<=-16'd3491;
      24615:data<=-16'd2757;
      24616:data<=-16'd2996;
      24617:data<=-16'd3297;
      24618:data<=-16'd2949;
      24619:data<=-16'd4073;
      24620:data<=-16'd4962;
      24621:data<=-16'd4581;
      24622:data<=-16'd4629;
      24623:data<=-16'd4575;
      24624:data<=-16'd4026;
      24625:data<=-16'd2881;
      24626:data<=-16'd1886;
      24627:data<=-16'd1986;
      24628:data<=-16'd1269;
      24629:data<=-16'd1186;
      24630:data<=-16'd2226;
      24631:data<=-16'd1256;
      24632:data<=-16'd5013;
      24633:data<=-16'd15013;
      24634:data<=-16'd18175;
      24635:data<=-16'd15386;
      24636:data<=-16'd15600;
      24637:data<=-16'd15617;
      24638:data<=-16'd14510;
      24639:data<=-16'd14509;
      24640:data<=-16'd13678;
      24641:data<=-16'd12834;
      24642:data<=-16'd12675;
      24643:data<=-16'd12624;
      24644:data<=-16'd13212;
      24645:data<=-16'd13220;
      24646:data<=-16'd12903;
      24647:data<=-16'd12768;
      24648:data<=-16'd11720;
      24649:data<=-16'd11189;
      24650:data<=-16'd11112;
      24651:data<=-16'd10107;
      24652:data<=-16'd9744;
      24653:data<=-16'd9856;
      24654:data<=-16'd9075;
      24655:data<=-16'd8410;
      24656:data<=-16'd8995;
      24657:data<=-16'd10237;
      24658:data<=-16'd10228;
      24659:data<=-16'd9368;
      24660:data<=-16'd9291;
      24661:data<=-16'd8875;
      24662:data<=-16'd8028;
      24663:data<=-16'd7623;
      24664:data<=-16'd6902;
      24665:data<=-16'd6246;
      24666:data<=-16'd5934;
      24667:data<=-16'd5724;
      24668:data<=-16'd6225;
      24669:data<=-16'd6916;
      24670:data<=-16'd7127;
      24671:data<=-16'd6686;
      24672:data<=-16'd5999;
      24673:data<=-16'd5824;
      24674:data<=-16'd5362;
      24675:data<=-16'd5062;
      24676:data<=-16'd5236;
      24677:data<=-16'd4608;
      24678:data<=-16'd4748;
      24679:data<=-16'd4400;
      24680:data<=-16'd2685;
      24681:data<=-16'd4584;
      24682:data<=-16'd4381;
      24683:data<=16'd4325;
      24684:data<=16'd10009;
      24685:data<=16'd8505;
      24686:data<=16'd8149;
      24687:data<=16'd8454;
      24688:data<=16'd7835;
      24689:data<=16'd8264;
      24690:data<=16'd8331;
      24691:data<=16'd7550;
      24692:data<=16'd6611;
      24693:data<=16'd5726;
      24694:data<=16'd4869;
      24695:data<=16'd3797;
      24696:data<=16'd3808;
      24697:data<=16'd3990;
      24698:data<=16'd3095;
      24699:data<=16'd3240;
      24700:data<=16'd3492;
      24701:data<=16'd2919;
      24702:data<=16'd3427;
      24703:data<=16'd3609;
      24704:data<=16'd3137;
      24705:data<=16'd3307;
      24706:data<=16'd2725;
      24707:data<=16'd1838;
      24708:data<=16'd1547;
      24709:data<=16'd1316;
      24710:data<=16'd1459;
      24711:data<=16'd1177;
      24712:data<=16'd584;
      24713:data<=16'd760;
      24714:data<=16'd1080;
      24715:data<=16'd1377;
      24716:data<=16'd1039;
      24717:data<=16'd641;
      24718:data<=16'd1700;
      24719:data<=16'd1354;
      24720:data<=-16'd608;
      24721:data<=-16'd701;
      24722:data<=-16'd352;
      24723:data<=-16'd409;
      24724:data<=-16'd6;
      24725:data<=-16'd202;
      24726:data<=16'd86;
      24727:data<=16'd682;
      24728:data<=16'd379;
      24729:data<=16'd409;
      24730:data<=16'd303;
      24731:data<=16'd415;
      24732:data<=-16'd1090;
      24733:data<=-16'd8733;
      24734:data<=-16'd15524;
      24735:data<=-16'd14574;
      24736:data<=-16'd12595;
      24737:data<=-16'd12398;
      24738:data<=-16'd11629;
      24739:data<=-16'd11471;
      24740:data<=-16'd11100;
      24741:data<=-16'd10299;
      24742:data<=-16'd9962;
      24743:data<=-16'd9362;
      24744:data<=-16'd9888;
      24745:data<=-16'd10942;
      24746:data<=-16'd10557;
      24747:data<=-16'd10013;
      24748:data<=-16'd9175;
      24749:data<=-16'd8047;
      24750:data<=-16'd7741;
      24751:data<=-16'd7156;
      24752:data<=-16'd6684;
      24753:data<=-16'd6865;
      24754:data<=-16'd6276;
      24755:data<=-16'd5236;
      24756:data<=-16'd4817;
      24757:data<=-16'd5057;
      24758:data<=-16'd4396;
      24759:data<=-16'd2309;
      24760:data<=-16'd1400;
      24761:data<=-16'd1278;
      24762:data<=-16'd419;
      24763:data<=-16'd314;
      24764:data<=-16'd329;
      24765:data<=16'd203;
      24766:data<=16'd629;
      24767:data<=16'd1155;
      24768:data<=16'd795;
      24769:data<=16'd1272;
      24770:data<=16'd3438;
      24771:data<=16'd3639;
      24772:data<=16'd3474;
      24773:data<=16'd4332;
      24774:data<=16'd3645;
      24775:data<=16'd3550;
      24776:data<=16'd4034;
      24777:data<=16'd3410;
      24778:data<=16'd3641;
      24779:data<=16'd3798;
      24780:data<=16'd4082;
      24781:data<=16'd4676;
      24782:data<=16'd4813;
      24783:data<=16'd10546;
      24784:data<=16'd18983;
      24785:data<=16'd19873;
      24786:data<=16'd17841;
      24787:data<=16'd17884;
      24788:data<=16'd17478;
      24789:data<=16'd17569;
      24790:data<=16'd16810;
      24791:data<=16'd15356;
      24792:data<=16'd15602;
      24793:data<=16'd14906;
      24794:data<=16'd14766;
      24795:data<=16'd16521;
      24796:data<=16'd16104;
      24797:data<=16'd15065;
      24798:data<=16'd14959;
      24799:data<=16'd14119;
      24800:data<=16'd13761;
      24801:data<=16'd13309;
      24802:data<=16'd12377;
      24803:data<=16'd12331;
      24804:data<=16'd11862;
      24805:data<=16'd10988;
      24806:data<=16'd11239;
      24807:data<=16'd12354;
      24808:data<=16'd12847;
      24809:data<=16'd11966;
      24810:data<=16'd11471;
      24811:data<=16'd11163;
      24812:data<=16'd9996;
      24813:data<=16'd9973;
      24814:data<=16'd10076;
      24815:data<=16'd9083;
      24816:data<=16'd8484;
      24817:data<=16'd7321;
      24818:data<=16'd6768;
      24819:data<=16'd8153;
      24820:data<=16'd8992;
      24821:data<=16'd9142;
      24822:data<=16'd8536;
      24823:data<=16'd7729;
      24824:data<=16'd8187;
      24825:data<=16'd6981;
      24826:data<=16'd4983;
      24827:data<=16'd4693;
      24828:data<=16'd3938;
      24829:data<=16'd3947;
      24830:data<=16'd3803;
      24831:data<=16'd2978;
      24832:data<=16'd5422;
      24833:data<=16'd3039;
      24834:data<=-16'd6661;
      24835:data<=-16'd9511;
      24836:data<=-16'd7233;
      24837:data<=-16'd8170;
      24838:data<=-16'd7956;
      24839:data<=-16'd7207;
      24840:data<=-16'd7794;
      24841:data<=-16'd7083;
      24842:data<=-16'd6863;
      24843:data<=-16'd6954;
      24844:data<=-16'd5934;
      24845:data<=-16'd5216;
      24846:data<=-16'd4704;
      24847:data<=-16'd4475;
      24848:data<=-16'd4041;
      24849:data<=-16'd3294;
      24850:data<=-16'd3574;
      24851:data<=-16'd3262;
      24852:data<=-16'd2620;
      24853:data<=-16'd3310;
      24854:data<=-16'd3239;
      24855:data<=-16'd2728;
      24856:data<=-16'd2763;
      24857:data<=-16'd1718;
      24858:data<=-16'd443;
      24859:data<=-16'd123;
      24860:data<=-16'd306;
      24861:data<=-16'd343;
      24862:data<=16'd165;
      24863:data<=16'd262;
      24864:data<=-16'd53;
      24865:data<=-16'd290;
      24866:data<=-16'd359;
      24867:data<=16'd340;
      24868:data<=16'd440;
      24869:data<=16'd393;
      24870:data<=16'd1694;
      24871:data<=16'd1829;
      24872:data<=16'd1638;
      24873:data<=16'd2538;
      24874:data<=16'd1944;
      24875:data<=16'd1404;
      24876:data<=16'd1641;
      24877:data<=16'd1377;
      24878:data<=16'd1717;
      24879:data<=16'd698;
      24880:data<=16'd83;
      24881:data<=16'd1710;
      24882:data<=16'd1336;
      24883:data<=16'd5225;
      24884:data<=16'd14954;
      24885:data<=16'd16950;
      24886:data<=16'd14066;
      24887:data<=16'd14687;
      24888:data<=16'd13606;
      24889:data<=16'd12178;
      24890:data<=16'd12722;
      24891:data<=16'd11708;
      24892:data<=16'd11590;
      24893:data<=16'd12605;
      24894:data<=16'd12781;
      24895:data<=16'd13764;
      24896:data<=16'd14104;
      24897:data<=16'd13174;
      24898:data<=16'd12396;
      24899:data<=16'd11389;
      24900:data<=16'd10912;
      24901:data<=16'd10643;
      24902:data<=16'd9879;
      24903:data<=16'd9542;
      24904:data<=16'd8933;
      24905:data<=16'd8075;
      24906:data<=16'd8125;
      24907:data<=16'd8765;
      24908:data<=16'd8983;
      24909:data<=16'd8428;
      24910:data<=16'd8267;
      24911:data<=16'd7803;
      24912:data<=16'd6401;
      24913:data<=16'd6469;
      24914:data<=16'd6419;
      24915:data<=16'd5136;
      24916:data<=16'd5357;
      24917:data<=16'd4692;
      24918:data<=16'd2975;
      24919:data<=16'd3888;
      24920:data<=16'd5218;
      24921:data<=16'd5427;
      24922:data<=16'd5015;
      24923:data<=16'd4009;
      24924:data<=16'd4074;
      24925:data<=16'd3882;
      24926:data<=16'd3312;
      24927:data<=16'd3439;
      24928:data<=16'd2364;
      24929:data<=16'd2372;
      24930:data<=16'd2510;
      24931:data<=16'd672;
      24932:data<=16'd2394;
      24933:data<=16'd1441;
      24934:data<=-16'd7561;
      24935:data<=-16'd11210;
      24936:data<=-16'd9091;
      24937:data<=-16'd9867;
      24938:data<=-16'd9767;
      24939:data<=-16'd9374;
      24940:data<=-16'd10155;
      24941:data<=-16'd9033;
      24942:data<=-16'd8943;
      24943:data<=-16'd9486;
      24944:data<=-16'd8156;
      24945:data<=-16'd7213;
      24946:data<=-16'd6563;
      24947:data<=-16'd6150;
      24948:data<=-16'd6150;
      24949:data<=-16'd5771;
      24950:data<=-16'd6196;
      24951:data<=-16'd6175;
      24952:data<=-16'd5471;
      24953:data<=-16'd6026;
      24954:data<=-16'd6138;
      24955:data<=-16'd5803;
      24956:data<=-16'd6029;
      24957:data<=-16'd5550;
      24958:data<=-16'd5210;
      24959:data<=-16'd5858;
      24960:data<=-16'd7144;
      24961:data<=-16'd7834;
      24962:data<=-16'd6842;
      24963:data<=-16'd6575;
      24964:data<=-16'd7066;
      24965:data<=-16'd6672;
      24966:data<=-16'd6784;
      24967:data<=-16'd6367;
      24968:data<=-16'd5439;
      24969:data<=-16'd6190;
      24970:data<=-16'd7268;
      24971:data<=-16'd8102;
      24972:data<=-16'd8211;
      24973:data<=-16'd7418;
      24974:data<=-16'd7696;
      24975:data<=-16'd7427;
      24976:data<=-16'd6670;
      24977:data<=-16'd6839;
      24978:data<=-16'd6003;
      24979:data<=-16'd6209;
      24980:data<=-16'd6357;
      24981:data<=-16'd4579;
      24982:data<=-16'd6499;
      24983:data<=-16'd5846;
      24984:data<=16'd3092;
      24985:data<=16'd7094;
      24986:data<=16'd4819;
      24987:data<=16'd5275;
      24988:data<=16'd5310;
      24989:data<=16'd4300;
      24990:data<=16'd4821;
      24991:data<=16'd4698;
      24992:data<=16'd4356;
      24993:data<=16'd4006;
      24994:data<=16'd3036;
      24995:data<=16'd2350;
      24996:data<=16'd1610;
      24997:data<=16'd1222;
      24998:data<=16'd1014;
      24999:data<=16'd516;
      25000:data<=16'd878;
      25001:data<=16'd1077;
      25002:data<=16'd596;
      25003:data<=16'd690;
      25004:data<=16'd755;
      25005:data<=16'd634;
      25006:data<=16'd446;
      25007:data<=-16'd506;
      25008:data<=-16'd1876;
      25009:data<=-16'd2416;
      25010:data<=-16'd1603;
      25011:data<=-16'd1541;
      25012:data<=-16'd2679;
      25013:data<=-16'd2488;
      25014:data<=-16'd2155;
      25015:data<=-16'd2540;
      25016:data<=-16'd1865;
      25017:data<=-16'd1457;
      25018:data<=-16'd1794;
      25019:data<=-16'd2278;
      25020:data<=-16'd3536;
      25021:data<=-16'd4050;
      25022:data<=-16'd3776;
      25023:data<=-16'd3789;
      25024:data<=-16'd3577;
      25025:data<=-16'd3571;
      25026:data<=-16'd2569;
      25027:data<=-16'd879;
      25028:data<=-16'd1025;
      25029:data<=-16'd1071;
      25030:data<=-16'd1083;
      25031:data<=-16'd1751;
      25032:data<=-16'd789;
      25033:data<=-16'd3977;
      25034:data<=-16'd13053;
      25035:data<=-16'd17243;
      25036:data<=-16'd15649;
      25037:data<=-16'd14697;
      25038:data<=-16'd13957;
      25039:data<=-16'd13597;
      25040:data<=-16'd13826;
      25041:data<=-16'd12851;
      25042:data<=-16'd11975;
      25043:data<=-16'd11652;
      25044:data<=-16'd11229;
      25045:data<=-16'd11806;
      25046:data<=-16'd12698;
      25047:data<=-16'd12402;
      25048:data<=-16'd11512;
      25049:data<=-16'd10757;
      25050:data<=-16'd9903;
      25051:data<=-16'd9162;
      25052:data<=-16'd8907;
      25053:data<=-16'd8498;
      25054:data<=-16'd8103;
      25055:data<=-16'd8185;
      25056:data<=-16'd7685;
      25057:data<=-16'd7474;
      25058:data<=-16'd8695;
      25059:data<=-16'd9332;
      25060:data<=-16'd8953;
      25061:data<=-16'd8345;
      25062:data<=-16'd7151;
      25063:data<=-16'd6643;
      25064:data<=-16'd6802;
      25065:data<=-16'd6115;
      25066:data<=-16'd5635;
      25067:data<=-16'd5535;
      25068:data<=-16'd4775;
      25069:data<=-16'd4275;
      25070:data<=-16'd4836;
      25071:data<=-16'd5940;
      25072:data<=-16'd6112;
      25073:data<=-16'd5086;
      25074:data<=-16'd4458;
      25075:data<=-16'd4179;
      25076:data<=-16'd4115;
      25077:data<=-16'd4215;
      25078:data<=-16'd3234;
      25079:data<=-16'd3008;
      25080:data<=-16'd3315;
      25081:data<=-16'd1780;
      25082:data<=-16'd2414;
      25083:data<=-16'd3016;
      25084:data<=16'd3659;
      25085:data<=16'd9996;
      25086:data<=16'd9591;
      25087:data<=16'd9103;
      25088:data<=16'd9588;
      25089:data<=16'd8990;
      25090:data<=16'd9222;
      25091:data<=16'd9480;
      25092:data<=16'd9138;
      25093:data<=16'd8222;
      25094:data<=16'd6135;
      25095:data<=16'd4673;
      25096:data<=16'd4199;
      25097:data<=16'd3885;
      25098:data<=16'd3838;
      25099:data<=16'd3345;
      25100:data<=16'd3239;
      25101:data<=16'd3747;
      25102:data<=16'd3327;
      25103:data<=16'd2992;
      25104:data<=16'd3418;
      25105:data<=16'd3662;
      25106:data<=16'd3430;
      25107:data<=16'd2296;
      25108:data<=16'd1113;
      25109:data<=16'd890;
      25110:data<=16'd1186;
      25111:data<=16'd1427;
      25112:data<=16'd905;
      25113:data<=16'd620;
      25114:data<=16'd1178;
      25115:data<=16'd1199;
      25116:data<=16'd1592;
      25117:data<=16'd1929;
      25118:data<=16'd869;
      25119:data<=16'd684;
      25120:data<=16'd540;
      25121:data<=-16'd713;
      25122:data<=-16'd710;
      25123:data<=-16'd805;
      25124:data<=-16'd1312;
      25125:data<=-16'd514;
      25126:data<=-16'd196;
      25127:data<=-16'd183;
      25128:data<=-16'd124;
      25129:data<=-16'd487;
      25130:data<=16'd79;
      25131:data<=-16'd285;
      25132:data<=-16'd913;
      25133:data<=-16'd1192;
      25134:data<=-16'd7386;
      25135:data<=-16'd14815;
      25136:data<=-16'd14689;
      25137:data<=-16'd13298;
      25138:data<=-16'd13759;
      25139:data<=-16'd12736;
      25140:data<=-16'd12319;
      25141:data<=-16'd11909;
      25142:data<=-16'd10887;
      25143:data<=-16'd10807;
      25144:data<=-16'd9693;
      25145:data<=-16'd9115;
      25146:data<=-16'd10681;
      25147:data<=-16'd11101;
      25148:data<=-16'd10443;
      25149:data<=-16'd9706;
      25150:data<=-16'd8557;
      25151:data<=-16'd8011;
      25152:data<=-16'd7494;
      25153:data<=-16'd6798;
      25154:data<=-16'd6519;
      25155:data<=-16'd6037;
      25156:data<=-16'd5711;
      25157:data<=-16'd5321;
      25158:data<=-16'd4651;
      25159:data<=-16'd4496;
      25160:data<=-16'd3767;
      25161:data<=-16'd2322;
      25162:data<=-16'd1381;
      25163:data<=-16'd745;
      25164:data<=-16'd532;
      25165:data<=-16'd558;
      25166:data<=-16'd335;
      25167:data<=-16'd15;
      25168:data<=16'd517;
      25169:data<=16'd884;
      25170:data<=16'd1645;
      25171:data<=16'd2907;
      25172:data<=16'd3083;
      25173:data<=16'd3159;
      25174:data<=16'd3548;
      25175:data<=16'd3377;
      25176:data<=16'd3864;
      25177:data<=16'd3965;
      25178:data<=16'd3618;
      25179:data<=16'd4076;
      25180:data<=16'd3394;
      25181:data<=16'd3792;
      25182:data<=16'd5024;
      25183:data<=16'd3777;
      25184:data<=16'd8557;
      25185:data<=16'd18639;
      25186:data<=16'd20102;
      25187:data<=16'd17613;
      25188:data<=16'd18689;
      25189:data<=16'd17755;
      25190:data<=16'd16393;
      25191:data<=16'd16868;
      25192:data<=16'd16093;
      25193:data<=16'd15379;
      25194:data<=16'd14816;
      25195:data<=16'd14574;
      25196:data<=16'd15941;
      25197:data<=16'd16126;
      25198:data<=16'd15353;
      25199:data<=16'd15074;
      25200:data<=16'd13961;
      25201:data<=16'd13400;
      25202:data<=16'd13383;
      25203:data<=16'd12214;
      25204:data<=16'd11309;
      25205:data<=16'd11135;
      25206:data<=16'd10839;
      25207:data<=16'd10575;
      25208:data<=16'd10975;
      25209:data<=16'd12040;
      25210:data<=16'd12023;
      25211:data<=16'd11056;
      25212:data<=16'd10666;
      25213:data<=16'd10207;
      25214:data<=16'd9729;
      25215:data<=16'd9433;
      25216:data<=16'd8810;
      25217:data<=16'd8426;
      25218:data<=16'd7755;
      25219:data<=16'd6928;
      25220:data<=16'd7511;
      25221:data<=16'd8840;
      25222:data<=16'd9388;
      25223:data<=16'd8610;
      25224:data<=16'd7630;
      25225:data<=16'd7413;
      25226:data<=16'd6877;
      25227:data<=16'd6090;
      25228:data<=16'd4645;
      25229:data<=16'd3134;
      25230:data<=16'd4161;
      25231:data<=16'd4000;
      25232:data<=16'd2728;
      25233:data<=16'd5356;
      25234:data<=16'd2889;
      25235:data<=-16'd6801;
      25236:data<=-16'd9456;
      25237:data<=-16'd7247;
      25238:data<=-16'd8381;
      25239:data<=-16'd8352;
      25240:data<=-16'd7533;
      25241:data<=-16'd8178;
      25242:data<=-16'd7915;
      25243:data<=-16'd7691;
      25244:data<=-16'd7424;
      25245:data<=-16'd6193;
      25246:data<=-16'd5048;
      25247:data<=-16'd4197;
      25248:data<=-16'd4114;
      25249:data<=-16'd3906;
      25250:data<=-16'd3354;
      25251:data<=-16'd3997;
      25252:data<=-16'd4197;
      25253:data<=-16'd3657;
      25254:data<=-16'd3761;
      25255:data<=-16'd3313;
      25256:data<=-16'd2874;
      25257:data<=-16'd2878;
      25258:data<=-16'd1882;
      25259:data<=-16'd526;
      25260:data<=16'd120;
      25261:data<=-16'd130;
      25262:data<=-16'd414;
      25263:data<=-16'd323;
      25264:data<=-16'd817;
      25265:data<=-16'd728;
      25266:data<=-16'd212;
      25267:data<=-16'd637;
      25268:data<=-16'd334;
      25269:data<=16'd38;
      25270:data<=-16'd24;
      25271:data<=16'd1090;
      25272:data<=16'd1524;
      25273:data<=16'd1474;
      25274:data<=16'd2018;
      25275:data<=16'd1685;
      25276:data<=16'd1525;
      25277:data<=16'd1115;
      25278:data<=16'd795;
      25279:data<=16'd1964;
      25280:data<=16'd970;
      25281:data<=-16'd61;
      25282:data<=16'd814;
      25283:data<=-16'd252;
      25284:data<=16'd4311;
      25285:data<=16'd14609;
      25286:data<=16'd16395;
      25287:data<=16'd13541;
      25288:data<=16'd14088;
      25289:data<=16'd13479;
      25290:data<=16'd12542;
      25291:data<=16'd12511;
      25292:data<=16'd11523;
      25293:data<=16'd11150;
      25294:data<=16'd11038;
      25295:data<=16'd11746;
      25296:data<=16'd13321;
      25297:data<=16'd13204;
      25298:data<=16'd12862;
      25299:data<=16'd12417;
      25300:data<=16'd10831;
      25301:data<=16'd10120;
      25302:data<=16'd9705;
      25303:data<=16'd9200;
      25304:data<=16'd8930;
      25305:data<=16'd7834;
      25306:data<=16'd6969;
      25307:data<=16'd6425;
      25308:data<=16'd6586;
      25309:data<=16'd8032;
      25310:data<=16'd7818;
      25311:data<=16'd6953;
      25312:data<=16'd6993;
      25313:data<=16'd5852;
      25314:data<=16'd5316;
      25315:data<=16'd5095;
      25316:data<=16'd3667;
      25317:data<=16'd3853;
      25318:data<=16'd3833;
      25319:data<=16'd2356;
      25320:data<=16'd2880;
      25321:data<=16'd4399;
      25322:data<=16'd5080;
      25323:data<=16'd4822;
      25324:data<=16'd3976;
      25325:data<=16'd3659;
      25326:data<=16'd2908;
      25327:data<=16'd2566;
      25328:data<=16'd2711;
      25329:data<=16'd1536;
      25330:data<=16'd2002;
      25331:data<=16'd2332;
      25332:data<=16'd851;
      25333:data<=16'd2954;
      25334:data<=16'd1424;
      25335:data<=-16'd7947;
      25336:data<=-16'd11612;
      25337:data<=-16'd9903;
      25338:data<=-16'd10880;
      25339:data<=-16'd10695;
      25340:data<=-16'd9867;
      25341:data<=-16'd10357;
      25342:data<=-16'd9703;
      25343:data<=-16'd9599;
      25344:data<=-16'd9984;
      25345:data<=-16'd9153;
      25346:data<=-16'd7924;
      25347:data<=-16'd6796;
      25348:data<=-16'd6893;
      25349:data<=-16'd7162;
      25350:data<=-16'd6501;
      25351:data<=-16'd6722;
      25352:data<=-16'd6637;
      25353:data<=-16'd5971;
      25354:data<=-16'd6322;
      25355:data<=-16'd5911;
      25356:data<=-16'd5213;
      25357:data<=-16'd5509;
      25358:data<=-16'd5327;
      25359:data<=-16'd5059;
      25360:data<=-16'd5100;
      25361:data<=-16'd5641;
      25362:data<=-16'd7066;
      25363:data<=-16'd7345;
      25364:data<=-16'd6681;
      25365:data<=-16'd6567;
      25366:data<=-16'd6179;
      25367:data<=-16'd6065;
      25368:data<=-16'd6282;
      25369:data<=-16'd5695;
      25370:data<=-16'd5550;
      25371:data<=-16'd6704;
      25372:data<=-16'd7773;
      25373:data<=-16'd7670;
      25374:data<=-16'd7383;
      25375:data<=-16'd7520;
      25376:data<=-16'd7022;
      25377:data<=-16'd6880;
      25378:data<=-16'd6928;
      25379:data<=-16'd5780;
      25380:data<=-16'd5955;
      25381:data<=-16'd6109;
      25382:data<=-16'd4848;
      25383:data<=-16'd6822;
      25384:data<=-16'd6223;
      25385:data<=16'd2246;
      25386:data<=16'd6792;
      25387:data<=16'd4977;
      25388:data<=16'd5192;
      25389:data<=16'd5350;
      25390:data<=16'd4420;
      25391:data<=16'd4945;
      25392:data<=16'd4637;
      25393:data<=16'd4337;
      25394:data<=16'd4913;
      25395:data<=16'd3871;
      25396:data<=16'd2275;
      25397:data<=16'd1495;
      25398:data<=16'd1166;
      25399:data<=16'd1300;
      25400:data<=16'd1213;
      25401:data<=16'd999;
      25402:data<=16'd851;
      25403:data<=16'd514;
      25404:data<=16'd490;
      25405:data<=16'd312;
      25406:data<=16'd6;
      25407:data<=16'd36;
      25408:data<=-16'd963;
      25409:data<=-16'd2611;
      25410:data<=-16'd2960;
      25411:data<=-16'd2344;
      25412:data<=-16'd2015;
      25413:data<=-16'd2246;
      25414:data<=-16'd2405;
      25415:data<=-16'd2284;
      25416:data<=-16'd2285;
      25417:data<=-16'd2076;
      25418:data<=-16'd1744;
      25419:data<=-16'd1783;
      25420:data<=-16'd2355;
      25421:data<=-16'd3615;
      25422:data<=-16'd4396;
      25423:data<=-16'd4003;
      25424:data<=-16'd3524;
      25425:data<=-16'd3409;
      25426:data<=-16'd3642;
      25427:data<=-16'd3400;
      25428:data<=-16'd2423;
      25429:data<=-16'd2005;
      25430:data<=-16'd1331;
      25431:data<=-16'd775;
      25432:data<=-16'd1371;
      25433:data<=-16'd961;
      25434:data<=-16'd3475;
      25435:data<=-16'd11867;
      25436:data<=-16'd16822;
      25437:data<=-16'd15756;
      25438:data<=-16'd15103;
      25439:data<=-16'd14577;
      25440:data<=-16'd13794;
      25441:data<=-16'd13564;
      25442:data<=-16'd12298;
      25443:data<=-16'd11932;
      25444:data<=-16'd12466;
      25445:data<=-16'd11747;
      25446:data<=-16'd11832;
      25447:data<=-16'd12604;
      25448:data<=-16'd12420;
      25449:data<=-16'd12328;
      25450:data<=-16'd11872;
      25451:data<=-16'd10689;
      25452:data<=-16'd9967;
      25453:data<=-16'd9670;
      25454:data<=-16'd9124;
      25455:data<=-16'd8200;
      25456:data<=-16'd7426;
      25457:data<=-16'd6893;
      25458:data<=-16'd7063;
      25459:data<=-16'd8411;
      25460:data<=-16'd8715;
      25461:data<=-16'd7865;
      25462:data<=-16'd8059;
      25463:data<=-16'd7793;
      25464:data<=-16'd6909;
      25465:data<=-16'd6751;
      25466:data<=-16'd6020;
      25467:data<=-16'd5603;
      25468:data<=-16'd5805;
      25469:data<=-16'd4852;
      25470:data<=-16'd4264;
      25471:data<=-16'd4757;
      25472:data<=-16'd5379;
      25473:data<=-16'd5839;
      25474:data<=-16'd5348;
      25475:data<=-16'd5145;
      25476:data<=-16'd5306;
      25477:data<=-16'd4451;
      25478:data<=-16'd4044;
      25479:data<=-16'd3532;
      25480:data<=-16'd2958;
      25481:data<=-16'd3553;
      25482:data<=-16'd2604;
      25483:data<=-16'd2720;
      25484:data<=-16'd4346;
      25485:data<=16'd1284;
      25486:data<=16'd9218;
      25487:data<=16'd9567;
      25488:data<=16'd8266;
      25489:data<=16'd8837;
      25490:data<=16'd8636;
      25491:data<=16'd8686;
      25492:data<=16'd8275;
      25493:data<=16'd8003;
      25494:data<=16'd8807;
      25495:data<=16'd7762;
      25496:data<=16'd5388;
      25497:data<=16'd3679;
      25498:data<=16'd3021;
      25499:data<=16'd3704;
      25500:data<=16'd3703;
      25501:data<=16'd3045;
      25502:data<=16'd3260;
      25503:data<=16'd3169;
      25504:data<=16'd3074;
      25505:data<=16'd3078;
      25506:data<=16'd2628;
      25507:data<=16'd2866;
      25508:data<=16'd2331;
      25509:data<=16'd594;
      25510:data<=16'd143;
      25511:data<=16'd426;
      25512:data<=16'd623;
      25513:data<=16'd1057;
      25514:data<=16'd1274;
      25515:data<=16'd1400;
      25516:data<=16'd1287;
      25517:data<=16'd1256;
      25518:data<=16'd1489;
      25519:data<=16'd1400;
      25520:data<=16'd1489;
      25521:data<=16'd552;
      25522:data<=-16'd1234;
      25523:data<=-16'd1077;
      25524:data<=-16'd593;
      25525:data<=-16'd529;
      25526:data<=16'd299;
      25527:data<=16'd64;
      25528:data<=16'd102;
      25529:data<=16'd550;
      25530:data<=-16'd344;
      25531:data<=16'd355;
      25532:data<=16'd596;
      25533:data<=-16'd629;
      25534:data<=16'd240;
      25535:data<=-16'd4240;
      25536:data<=-16'd13706;
      25537:data<=-16'd14989;
      25538:data<=-16'd12000;
      25539:data<=-16'd12286;
      25540:data<=-16'd11782;
      25541:data<=-16'd11051;
      25542:data<=-16'd11106;
      25543:data<=-16'd10369;
      25544:data<=-16'd10053;
      25545:data<=-16'd9324;
      25546:data<=-16'd8934;
      25547:data<=-16'd9911;
      25548:data<=-16'd9741;
      25549:data<=-16'd9213;
      25550:data<=-16'd8863;
      25551:data<=-16'd7644;
      25552:data<=-16'd7181;
      25553:data<=-16'd7025;
      25554:data<=-16'd6495;
      25555:data<=-16'd6093;
      25556:data<=-16'd4919;
      25557:data<=-16'd4091;
      25558:data<=-16'd3759;
      25559:data<=-16'd2793;
      25560:data<=-16'd2830;
      25561:data<=-16'd3093;
      25562:data<=-16'd1739;
      25563:data<=-16'd346;
      25564:data<=-16'd64;
      25565:data<=-16'd291;
      25566:data<=16'd92;
      25567:data<=16'd775;
      25568:data<=16'd804;
      25569:data<=16'd1087;
      25570:data<=16'd1577;
      25571:data<=16'd2397;
      25572:data<=16'd3864;
      25573:data<=16'd4029;
      25574:data<=16'd3858;
      25575:data<=16'd4267;
      25576:data<=16'd3767;
      25577:data<=16'd3849;
      25578:data<=16'd3930;
      25579:data<=16'd3594;
      25580:data<=16'd4619;
      25581:data<=16'd4115;
      25582:data<=16'd3730;
      25583:data<=16'd5116;
      25584:data<=16'd3956;
      25585:data<=16'd7752;
      25586:data<=16'd17995;
      25587:data<=16'd20069;
      25588:data<=16'd17105;
      25589:data<=16'd17807;
      25590:data<=16'd17086;
      25591:data<=16'd16175;
      25592:data<=16'd16598;
      25593:data<=16'd15302;
      25594:data<=16'd15145;
      25595:data<=16'd15201;
      25596:data<=16'd14175;
      25597:data<=16'd15057;
      25598:data<=16'd15412;
      25599:data<=16'd14575;
      25600:data<=16'd14665;
      25601:data<=16'd13873;
      25602:data<=16'd12772;
      25603:data<=16'd12625;
      25604:data<=16'd12254;
      25605:data<=16'd11677;
      25606:data<=16'd10977;
      25607:data<=16'd10191;
      25608:data<=16'd9662;
      25609:data<=16'd10003;
      25610:data<=16'd11309;
      25611:data<=16'd11362;
      25612:data<=16'd10307;
      25613:data<=16'd10049;
      25614:data<=16'd9718;
      25615:data<=16'd9401;
      25616:data<=16'd9236;
      25617:data<=16'd8442;
      25618:data<=16'd8172;
      25619:data<=16'd7947;
      25620:data<=16'd7021;
      25621:data<=16'd7172;
      25622:data<=16'd8385;
      25623:data<=16'd8825;
      25624:data<=16'd8109;
      25625:data<=16'd7847;
      25626:data<=16'd7953;
      25627:data<=16'd6963;
      25628:data<=16'd6576;
      25629:data<=16'd5926;
      25630:data<=16'd3836;
      25631:data<=16'd4094;
      25632:data<=16'd3896;
      25633:data<=16'd2431;
      25634:data<=16'd5421;
      25635:data<=16'd3802;
      25636:data<=-16'd6308;
      25637:data<=-16'd9571;
      25638:data<=-16'd6587;
      25639:data<=-16'd7050;
      25640:data<=-16'd7398;
      25641:data<=-16'd7021;
      25642:data<=-16'd7438;
      25643:data<=-16'd6534;
      25644:data<=-16'd6501;
      25645:data<=-16'd7269;
      25646:data<=-16'd6155;
      25647:data<=-16'd4296;
      25648:data<=-16'd3163;
      25649:data<=-16'd3187;
      25650:data<=-16'd3245;
      25651:data<=-16'd2613;
      25652:data<=-16'd2776;
      25653:data<=-16'd3168;
      25654:data<=-16'd2890;
      25655:data<=-16'd2563;
      25656:data<=-16'd2124;
      25657:data<=-16'd2050;
      25658:data<=-16'd1986;
      25659:data<=-16'd839;
      25660:data<=16'd685;
      25661:data<=16'd1283;
      25662:data<=16'd719;
      25663:data<=16'd564;
      25664:data<=16'd746;
      25665:data<=-16'd123;
      25666:data<=-16'd86;
      25667:data<=16'd494;
      25668:data<=-16'd349;
      25669:data<=-16'd505;
      25670:data<=-16'd224;
      25671:data<=16'd138;
      25672:data<=16'd1953;
      25673:data<=16'd2575;
      25674:data<=16'd2067;
      25675:data<=16'd2053;
      25676:data<=16'd1325;
      25677:data<=16'd1365;
      25678:data<=16'd1665;
      25679:data<=16'd1347;
      25680:data<=16'd1791;
      25681:data<=16'd746;
      25682:data<=16'd388;
      25683:data<=16'd1601;
      25684:data<=16'd183;
      25685:data<=16'd4090;
      25686:data<=16'd14111;
      25687:data<=16'd16375;
      25688:data<=16'd14031;
      25689:data<=16'd14223;
      25690:data<=16'd13100;
      25691:data<=16'd12326;
      25692:data<=16'd12214;
      25693:data<=16'd10857;
      25694:data<=16'd10655;
      25695:data<=16'd10539;
      25696:data<=16'd11245;
      25697:data<=16'd13212;
      25698:data<=16'd12554;
      25699:data<=16'd11526;
      25700:data<=16'd11664;
      25701:data<=16'd10757;
      25702:data<=16'd10307;
      25703:data<=16'd9846;
      25704:data<=16'd8772;
      25705:data<=16'd8316;
      25706:data<=16'd7603;
      25707:data<=16'd7068;
      25708:data<=16'd6517;
      25709:data<=16'd6158;
      25710:data<=16'd7445;
      25711:data<=16'd7626;
      25712:data<=16'd6587;
      25713:data<=16'd6510;
      25714:data<=16'd6012;
      25715:data<=16'd5770;
      25716:data<=16'd5262;
      25717:data<=16'd3717;
      25718:data<=16'd3914;
      25719:data<=16'd4071;
      25720:data<=16'd3200;
      25721:data<=16'd3647;
      25722:data<=16'd4100;
      25723:data<=16'd4673;
      25724:data<=16'd5033;
      25725:data<=16'd4009;
      25726:data<=16'd3694;
      25727:data<=16'd2892;
      25728:data<=16'd1798;
      25729:data<=16'd2165;
      25730:data<=16'd1469;
      25731:data<=16'd1290;
      25732:data<=16'd1310;
      25733:data<=-16'd130;
      25734:data<=16'd1844;
      25735:data<=16'd1048;
      25736:data<=-16'd7732;
      25737:data<=-16'd12076;
      25738:data<=-16'd10534;
      25739:data<=-16'd10740;
      25740:data<=-16'd10696;
      25741:data<=-16'd10534;
      25742:data<=-16'd10900;
      25743:data<=-16'd10009;
      25744:data<=-16'd9671;
      25745:data<=-16'd9696;
      25746:data<=-16'd9291;
      25747:data<=-16'd8567;
      25748:data<=-16'd7072;
      25749:data<=-16'd6573;
      25750:data<=-16'd6664;
      25751:data<=-16'd6552;
      25752:data<=-16'd7142;
      25753:data<=-16'd6777;
      25754:data<=-16'd6326;
      25755:data<=-16'd6666;
      25756:data<=-16'd5802;
      25757:data<=-16'd5532;
      25758:data<=-16'd5924;
      25759:data<=-16'd5413;
      25760:data<=-16'd5612;
      25761:data<=-16'd5344;
      25762:data<=-16'd4751;
      25763:data<=-16'd6117;
      25764:data<=-16'd7363;
      25765:data<=-16'd7476;
      25766:data<=-16'd7012;
      25767:data<=-16'd6220;
      25768:data<=-16'd6466;
      25769:data<=-16'd6546;
      25770:data<=-16'd6000;
      25771:data<=-16'd6284;
      25772:data<=-16'd6862;
      25773:data<=-16'd7870;
      25774:data<=-16'd8229;
      25775:data<=-16'd7112;
      25776:data<=-16'd7048;
      25777:data<=-16'd7313;
      25778:data<=-16'd6902;
      25779:data<=-16'd7047;
      25780:data<=-16'd6717;
      25781:data<=-16'd6514;
      25782:data<=-16'd6173;
      25783:data<=-16'd5021;
      25784:data<=-16'd6435;
      25785:data<=-16'd5981;
      25786:data<=16'd1469;
      25787:data<=16'd6983;
      25788:data<=16'd6369;
      25789:data<=16'd5456;
      25790:data<=16'd5109;
      25791:data<=16'd4955;
      25792:data<=16'd5154;
      25793:data<=16'd4337;
      25794:data<=16'd3961;
      25795:data<=16'd4369;
      25796:data<=16'd4027;
      25797:data<=16'd3118;
      25798:data<=16'd1673;
      25799:data<=16'd987;
      25800:data<=16'd1663;
      25801:data<=16'd1381;
      25802:data<=16'd667;
      25803:data<=16'd969;
      25804:data<=16'd1037;
      25805:data<=16'd848;
      25806:data<=16'd754;
      25807:data<=16'd490;
      25808:data<=16'd402;
      25809:data<=-16'd305;
      25810:data<=-16'd1929;
      25811:data<=-16'd2927;
      25812:data<=-16'd2514;
      25813:data<=-16'd1741;
      25814:data<=-16'd2041;
      25815:data<=-16'd2743;
      25816:data<=-16'd2717;
      25817:data<=-16'd2461;
      25818:data<=-16'd2012;
      25819:data<=-16'd1829;
      25820:data<=-16'd1868;
      25821:data<=-16'd1246;
      25822:data<=-16'd2187;
      25823:data<=-16'd4137;
      25824:data<=-16'd3539;
      25825:data<=-16'd2767;
      25826:data<=-16'd3186;
      25827:data<=-16'd2886;
      25828:data<=-16'd3157;
      25829:data<=-16'd3101;
      25830:data<=-16'd1709;
      25831:data<=-16'd1033;
      25832:data<=-16'd740;
      25833:data<=-16'd896;
      25834:data<=-16'd1266;
      25835:data<=-16'd2776;
      25836:data<=-16'd9643;
      25837:data<=-16'd16311;
      25838:data<=-16'd16046;
      25839:data<=-16'd14922;
      25840:data<=-16'd15032;
      25841:data<=-16'd13855;
      25842:data<=-16'd13464;
      25843:data<=-16'd12807;
      25844:data<=-16'd11761;
      25845:data<=-16'd11626;
      25846:data<=-16'd10502;
      25847:data<=-16'd10622;
      25848:data<=-16'd12395;
      25849:data<=-16'd11947;
      25850:data<=-16'd10953;
      25851:data<=-16'd10860;
      25852:data<=-16'd10458;
      25853:data<=-16'd10214;
      25854:data<=-16'd9561;
      25855:data<=-16'd8904;
      25856:data<=-16'd8780;
      25857:data<=-16'd7794;
      25858:data<=-16'd6696;
      25859:data<=-16'd6699;
      25860:data<=-16'd7649;
      25861:data<=-16'd8307;
      25862:data<=-16'd7500;
      25863:data<=-16'd7166;
      25864:data<=-16'd7401;
      25865:data<=-16'd6404;
      25866:data<=-16'd6023;
      25867:data<=-16'd6337;
      25868:data<=-16'd5894;
      25869:data<=-16'd5673;
      25870:data<=-16'd5225;
      25871:data<=-16'd4623;
      25872:data<=-16'd5239;
      25873:data<=-16'd6537;
      25874:data<=-16'd7068;
      25875:data<=-16'd6037;
      25876:data<=-16'd5627;
      25877:data<=-16'd6285;
      25878:data<=-16'd5125;
      25879:data<=-16'd4249;
      25880:data<=-16'd4589;
      25881:data<=-16'd3817;
      25882:data<=-16'd3720;
      25883:data<=-16'd2902;
      25884:data<=-16'd2129;
      25885:data<=-16'd4775;
      25886:data<=-16'd1389;
      25887:data<=16'd8340;
      25888:data<=16'd10088;
      25889:data<=16'd7680;
      25890:data<=16'd8772;
      25891:data<=16'd8273;
      25892:data<=16'd7591;
      25893:data<=16'd8343;
      25894:data<=16'd7354;
      25895:data<=16'd7036;
      25896:data<=16'd7121;
      25897:data<=16'd4930;
      25898:data<=16'd2740;
      25899:data<=16'd2049;
      25900:data<=16'd2244;
      25901:data<=16'd2564;
      25902:data<=16'd2637;
      25903:data<=16'd2723;
      25904:data<=16'd2517;
      25905:data<=16'd2532;
      25906:data<=16'd2444;
      25907:data<=16'd1692;
      25908:data<=16'd1947;
      25909:data<=16'd1794;
      25910:data<=-16'd138;
      25911:data<=-16'd811;
      25912:data<=-16'd328;
      25913:data<=-16'd276;
      25914:data<=16'd77;
      25915:data<=16'd153;
      25916:data<=16'd94;
      25917:data<=16'd785;
      25918:data<=16'd1259;
      25919:data<=16'd914;
      25920:data<=16'd702;
      25921:data<=16'd1266;
      25922:data<=16'd741;
      25923:data<=-16'd1113;
      25924:data<=-16'd1416;
      25925:data<=-16'd767;
      25926:data<=-16'd64;
      25927:data<=16'd1066;
      25928:data<=16'd473;
      25929:data<=-16'd284;
      25930:data<=16'd449;
      25931:data<=16'd493;
      25932:data<=16'd829;
      25933:data<=16'd265;
      25934:data<=-16'd1158;
      25935:data<=16'd144;
      25936:data<=-16'd3441;
      25937:data<=-16'd13400;
      25938:data<=-16'd16075;
      25939:data<=-16'd13069;
      25940:data<=-16'd12959;
      25941:data<=-16'd12214;
      25942:data<=-16'd10860;
      25943:data<=-16'd10972;
      25944:data<=-16'd10398;
      25945:data<=-16'd9919;
      25946:data<=-16'd9479;
      25947:data<=-16'd9113;
      25948:data<=-16'd10122;
      25949:data<=-16'd10009;
      25950:data<=-16'd8790;
      25951:data<=-16'd8705;
      25952:data<=-16'd8301;
      25953:data<=-16'd7379;
      25954:data<=-16'd6863;
      25955:data<=-16'd6038;
      25956:data<=-16'd5350;
      25957:data<=-16'd5095;
      25958:data<=-16'd4461;
      25959:data<=-16'd3580;
      25960:data<=-16'd2881;
      25961:data<=-16'd2419;
      25962:data<=-16'd2391;
      25963:data<=-16'd2052;
      25964:data<=-16'd373;
      25965:data<=16'd981;
      25966:data<=16'd870;
      25967:data<=16'd1118;
      25968:data<=16'd1384;
      25969:data<=16'd995;
      25970:data<=16'd1274;
      25971:data<=16'd1342;
      25972:data<=16'd1721;
      25973:data<=16'd3617;
      25974:data<=16'd4341;
      25975:data<=16'd3858;
      25976:data<=16'd3550;
      25977:data<=16'd2969;
      25978:data<=16'd3753;
      25979:data<=16'd4752;
      25980:data<=16'd4217;
      25981:data<=16'd4156;
      25982:data<=16'd3971;
      25983:data<=16'd4338;
      25984:data<=16'd5210;
      25985:data<=16'd4047;
      25986:data<=16'd8234;
      25987:data<=16'd18330;
      25988:data<=16'd20882;
      25989:data<=16'd18327;
      25990:data<=16'd18766;
      25991:data<=16'd17992;
      25992:data<=16'd17036;
      25993:data<=16'd17509;
      25994:data<=16'd16075;
      25995:data<=16'd15151;
      25996:data<=16'd15062;
      25997:data<=16'd14640;
      25998:data<=16'd15837;
      25999:data<=16'd16169;
      26000:data<=16'd14778;
      26001:data<=16'd14064;
      26002:data<=16'd13482;
      26003:data<=16'd13538;
      26004:data<=16'd13863;
      26005:data<=16'd12690;
      26006:data<=16'd11389;
      26007:data<=16'd10947;
      26008:data<=16'd10646;
      26009:data<=16'd9867;
      26010:data<=16'd9635;
      26011:data<=16'd11051;
      26012:data<=16'd11433;
      26013:data<=16'd10316;
      26014:data<=16'd9868;
      26015:data<=16'd9321;
      26016:data<=16'd9339;
      26017:data<=16'd9659;
      26018:data<=16'd8613;
      26019:data<=16'd8420;
      26020:data<=16'd8067;
      26021:data<=16'd6341;
      26022:data<=16'd7069;
      26023:data<=16'd9003;
      26024:data<=16'd9045;
      26025:data<=16'd8526;
      26026:data<=16'd8334;
      26027:data<=16'd8087;
      26028:data<=16'd7312;
      26029:data<=16'd7081;
      26030:data<=16'd6702;
      26031:data<=16'd4461;
      26032:data<=16'd3941;
      26033:data<=16'd3833;
      26034:data<=16'd2006;
      26035:data<=16'd4131;
      26036:data<=16'd3401;
      26037:data<=-16'd5718;
      26038:data<=-16'd9690;
      26039:data<=-16'd8043;
      26040:data<=-16'd8872;
      26041:data<=-16'd7940;
      26042:data<=-16'd6910;
      26043:data<=-16'd8425;
      26044:data<=-16'd8029;
      26045:data<=-16'd7421;
      26046:data<=-16'd7782;
      26047:data<=-16'd6771;
      26048:data<=-16'd5286;
      26049:data<=-16'd4293;
      26050:data<=-16'd3949;
      26051:data<=-16'd3485;
      26052:data<=-16'd3333;
      26053:data<=-16'd4228;
      26054:data<=-16'd3668;
      26055:data<=-16'd2792;
      26056:data<=-16'd3297;
      26057:data<=-16'd2757;
      26058:data<=-16'd2497;
      26059:data<=-16'd2870;
      26060:data<=-16'd1218;
      26061:data<=16'd793;
      26062:data<=16'd1322;
      26063:data<=16'd735;
      26064:data<=16'd277;
      26065:data<=16'd582;
      26066:data<=16'd168;
      26067:data<=16'd2;
      26068:data<=16'd502;
      26069:data<=16'd153;
      26070:data<=16'd209;
      26071:data<=16'd59;
      26072:data<=-16'd226;
      26073:data<=16'd1313;
      26074:data<=16'd2043;
      26075:data<=16'd1519;
      26076:data<=16'd1239;
      26077:data<=16'd511;
      26078:data<=16'd785;
      26079:data<=16'd1052;
      26080:data<=16'd602;
      26081:data<=16'd961;
      26082:data<=-16'd23;
      26083:data<=-16'd265;
      26084:data<=16'd734;
      26085:data<=-16'd578;
      26086:data<=16'd3486;
      26087:data<=16'd13254;
      26088:data<=16'd16211;
      26089:data<=16'd14468;
      26090:data<=16'd14085;
      26091:data<=16'd12847;
      26092:data<=16'd12020;
      26093:data<=16'd12116;
      26094:data<=16'd12066;
      26095:data<=16'd12070;
      26096:data<=16'd10712;
      26097:data<=16'd10257;
      26098:data<=16'd12395;
      26099:data<=16'd13452;
      26100:data<=16'd12790;
      26101:data<=16'd11776;
      26102:data<=16'd10392;
      26103:data<=16'd9843;
      26104:data<=16'd10026;
      26105:data<=16'd9115;
      26106:data<=16'd7591;
      26107:data<=16'd6945;
      26108:data<=16'd6276;
      26109:data<=16'd5318;
      26110:data<=16'd5776;
      26111:data<=16'd6869;
      26112:data<=16'd7185;
      26113:data<=16'd6968;
      26114:data<=16'd5965;
      26115:data<=16'd5131;
      26116:data<=16'd5110;
      26117:data<=16'd4933;
      26118:data<=16'd4969;
      26119:data<=16'd4534;
      26120:data<=16'd3130;
      26121:data<=16'd2663;
      26122:data<=16'd3099;
      26123:data<=16'd3923;
      26124:data<=16'd4874;
      26125:data<=16'd4646;
      26126:data<=16'd4202;
      26127:data<=16'd3961;
      26128:data<=16'd3109;
      26129:data<=16'd2907;
      26130:data<=16'd2811;
      26131:data<=16'd2112;
      26132:data<=16'd2106;
      26133:data<=16'd1307;
      26134:data<=16'd187;
      26135:data<=16'd1698;
      26136:data<=16'd1107;
      26137:data<=-16'd5844;
      26138:data<=-16'd11685;
      26139:data<=-16'd11650;
      26140:data<=-16'd10909;
      26141:data<=-16'd10939;
      26142:data<=-16'd10170;
      26143:data<=-16'd10207;
      26144:data<=-16'd10404;
      26145:data<=-16'd10017;
      26146:data<=-16'd10187;
      26147:data<=-16'd9797;
      26148:data<=-16'd8739;
      26149:data<=-16'd7767;
      26150:data<=-16'd6895;
      26151:data<=-16'd7098;
      26152:data<=-16'd7142;
      26153:data<=-16'd6590;
      26154:data<=-16'd6993;
      26155:data<=-16'd6652;
      26156:data<=-16'd5815;
      26157:data<=-16'd6150;
      26158:data<=-16'd5812;
      26159:data<=-16'd5153;
      26160:data<=-16'd5145;
      26161:data<=-16'd4927;
      26162:data<=-16'd5022;
      26163:data<=-16'd5089;
      26164:data<=-16'd5510;
      26165:data<=-16'd6819;
      26166:data<=-16'd7063;
      26167:data<=-16'd6977;
      26168:data<=-16'd7332;
      26169:data<=-16'd6649;
      26170:data<=-16'd6117;
      26171:data<=-16'd6105;
      26172:data<=-16'd5946;
      26173:data<=-16'd6919;
      26174:data<=-16'd8422;
      26175:data<=-16'd8831;
      26176:data<=-16'd8264;
      26177:data<=-16'd7862;
      26178:data<=-16'd8199;
      26179:data<=-16'd8281;
      26180:data<=-16'd7984;
      26181:data<=-16'd7843;
      26182:data<=-16'd7899;
      26183:data<=-16'd7817;
      26184:data<=-16'd6699;
      26185:data<=-16'd7001;
      26186:data<=-16'd7887;
      26187:data<=-16'd2317;
      26188:data<=16'd4881;
      26189:data<=16'd5080;
      26190:data<=16'd3891;
      26191:data<=16'd4341;
      26192:data<=16'd3444;
      26193:data<=16'd3389;
      26194:data<=16'd3853;
      26195:data<=16'd3309;
      26196:data<=16'd3292;
      26197:data<=16'd3060;
      26198:data<=16'd1924;
      26199:data<=16'd431;
      26200:data<=-16'd431;
      26201:data<=16'd32;
      26202:data<=-16'd76;
      26203:data<=-16'd535;
      26204:data<=-16'd161;
      26205:data<=-16'd428;
      26206:data<=-16'd940;
      26207:data<=-16'd1192;
      26208:data<=-16'd1278;
      26209:data<=-16'd644;
      26210:data<=-16'd1407;
      26211:data<=-16'd3397;
      26212:data<=-16'd4064;
      26213:data<=-16'd4124;
      26214:data<=-16'd3795;
      26215:data<=-16'd3342;
      26216:data<=-16'd3660;
      26217:data<=-16'd3670;
      26218:data<=-16'd3521;
      26219:data<=-16'd3307;
      26220:data<=-16'd3099;
      26221:data<=-16'd3657;
      26222:data<=-16'd3351;
      26223:data<=-16'd3432;
      26224:data<=-16'd4904;
      26225:data<=-16'd4523;
      26226:data<=-16'd4215;
      26227:data<=-16'd4728;
      26228:data<=-16'd3257;
      26229:data<=-16'd3110;
      26230:data<=-16'd3902;
      26231:data<=-16'd2732;
      26232:data<=-16'd2247;
      26233:data<=-16'd1544;
      26234:data<=-16'd790;
      26235:data<=-16'd1770;
      26236:data<=-16'd2558;
      26237:data<=-16'd7485;
      26238:data<=-16'd15456;
      26239:data<=-16'd16416;
      26240:data<=-16'd14114;
      26241:data<=-16'd14331;
      26242:data<=-16'd13520;
      26243:data<=-16'd12866;
      26244:data<=-16'd12797;
      26245:data<=-16'd11729;
      26246:data<=-16'd11702;
      26247:data<=-16'd11315;
      26248:data<=-16'd10822;
      26249:data<=-16'd12380;
      26250:data<=-16'd12624;
      26251:data<=-16'd11351;
      26252:data<=-16'd10934;
      26253:data<=-16'd10173;
      26254:data<=-16'd9770;
      26255:data<=-16'd9902;
      26256:data<=-16'd8666;
      26257:data<=-16'd7582;
      26258:data<=-16'd7526;
      26259:data<=-16'd6666;
      26260:data<=-16'd6102;
      26261:data<=-16'd7406;
      26262:data<=-16'd8179;
      26263:data<=-16'd7512;
      26264:data<=-16'd7275;
      26265:data<=-16'd6698;
      26266:data<=-16'd5789;
      26267:data<=-16'd6132;
      26268:data<=-16'd6181;
      26269:data<=-16'd5618;
      26270:data<=-16'd5227;
      26271:data<=-16'd3997;
      26272:data<=-16'd3268;
      26273:data<=-16'd3971;
      26274:data<=-16'd5321;
      26275:data<=-16'd6563;
      26276:data<=-16'd5694;
      26277:data<=-16'd4842;
      26278:data<=-16'd5691;
      26279:data<=-16'd4905;
      26280:data<=-16'd4558;
      26281:data<=-16'd5251;
      26282:data<=-16'd3712;
      26283:data<=-16'd3312;
      26284:data<=-16'd3001;
      26285:data<=-16'd1715;
      26286:data<=-16'd4243;
      26287:data<=-16'd1930;
      26288:data<=16'd7899;
      26289:data<=16'd10337;
      26290:data<=16'd7829;
      26291:data<=16'd9389;
      26292:data<=16'd9456;
      26293:data<=16'd8170;
      26294:data<=16'd8384;
      26295:data<=16'd7511;
      26296:data<=16'd7711;
      26297:data<=16'd8834;
      26298:data<=16'd7009;
      26299:data<=16'd4222;
      26300:data<=16'd3418;
      26301:data<=16'd3782;
      26302:data<=16'd3803;
      26303:data<=16'd3585;
      26304:data<=16'd3751;
      26305:data<=16'd3883;
      26306:data<=16'd3842;
      26307:data<=16'd3482;
      26308:data<=16'd3077;
      26309:data<=16'd3389;
      26310:data<=16'd3109;
      26311:data<=16'd1701;
      26312:data<=16'd617;
      26313:data<=16'd585;
      26314:data<=16'd1468;
      26315:data<=16'd1579;
      26316:data<=16'd1087;
      26317:data<=16'd1663;
      26318:data<=16'd1736;
      26319:data<=16'd1777;
      26320:data<=16'd2497;
      26321:data<=16'd1651;
      26322:data<=16'd1444;
      26323:data<=16'd2047;
      26324:data<=16'd475;
      26325:data<=-16'd146;
      26326:data<=16'd591;
      26327:data<=16'd525;
      26328:data<=16'd1354;
      26329:data<=16'd1926;
      26330:data<=16'd1841;
      26331:data<=16'd2003;
      26332:data<=16'd1468;
      26333:data<=16'd2009;
      26334:data<=16'd2074;
      26335:data<=16'd1239;
      26336:data<=16'd2491;
      26337:data<=-16'd1645;
      26338:data<=-16'd11226;
      26339:data<=-16'd13540;
      26340:data<=-16'd11433;
      26341:data<=-16'd11509;
      26342:data<=-16'd10745;
      26343:data<=-16'd10258;
      26344:data<=-16'd9902;
      26345:data<=-16'd8628;
      26346:data<=-16'd8689;
      26347:data<=-16'd7893;
      26348:data<=-16'd6953;
      26349:data<=-16'd8249;
      26350:data<=-16'd8298;
      26351:data<=-16'd7415;
      26352:data<=-16'd7473;
      26353:data<=-16'd7095;
      26354:data<=-16'd6793;
      26355:data<=-16'd6341;
      26356:data<=-16'd5394;
      26357:data<=-16'd4889;
      26358:data<=-16'd4454;
      26359:data<=-16'd4185;
      26360:data<=-16'd3679;
      26361:data<=-16'd2726;
      26362:data<=-16'd2096;
      26363:data<=-16'd1290;
      26364:data<=-16'd1304;
      26365:data<=-16'd1568;
      26366:data<=16'd124;
      26367:data<=16'd1171;
      26368:data<=16'd767;
      26369:data<=16'd837;
      26370:data<=16'd804;
      26371:data<=16'd1519;
      26372:data<=16'd2331;
      26373:data<=16'd2265;
      26374:data<=16'd3597;
      26375:data<=16'd4610;
      26376:data<=16'd4199;
      26377:data<=16'd4557;
      26378:data<=16'd4417;
      26379:data<=16'd3991;
      26380:data<=16'd4229;
      26381:data<=16'd4102;
      26382:data<=16'd4343;
      26383:data<=16'd4455;
      26384:data<=16'd4590;
      26385:data<=16'd4416;
      26386:data<=16'd3186;
      26387:data<=16'd8103;
      26388:data<=16'd17837;
      26389:data<=16'd20052;
      26390:data<=16'd17929;
      26391:data<=16'd18122;
      26392:data<=16'd17226;
      26393:data<=16'd16343;
      26394:data<=16'd16125;
      26395:data<=16'd15303;
      26396:data<=16'd15594;
      26397:data<=16'd14736;
      26398:data<=16'd13476;
      26399:data<=16'd14950;
      26400:data<=16'd15626;
      26401:data<=16'd14643;
      26402:data<=16'd14164;
      26403:data<=16'd13635;
      26404:data<=16'd13238;
      26405:data<=16'd12765;
      26406:data<=16'd12239;
      26407:data<=16'd12022;
      26408:data<=16'd11590;
      26409:data<=16'd11424;
      26410:data<=16'd10566;
      26411:data<=16'd9697;
      26412:data<=16'd11041;
      26413:data<=16'd11385;
      26414:data<=16'd10285;
      26415:data<=16'd10662;
      26416:data<=16'd10243;
      26417:data<=16'd9100;
      26418:data<=16'd9301;
      26419:data<=16'd9297;
      26420:data<=16'd8965;
      26421:data<=16'd8320;
      26422:data<=16'd7169;
      26423:data<=16'd7207;
      26424:data<=16'd8287;
      26425:data<=16'd8942;
      26426:data<=16'd8317;
      26427:data<=16'd7564;
      26428:data<=16'd7968;
      26429:data<=16'd7603;
      26430:data<=16'd6942;
      26431:data<=16'd7021;
      26432:data<=16'd5823;
      26433:data<=16'd4661;
      26434:data<=16'd3530;
      26435:data<=16'd2473;
      26436:data<=16'd4955;
      26437:data<=16'd3968;
      26438:data<=-16'd4605;
      26439:data<=-16'd8757;
      26440:data<=-16'd7010;
      26441:data<=-16'd7163;
      26442:data<=-16'd7119;
      26443:data<=-16'd6241;
      26444:data<=-16'd6686;
      26445:data<=-16'd6536;
      26446:data<=-16'd6269;
      26447:data<=-16'd6648;
      26448:data<=-16'd5982;
      26449:data<=-16'd4299;
      26450:data<=-16'd3151;
      26451:data<=-16'd3227;
      26452:data<=-16'd3277;
      26453:data<=-16'd2955;
      26454:data<=-16'd3146;
      26455:data<=-16'd2913;
      26456:data<=-16'd2590;
      26457:data<=-16'd3218;
      26458:data<=-16'd3297;
      26459:data<=-16'd2804;
      26460:data<=-16'd2687;
      26461:data<=-16'd1768;
      26462:data<=16'd97;
      26463:data<=16'd1131;
      26464:data<=16'd810;
      26465:data<=16'd343;
      26466:data<=-16'd2;
      26467:data<=-16'd344;
      26468:data<=-16'd117;
      26469:data<=-16'd273;
      26470:data<=-16'd714;
      26471:data<=-16'd150;
      26472:data<=-16'd100;
      26473:data<=-16'd230;
      26474:data<=16'd1093;
      26475:data<=16'd2012;
      26476:data<=16'd2103;
      26477:data<=16'd2005;
      26478:data<=16'd1609;
      26479:data<=16'd1635;
      26480:data<=16'd1089;
      26481:data<=16'd902;
      26482:data<=16'd1924;
      26483:data<=16'd1174;
      26484:data<=16'd920;
      26485:data<=16'd1726;
      26486:data<=16'd144;
      26487:data<=16'd3338;
      26488:data<=16'd12283;
      26489:data<=16'd15609;
      26490:data<=16'd14835;
      26491:data<=16'd15417;
      26492:data<=16'd14795;
      26493:data<=16'd14231;
      26494:data<=16'd14148;
      26495:data<=16'd13022;
      26496:data<=16'd12869;
      26497:data<=16'd12610;
      26498:data<=16'd11496;
      26499:data<=16'd11697;
      26500:data<=16'd12110;
      26501:data<=16'd11711;
      26502:data<=16'd11139;
      26503:data<=16'd10246;
      26504:data<=16'd9495;
      26505:data<=16'd9218;
      26506:data<=16'd8886;
      26507:data<=16'd8144;
      26508:data<=16'd7741;
      26509:data<=16'd7884;
      26510:data<=16'd7204;
      26511:data<=16'd6845;
      26512:data<=16'd7829;
      26513:data<=16'd7787;
      26514:data<=16'd6983;
      26515:data<=16'd6652;
      26516:data<=16'd5891;
      26517:data<=16'd5278;
      26518:data<=16'd5106;
      26519:data<=16'd5181;
      26520:data<=16'd5421;
      26521:data<=16'd4531;
      26522:data<=16'd3535;
      26523:data<=16'd3398;
      26524:data<=16'd3385;
      26525:data<=16'd4394;
      26526:data<=16'd5007;
      26527:data<=16'd4040;
      26528:data<=16'd3832;
      26529:data<=16'd3755;
      26530:data<=16'd3083;
      26531:data<=16'd2693;
      26532:data<=16'd1956;
      26533:data<=16'd2087;
      26534:data<=16'd2117;
      26535:data<=16'd732;
      26536:data<=16'd1858;
      26537:data<=16'd2494;
      26538:data<=-16'd3083;
      26539:data<=-16'd8545;
      26540:data<=-16'd8784;
      26541:data<=-16'd7937;
      26542:data<=-16'd8237;
      26543:data<=-16'd8490;
      26544:data<=-16'd8137;
      26545:data<=-16'd7935;
      26546:data<=-16'd8149;
      26547:data<=-16'd7984;
      26548:data<=-16'd7938;
      26549:data<=-16'd7506;
      26550:data<=-16'd5749;
      26551:data<=-16'd5009;
      26552:data<=-16'd5615;
      26553:data<=-16'd5215;
      26554:data<=-16'd4777;
      26555:data<=-16'd5586;
      26556:data<=-16'd6109;
      26557:data<=-16'd5688;
      26558:data<=-16'd5564;
      26559:data<=-16'd5964;
      26560:data<=-16'd6082;
      26561:data<=-16'd6273;
      26562:data<=-16'd6061;
      26563:data<=-16'd4772;
      26564:data<=-16'd4575;
      26565:data<=-16'd5288;
      26566:data<=-16'd4643;
      26567:data<=-16'd4444;
      26568:data<=-16'd5310;
      26569:data<=-16'd5325;
      26570:data<=-16'd5297;
      26571:data<=-16'd5588;
      26572:data<=-16'd5614;
      26573:data<=-16'd5818;
      26574:data<=-16'd6047;
      26575:data<=-16'd6818;
      26576:data<=-16'd7589;
      26577:data<=-16'd6907;
      26578:data<=-16'd6614;
      26579:data<=-16'd7253;
      26580:data<=-16'd7028;
      26581:data<=-16'd6479;
      26582:data<=-16'd5953;
      26583:data<=-16'd5912;
      26584:data<=-16'd6551;
      26585:data<=-16'd6138;
      26586:data<=-16'd6878;
      26587:data<=-16'd8675;
      26588:data<=-16'd4599;
      26589:data<=16'd2350;
      26590:data<=16'd3196;
      26591:data<=16'd1468;
      26592:data<=16'd2234;
      26593:data<=16'd2434;
      26594:data<=16'd1609;
      26595:data<=16'd1653;
      26596:data<=16'd1441;
      26597:data<=16'd914;
      26598:data<=16'd881;
      26599:data<=16'd73;
      26600:data<=-16'd1538;
      26601:data<=-16'd2228;
      26602:data<=-16'd2106;
      26603:data<=-16'd2033;
      26604:data<=-16'd2194;
      26605:data<=-16'd2560;
      26606:data<=-16'd2215;
      26607:data<=-16'd1597;
      26608:data<=-16'd2261;
      26609:data<=-16'd2998;
      26610:data<=-16'd2870;
      26611:data<=-16'd3193;
      26612:data<=-16'd4131;
      26613:data<=-16'd5113;
      26614:data<=-16'd5435;
      26615:data<=-16'd5075;
      26616:data<=-16'd5115;
      26617:data<=-16'd4871;
      26618:data<=-16'd4338;
      26619:data<=-16'd4563;
      26620:data<=-16'd4387;
      26621:data<=-16'd4441;
      26622:data<=-16'd5009;
      26623:data<=-16'd4235;
      26624:data<=-16'd4787;
      26625:data<=-16'd7013;
      26626:data<=-16'd6846;
      26627:data<=-16'd6213;
      26628:data<=-16'd6719;
      26629:data<=-16'd6443;
      26630:data<=-16'd6304;
      26631:data<=-16'd6020;
      26632:data<=-16'd5595;
      26633:data<=-16'd6035;
      26634:data<=-16'd5692;
      26635:data<=-16'd6002;
      26636:data<=-16'd6787;
      26637:data<=-16'd5862;
      26638:data<=-16'd9273;
      26639:data<=-16'd16533;
      26640:data<=-16'd18057;
      26641:data<=-16'd16143;
      26642:data<=-16'd16031;
      26643:data<=-16'd15611;
      26644:data<=-16'd14850;
      26645:data<=-16'd14081;
      26646:data<=-16'd13694;
      26647:data<=-16'd14292;
      26648:data<=-16'd13379;
      26649:data<=-16'd12798;
      26650:data<=-16'd14431;
      26651:data<=-16'd14041;
      26652:data<=-16'd12522;
      26653:data<=-16'd12486;
      26654:data<=-16'd11564;
      26655:data<=-16'd10754;
      26656:data<=-16'd11259;
      26657:data<=-16'd10924;
      26658:data<=-16'd10387;
      26659:data<=-16'd10056;
      26660:data<=-16'd8915;
      26661:data<=-16'd8645;
      26662:data<=-16'd9923;
      26663:data<=-16'd10543;
      26664:data<=-16'd9776;
      26665:data<=-16'd8865;
      26666:data<=-16'd8290;
      26667:data<=-16'd7783;
      26668:data<=-16'd7395;
      26669:data<=-16'd6943;
      26670:data<=-16'd6513;
      26671:data<=-16'd6335;
      26672:data<=-16'd5797;
      26673:data<=-16'd5248;
      26674:data<=-16'd5576;
      26675:data<=-16'd6166;
      26676:data<=-16'd6407;
      26677:data<=-16'd6175;
      26678:data<=-16'd5535;
      26679:data<=-16'd4954;
      26680:data<=-16'd4657;
      26681:data<=-16'd4649;
      26682:data<=-16'd4335;
      26683:data<=-16'd3889;
      26684:data<=-16'd3918;
      26685:data<=-16'd2836;
      26686:data<=-16'd2490;
      26687:data<=-16'd4857;
      26688:data<=-16'd2420;
      26689:data<=16'd5462;
      26690:data<=16'd7846;
      26691:data<=16'd6044;
      26692:data<=16'd6989;
      26693:data<=16'd7310;
      26694:data<=16'd6404;
      26695:data<=16'd7003;
      26696:data<=16'd6871;
      26697:data<=16'd6087;
      26698:data<=16'd6193;
      26699:data<=16'd5559;
      26700:data<=16'd4193;
      26701:data<=16'd3711;
      26702:data<=16'd4071;
      26703:data<=16'd4331;
      26704:data<=16'd4047;
      26705:data<=16'd3826;
      26706:data<=16'd4256;
      26707:data<=16'd4740;
      26708:data<=16'd4440;
      26709:data<=16'd3968;
      26710:data<=16'd4090;
      26711:data<=16'd3852;
      26712:data<=16'd3092;
      26713:data<=16'd2692;
      26714:data<=16'd2273;
      26715:data<=16'd2117;
      26716:data<=16'd2635;
      26717:data<=16'd2693;
      26718:data<=16'd2302;
      26719:data<=16'd2402;
      26720:data<=16'd2810;
      26721:data<=16'd2704;
      26722:data<=16'd2262;
      26723:data<=16'd2711;
      26724:data<=16'd2537;
      26725:data<=16'd419;
      26726:data<=-16'd146;
      26727:data<=16'd1104;
      26728:data<=16'd657;
      26729:data<=-16'd158;
      26730:data<=16'd443;
      26731:data<=16'd1142;
      26732:data<=16'd1339;
      26733:data<=16'd1119;
      26734:data<=16'd954;
      26735:data<=16'd969;
      26736:data<=16'd1732;
      26737:data<=16'd2599;
      26738:data<=-16'd1898;
      26739:data<=-16'd9887;
      26740:data<=-16'd11436;
      26741:data<=-16'd9171;
      26742:data<=-16'd9826;
      26743:data<=-16'd9583;
      26744:data<=-16'd7978;
      26745:data<=-16'd8100;
      26746:data<=-16'd8038;
      26747:data<=-16'd7339;
      26748:data<=-16'd6714;
      26749:data<=-16'd6476;
      26750:data<=-16'd7412;
      26751:data<=-16'd7524;
      26752:data<=-16'd6854;
      26753:data<=-16'd7401;
      26754:data<=-16'd7400;
      26755:data<=-16'd6626;
      26756:data<=-16'd6222;
      26757:data<=-16'd5327;
      26758:data<=-16'd4852;
      26759:data<=-16'd4737;
      26760:data<=-16'd3767;
      26761:data<=-16'd3348;
      26762:data<=-16'd3309;
      26763:data<=-16'd2696;
      26764:data<=-16'd2406;
      26765:data<=-16'd2126;
      26766:data<=-16'd2056;
      26767:data<=-16'd2434;
      26768:data<=-16'd1444;
      26769:data<=-16'd92;
      26770:data<=-16'd500;
      26771:data<=-16'd866;
      26772:data<=-16'd32;
      26773:data<=16'd611;
      26774:data<=16'd1345;
      26775:data<=16'd2892;
      26776:data<=16'd4026;
      26777:data<=16'd4316;
      26778:data<=16'd4390;
      26779:data<=16'd3956;
      26780:data<=16'd3548;
      26781:data<=16'd4155;
      26782:data<=16'd4716;
      26783:data<=16'd4238;
      26784:data<=16'd3896;
      26785:data<=16'd4675;
      26786:data<=16'd4723;
      26787:data<=16'd4029;
      26788:data<=16'd8273;
      26789:data<=16'd16510;
      26790:data<=16'd19038;
      26791:data<=16'd16519;
      26792:data<=16'd16243;
      26793:data<=16'd16525;
      26794:data<=16'd15620;
      26795:data<=16'd15693;
      26796:data<=16'd15579;
      26797:data<=16'd14744;
      26798:data<=16'd14342;
      26799:data<=16'd14302;
      26800:data<=16'd14921;
      26801:data<=16'd15528;
      26802:data<=16'd15220;
      26803:data<=16'd14795;
      26804:data<=16'd14358;
      26805:data<=16'd13800;
      26806:data<=16'd13620;
      26807:data<=16'd13229;
      26808:data<=16'd12471;
      26809:data<=16'd12222;
      26810:data<=16'd11794;
      26811:data<=16'd10615;
      26812:data<=16'd10733;
      26813:data<=16'd12266;
      26814:data<=16'd12414;
      26815:data<=16'd11627;
      26816:data<=16'd11705;
      26817:data<=16'd11461;
      26818:data<=16'd10466;
      26819:data<=16'd9964;
      26820:data<=16'd9947;
      26821:data<=16'd9608;
      26822:data<=16'd9197;
      26823:data<=16'd9354;
      26824:data<=16'd8974;
      26825:data<=16'd8187;
      26826:data<=16'd8889;
      26827:data<=16'd9341;
      26828:data<=16'd8305;
      26829:data<=16'd7912;
      26830:data<=16'd7768;
      26831:data<=16'd7059;
      26832:data<=16'd6181;
      26833:data<=16'd5480;
      26834:data<=16'd6235;
      26835:data<=16'd6216;
      26836:data<=16'd4831;
      26837:data<=16'd6112;
      26838:data<=16'd5432;
      26839:data<=-16'd1096;
      26840:data<=-16'd5012;
      26841:data<=-16'd4335;
      26842:data<=-16'd4322;
      26843:data<=-16'd4156;
      26844:data<=-16'd3545;
      26845:data<=-16'd3700;
      26846:data<=-16'd3730;
      26847:data<=-16'd3789;
      26848:data<=-16'd3407;
      26849:data<=-16'd2914;
      26850:data<=-16'd3072;
      26851:data<=-16'd1591;
      26852:data<=16'd115;
      26853:data<=-16'd993;
      26854:data<=-16'd1612;
      26855:data<=-16'd532;
      26856:data<=-16'd792;
      26857:data<=-16'd1783;
      26858:data<=-16'd2194;
      26859:data<=-16'd1871;
      26860:data<=-16'd682;
      26861:data<=-16'd610;
      26862:data<=-16'd1290;
      26863:data<=16'd20;
      26864:data<=16'd1776;
      26865:data<=16'd1809;
      26866:data<=16'd996;
      26867:data<=16'd425;
      26868:data<=16'd701;
      26869:data<=16'd746;
      26870:data<=-16'd100;
      26871:data<=16'd14;
      26872:data<=16'd293;
      26873:data<=-16'd855;
      26874:data<=-16'd823;
      26875:data<=16'd1515;
      26876:data<=16'd2881;
      26877:data<=16'd1753;
      26878:data<=16'd964;
      26879:data<=16'd1898;
      26880:data<=16'd2026;
      26881:data<=16'd1234;
      26882:data<=16'd1290;
      26883:data<=16'd1340;
      26884:data<=16'd1553;
      26885:data<=16'd2306;
      26886:data<=16'd1528;
      26887:data<=16'd220;
      26888:data<=16'd2987;
      26889:data<=16'd9809;
      26890:data<=16'd13553;
      26891:data<=16'd11776;
      26892:data<=16'd10983;
      26893:data<=16'd11956;
      26894:data<=16'd10933;
      26895:data<=16'd10120;
      26896:data<=16'd9782;
      26897:data<=16'd8595;
      26898:data<=16'd8707;
      26899:data<=16'd9279;
      26900:data<=16'd9843;
      26901:data<=16'd10887;
      26902:data<=16'd9680;
      26903:data<=16'd7862;
      26904:data<=16'd8144;
      26905:data<=16'd8023;
      26906:data<=16'd6953;
      26907:data<=16'd6475;
      26908:data<=16'd6922;
      26909:data<=16'd7215;
      26910:data<=16'd5339;
      26911:data<=16'd3783;
      26912:data<=16'd5580;
      26913:data<=16'd7142;
      26914:data<=16'd5964;
      26915:data<=16'd4848;
      26916:data<=16'd5037;
      26917:data<=16'd4881;
      26918:data<=16'd4256;
      26919:data<=16'd4170;
      26920:data<=16'd4102;
      26921:data<=16'd3748;
      26922:data<=16'd3065;
      26923:data<=16'd1798;
      26924:data<=16'd1319;
      26925:data<=16'd1835;
      26926:data<=16'd2162;
      26927:data<=16'd2149;
      26928:data<=16'd1789;
      26929:data<=16'd2238;
      26930:data<=16'd2875;
      26931:data<=16'd1673;
      26932:data<=16'd623;
      26933:data<=16'd296;
      26934:data<=-16'd115;
      26935:data<=-16'd88;
      26936:data<=-16'd1251;
      26937:data<=-16'd356;
      26938:data<=16'd2193;
      26939:data<=-16'd3290;
      26940:data<=-16'd10329;
      26941:data<=-16'd8715;
      26942:data<=-16'd7567;
      26943:data<=-16'd9726;
      26944:data<=-16'd9477;
      26945:data<=-16'd9248;
      26946:data<=-16'd9359;
      26947:data<=-16'd8939;
      26948:data<=-16'd9724;
      26949:data<=-16'd10169;
      26950:data<=-16'd9015;
      26951:data<=-16'd6915;
      26952:data<=-16'd6159;
      26953:data<=-16'd7160;
      26954:data<=-16'd6842;
      26955:data<=-16'd6833;
      26956:data<=-16'd7758;
      26957:data<=-16'd6704;
      26958:data<=-16'd6208;
      26959:data<=-16'd6554;
      26960:data<=-16'd5809;
      26961:data<=-16'd6205;
      26962:data<=-16'd6775;
      26963:data<=-16'd6602;
      26964:data<=-16'd6871;
      26965:data<=-16'd6478;
      26966:data<=-16'd6090;
      26967:data<=-16'd5788;
      26968:data<=-16'd5468;
      26969:data<=-16'd6263;
      26970:data<=-16'd5491;
      26971:data<=-16'd4149;
      26972:data<=-16'd5422;
      26973:data<=-16'd5874;
      26974:data<=-16'd4889;
      26975:data<=-16'd5172;
      26976:data<=-16'd6522;
      26977:data<=-16'd7815;
      26978:data<=-16'd6965;
      26979:data<=-16'd5694;
      26980:data<=-16'd6520;
      26981:data<=-16'd6630;
      26982:data<=-16'd6006;
      26983:data<=-16'd5723;
      26984:data<=-16'd5401;
      26985:data<=-16'd6244;
      26986:data<=-16'd5647;
      26987:data<=-16'd5239;
      26988:data<=-16'd8284;
      26989:data<=-16'd5529;
      26990:data<=16'd2672;
      26991:data<=16'd3574;
      26992:data<=16'd889;
      26993:data<=16'd1632;
      26994:data<=16'd1961;
      26995:data<=16'd1914;
      26996:data<=16'd2115;
      26997:data<=16'd895;
      26998:data<=16'd883;
      26999:data<=16'd1903;
      27000:data<=16'd802;
      27001:data<=-16'd1162;
      27002:data<=-16'd2190;
      27003:data<=-16'd2582;
      27004:data<=-16'd2009;
      27005:data<=-16'd1116;
      27006:data<=-16'd1653;
      27007:data<=-16'd2347;
      27008:data<=-16'd1350;
      27009:data<=-16'd701;
      27010:data<=-16'd1645;
      27011:data<=-16'd2352;
      27012:data<=-16'd2588;
      27013:data<=-16'd3187;
      27014:data<=-16'd3720;
      27015:data<=-16'd3788;
      27016:data<=-16'd3765;
      27017:data<=-16'd4037;
      27018:data<=-16'd4243;
      27019:data<=-16'd4517;
      27020:data<=-16'd5110;
      27021:data<=-16'd4849;
      27022:data<=-16'd4390;
      27023:data<=-16'd4523;
      27024:data<=-16'd3322;
      27025:data<=-16'd3007;
      27026:data<=-16'd6029;
      27027:data<=-16'd7511;
      27028:data<=-16'd6366;
      27029:data<=-16'd6578;
      27030:data<=-16'd6862;
      27031:data<=-16'd6020;
      27032:data<=-16'd5899;
      27033:data<=-16'd6253;
      27034:data<=-16'd6209;
      27035:data<=-16'd5870;
      27036:data<=-16'd6149;
      27037:data<=-16'd6246;
      27038:data<=-16'd5685;
      27039:data<=-16'd9636;
      27040:data<=-16'd16586;
      27041:data<=-16'd17693;
      27042:data<=-16'd16158;
      27043:data<=-16'd16698;
      27044:data<=-16'd15323;
      27045:data<=-16'd14425;
      27046:data<=-16'd16102;
      27047:data<=-16'd15511;
      27048:data<=-16'd13549;
      27049:data<=-16'd13174;
      27050:data<=-16'd13383;
      27051:data<=-16'd13268;
      27052:data<=-16'd12501;
      27053:data<=-16'd11869;
      27054:data<=-16'd11550;
      27055:data<=-16'd11018;
      27056:data<=-16'd10760;
      27057:data<=-16'd10119;
      27058:data<=-16'd9802;
      27059:data<=-16'd10584;
      27060:data<=-16'd10245;
      27061:data<=-16'd9224;
      27062:data<=-16'd8674;
      27063:data<=-16'd8012;
      27064:data<=-16'd8436;
      27065:data<=-16'd9389;
      27066:data<=-16'd9201;
      27067:data<=-16'd8096;
      27068:data<=-16'd7059;
      27069:data<=-16'd7864;
      27070:data<=-16'd8775;
      27071:data<=-16'd7551;
      27072:data<=-16'd6717;
      27073:data<=-16'd6428;
      27074:data<=-16'd6023;
      27075:data<=-16'd6739;
      27076:data<=-16'd6858;
      27077:data<=-16'd6438;
      27078:data<=-16'd6625;
      27079:data<=-16'd6147;
      27080:data<=-16'd5656;
      27081:data<=-16'd5325;
      27082:data<=-16'd4784;
      27083:data<=-16'd4783;
      27084:data<=-16'd4661;
      27085:data<=-16'd4396;
      27086:data<=-16'd3604;
      27087:data<=-16'd3391;
      27088:data<=-16'd4731;
      27089:data<=-16'd1131;
      27090:data<=16'd6278;
      27091:data<=16'd7753;
      27092:data<=16'd6601;
      27093:data<=16'd7322;
      27094:data<=16'd6628;
      27095:data<=16'd6176;
      27096:data<=16'd6563;
      27097:data<=16'd6478;
      27098:data<=16'd6902;
      27099:data<=16'd6328;
      27100:data<=16'd5946;
      27101:data<=16'd6361;
      27102:data<=16'd4399;
      27103:data<=16'd3250;
      27104:data<=16'd5016;
      27105:data<=16'd5236;
      27106:data<=16'd3723;
      27107:data<=16'd3130;
      27108:data<=16'd3536;
      27109:data<=16'd3789;
      27110:data<=16'd3544;
      27111:data<=16'd4008;
      27112:data<=16'd4726;
      27113:data<=16'd3899;
      27114:data<=16'd2067;
      27115:data<=16'd1588;
      27116:data<=16'd2770;
      27117:data<=16'd2877;
      27118:data<=16'd2127;
      27119:data<=16'd2220;
      27120:data<=16'd1859;
      27121:data<=16'd2432;
      27122:data<=16'd3756;
      27123:data<=16'd2457;
      27124:data<=16'd1695;
      27125:data<=16'd2379;
      27126:data<=16'd916;
      27127:data<=-16'd20;
      27128:data<=16'd561;
      27129:data<=16'd866;
      27130:data<=16'd1733;
      27131:data<=16'd1510;
      27132:data<=16'd748;
      27133:data<=16'd1707;
      27134:data<=16'd2651;
      27135:data<=16'd3215;
      27136:data<=16'd2687;
      27137:data<=16'd1207;
      27138:data<=16'd1389;
      27139:data<=-16'd1128;
      27140:data<=-16'd8158;
      27141:data<=-16'd11623;
      27142:data<=-16'd10084;
      27143:data<=-16'd8940;
      27144:data<=-16'd9169;
      27145:data<=-16'd8895;
      27146:data<=-16'd8040;
      27147:data<=-16'd8050;
      27148:data<=-16'd7515;
      27149:data<=-16'd6167;
      27150:data<=-16'd7424;
      27151:data<=-16'd8542;
      27152:data<=-16'd6551;
      27153:data<=-16'd5912;
      27154:data<=-16'd6463;
      27155:data<=-16'd5169;
      27156:data<=-16'd4432;
      27157:data<=-16'd5178;
      27158:data<=-16'd5127;
      27159:data<=-16'd3544;
      27160:data<=-16'd2670;
      27161:data<=-16'd4102;
      27162:data<=-16'd4686;
      27163:data<=-16'd3081;
      27164:data<=-16'd2149;
      27165:data<=-16'd2344;
      27166:data<=-16'd2578;
      27167:data<=-16'd1751;
      27168:data<=-16'd141;
      27169:data<=-16'd79;
      27170:data<=-16'd632;
      27171:data<=-16'd579;
      27172:data<=-16'd643;
      27173:data<=16'd264;
      27174:data<=16'd822;
      27175:data<=16'd696;
      27176:data<=16'd2685;
      27177:data<=16'd3823;
      27178:data<=16'd2769;
      27179:data<=16'd3494;
      27180:data<=16'd4845;
      27181:data<=16'd4748;
      27182:data<=16'd4205;
      27183:data<=16'd4297;
      27184:data<=16'd5127;
      27185:data<=16'd4475;
      27186:data<=16'd4173;
      27187:data<=16'd5597;
      27188:data<=16'd4773;
      27189:data<=16'd7045;
      27190:data<=16'd15421;
      27191:data<=16'd18883;
      27192:data<=16'd17009;
      27193:data<=16'd16756;
      27194:data<=16'd16841;
      27195:data<=16'd16877;
      27196:data<=16'd15982;
      27197:data<=16'd14199;
      27198:data<=16'd14502;
      27199:data<=16'd14096;
      27200:data<=16'd13650;
      27201:data<=16'd15781;
      27202:data<=16'd15837;
      27203:data<=16'd14771;
      27204:data<=16'd15076;
      27205:data<=16'd14324;
      27206:data<=16'd14474;
      27207:data<=16'd14751;
      27208:data<=16'd12568;
      27209:data<=16'd11508;
      27210:data<=16'd12308;
      27211:data<=16'd12698;
      27212:data<=16'd11976;
      27213:data<=16'd10988;
      27214:data<=16'd11976;
      27215:data<=16'd12872;
      27216:data<=16'd11859;
      27217:data<=16'd11171;
      27218:data<=16'd10470;
      27219:data<=16'd10210;
      27220:data<=16'd10572;
      27221:data<=16'd9574;
      27222:data<=16'd9420;
      27223:data<=16'd9849;
      27224:data<=16'd8354;
      27225:data<=16'd7896;
      27226:data<=16'd9165;
      27227:data<=16'd9814;
      27228:data<=16'd9844;
      27229:data<=16'd9646;
      27230:data<=16'd8992;
      27231:data<=16'd7292;
      27232:data<=16'd6557;
      27233:data<=16'd7230;
      27234:data<=16'd6062;
      27235:data<=16'd5988;
      27236:data<=16'd7426;
      27237:data<=16'd5988;
      27238:data<=16'd6604;
      27239:data<=16'd7752;
      27240:data<=16'd1707;
      27241:data<=-16'd3516;
      27242:data<=-16'd3207;
      27243:data<=-16'd3322;
      27244:data<=-16'd2617;
      27245:data<=-16'd1568;
      27246:data<=-16'd2877;
      27247:data<=-16'd3380;
      27248:data<=-16'd3328;
      27249:data<=-16'd3550;
      27250:data<=-16'd1924;
      27251:data<=-16'd466;
      27252:data<=-16'd476;
      27253:data<=16'd431;
      27254:data<=16'd1779;
      27255:data<=16'd870;
      27256:data<=-16'd989;
      27257:data<=-16'd341;
      27258:data<=16'd775;
      27259:data<=-16'd588;
      27260:data<=-16'd1242;
      27261:data<=16'd226;
      27262:data<=16'd848;
      27263:data<=16'd664;
      27264:data<=16'd1325;
      27265:data<=16'd2452;
      27266:data<=16'd3084;
      27267:data<=16'd2708;
      27268:data<=16'd1853;
      27269:data<=16'd1486;
      27270:data<=16'd1794;
      27271:data<=16'd2488;
      27272:data<=16'd2648;
      27273:data<=16'd1915;
      27274:data<=16'd1700;
      27275:data<=16'd1985;
      27276:data<=16'd1962;
      27277:data<=16'd3149;
      27278:data<=16'd4434;
      27279:data<=16'd3115;
      27280:data<=16'd2364;
      27281:data<=16'd4114;
      27282:data<=16'd4313;
      27283:data<=16'd2766;
      27284:data<=16'd2634;
      27285:data<=16'd3066;
      27286:data<=16'd2872;
      27287:data<=16'd3178;
      27288:data<=16'd3550;
      27289:data<=16'd4522;
      27290:data<=16'd9163;
      27291:data<=16'd14266;
      27292:data<=16'd14427;
      27293:data<=16'd13256;
      27294:data<=16'd13136;
      27295:data<=16'd11684;
      27296:data<=16'd10963;
      27297:data<=16'd10759;
      27298:data<=16'd9727;
      27299:data<=16'd10219;
      27300:data<=16'd9568;
      27301:data<=16'd7780;
      27302:data<=16'd9315;
      27303:data<=16'd10085;
      27304:data<=16'd8100;
      27305:data<=16'd7460;
      27306:data<=16'd7492;
      27307:data<=16'd7732;
      27308:data<=16'd7874;
      27309:data<=16'd6249;
      27310:data<=16'd5424;
      27311:data<=16'd6310;
      27312:data<=16'd6807;
      27313:data<=16'd6707;
      27314:data<=16'd6226;
      27315:data<=16'd6226;
      27316:data<=16'd6219;
      27317:data<=16'd5096;
      27318:data<=16'd4864;
      27319:data<=16'd5453;
      27320:data<=16'd4813;
      27321:data<=16'd4024;
      27322:data<=16'd4141;
      27323:data<=16'd3976;
      27324:data<=16'd2969;
      27325:data<=16'd2978;
      27326:data<=16'd4117;
      27327:data<=16'd3474;
      27328:data<=16'd2315;
      27329:data<=16'd3149;
      27330:data<=16'd3806;
      27331:data<=16'd3365;
      27332:data<=16'd2704;
      27333:data<=16'd1538;
      27334:data<=16'd843;
      27335:data<=16'd1773;
      27336:data<=16'd2736;
      27337:data<=16'd1374;
      27338:data<=16'd447;
      27339:data<=16'd2206;
      27340:data<=-16'd476;
      27341:data<=-16'd8401;
      27342:data<=-16'd11094;
      27343:data<=-16'd8895;
      27344:data<=-16'd9097;
      27345:data<=-16'd9855;
      27346:data<=-16'd8645;
      27347:data<=-16'd7523;
      27348:data<=-16'd7222;
      27349:data<=-16'd7366;
      27350:data<=-16'd8213;
      27351:data<=-16'd8434;
      27352:data<=-16'd6792;
      27353:data<=-16'd6191;
      27354:data<=-16'd7121;
      27355:data<=-16'd6150;
      27356:data<=-16'd5488;
      27357:data<=-16'd6893;
      27358:data<=-16'd6980;
      27359:data<=-16'd6275;
      27360:data<=-16'd6125;
      27361:data<=-16'd5976;
      27362:data<=-16'd6664;
      27363:data<=-16'd7086;
      27364:data<=-16'd6572;
      27365:data<=-16'd6199;
      27366:data<=-16'd5783;
      27367:data<=-16'd5981;
      27368:data<=-16'd6537;
      27369:data<=-16'd6529;
      27370:data<=-16'd6557;
      27371:data<=-16'd5996;
      27372:data<=-16'd5771;
      27373:data<=-16'd6968;
      27374:data<=-16'd6822;
      27375:data<=-16'd5598;
      27376:data<=-16'd5890;
      27377:data<=-16'd6811;
      27378:data<=-16'd7574;
      27379:data<=-16'd8052;
      27380:data<=-16'd7247;
      27381:data<=-16'd6147;
      27382:data<=-16'd6643;
      27383:data<=-16'd7503;
      27384:data<=-16'd6939;
      27385:data<=-16'd6610;
      27386:data<=-16'd7131;
      27387:data<=-16'd6478;
      27388:data<=-16'd5510;
      27389:data<=-16'd5238;
      27390:data<=-16'd1885;
      27391:data<=16'd4780;
      27392:data<=16'd6696;
      27393:data<=16'd4255;
      27394:data<=16'd5882;
      27395:data<=16'd5859;
      27396:data<=16'd1598;
      27397:data<=16'd2056;
      27398:data<=16'd805;
      27399:data<=16'd1577;
      27400:data<=16'd15262;
      27401:data<=16'd14360;
      27402:data<=-16'd5832;
      27403:data<=-16'd7918;
      27404:data<=16'd241;
      27405:data<=-16'd4478;
      27406:data<=-16'd8235;
      27407:data<=-16'd5903;
      27408:data<=-16'd3228;
      27409:data<=16'd663;
      27410:data<=16'd1836;
      27411:data<=-16'd1404;
      27412:data<=-16'd6196;
      27413:data<=-16'd7122;
      27414:data<=-16'd3682;
      27415:data<=-16'd3553;
      27416:data<=-16'd3991;
      27417:data<=-16'd2538;
      27418:data<=-16'd3956;
      27419:data<=-16'd2397;
      27420:data<=16'd2420;
      27421:data<=16'd628;
      27422:data<=-16'd6799;
      27423:data<=-16'd10442;
      27424:data<=-16'd8278;
      27425:data<=-16'd10663;
      27426:data<=-16'd15327;
      27427:data<=-16'd10373;
      27428:data<=-16'd5808;
      27429:data<=-16'd6837;
      27430:data<=-16'd6493;
      27431:data<=-16'd8674;
      27432:data<=-16'd8530;
      27433:data<=-16'd6090;
      27434:data<=-16'd10951;
      27435:data<=-16'd11402;
      27436:data<=-16'd3701;
      27437:data<=-16'd825;
      27438:data<=-16'd3786;
      27439:data<=-16'd7485;
      27440:data<=-16'd8088;
      27441:data<=-16'd12613;
      27442:data<=-16'd21995;
      27443:data<=-16'd20439;
      27444:data<=-16'd17164;
      27445:data<=-16'd23631;
      27446:data<=-16'd25335;
      27447:data<=-16'd21029;
      27448:data<=-16'd17371;
      27449:data<=-16'd16926;
      27450:data<=-16'd19446;
      27451:data<=-16'd17030;
      27452:data<=-16'd15221;
      27453:data<=-16'd14969;
      27454:data<=-16'd12330;
      27455:data<=-16'd18724;
      27456:data<=-16'd21842;
      27457:data<=-16'd15242;
      27458:data<=-16'd17658;
      27459:data<=-16'd16832;
      27460:data<=-16'd9511;
      27461:data<=-16'd10489;
      27462:data<=-16'd10560;
      27463:data<=-16'd12417;
      27464:data<=-16'd17209;
      27465:data<=-16'd16205;
      27466:data<=-16'd16877;
      27467:data<=-16'd12907;
      27468:data<=-16'd5600;
      27469:data<=-16'd6721;
      27470:data<=-16'd5662;
      27471:data<=-16'd7043;
      27472:data<=-16'd12122;
      27473:data<=-16'd7448;
      27474:data<=-16'd6015;
      27475:data<=-16'd9871;
      27476:data<=-16'd9896;
      27477:data<=-16'd10666;
      27478:data<=-16'd9338;
      27479:data<=-16'd9198;
      27480:data<=-16'd8343;
      27481:data<=-16'd3251;
      27482:data<=-16'd7776;
      27483:data<=-16'd12346;
      27484:data<=-16'd11368;
      27485:data<=-16'd13970;
      27486:data<=-16'd5545;
      27487:data<=-16'd414;
      27488:data<=-16'd13902;
      27489:data<=-16'd14648;
      27490:data<=-16'd3177;
      27491:data<=-16'd234;
      27492:data<=-16'd1394;
      27493:data<=-16'd2270;
      27494:data<=16'd2840;
      27495:data<=16'd8199;
      27496:data<=16'd7181;
      27497:data<=16'd9570;
      27498:data<=16'd8889;
      27499:data<=16'd5227;
      27500:data<=16'd8739;
      27501:data<=16'd8392;
      27502:data<=16'd7272;
      27503:data<=16'd11465;
      27504:data<=16'd7517;
      27505:data<=16'd4084;
      27506:data<=16'd13048;
      27507:data<=16'd16311;
      27508:data<=16'd6307;
      27509:data<=16'd3290;
      27510:data<=16'd10383;
      27511:data<=16'd10426;
      27512:data<=16'd6896;
      27513:data<=16'd5755;
      27514:data<=16'd5333;
      27515:data<=16'd11913;
      27516:data<=16'd13661;
      27517:data<=16'd9535;
      27518:data<=16'd14883;
      27519:data<=16'd12276;
      27520:data<=16'd7973;
      27521:data<=16'd19729;
      27522:data<=16'd18066;
      27523:data<=16'd9727;
      27524:data<=16'd16007;
      27525:data<=16'd14536;
      27526:data<=16'd12507;
      27527:data<=16'd17045;
      27528:data<=16'd11737;
      27529:data<=16'd12188;
      27530:data<=16'd16562;
      27531:data<=16'd8053;
      27532:data<=16'd6492;
      27533:data<=16'd15074;
      27534:data<=16'd13626;
      27535:data<=16'd9680;
      27536:data<=16'd15462;
      27537:data<=16'd15618;
      27538:data<=16'd7689;
      27539:data<=16'd11379;
      27540:data<=16'd12367;
      27541:data<=16'd914;
      27542:data<=16'd3701;
      27543:data<=16'd8771;
      27544:data<=16'd993;
      27545:data<=16'd2294;
      27546:data<=16'd6454;
      27547:data<=16'd6024;
      27548:data<=16'd6978;
      27549:data<=16'd425;
      27550:data<=-16'd1483;
      27551:data<=16'd3497;
      27552:data<=16'd281;
      27553:data<=16'd3724;
      27554:data<=16'd9809;
      27555:data<=16'd4188;
      27556:data<=16'd3385;
      27557:data<=16'd5034;
      27558:data<=16'd2185;
      27559:data<=16'd7210;
      27560:data<=16'd13007;
      27561:data<=16'd8558;
      27562:data<=16'd1947;
      27563:data<=16'd1137;
      27564:data<=16'd1289;
      27565:data<=-16'd667;
      27566:data<=16'd2995;
      27567:data<=16'd6467;
      27568:data<=16'd5494;
      27569:data<=16'd9157;
      27570:data<=16'd6777;
      27571:data<=16'd3723;
      27572:data<=16'd16316;
      27573:data<=16'd14915;
      27574:data<=-16'd3037;
      27575:data<=-16'd1192;
      27576:data<=16'd8921;
      27577:data<=16'd9614;
      27578:data<=16'd8214;
      27579:data<=16'd4425;
      27580:data<=16'd5676;
      27581:data<=16'd10295;
      27582:data<=16'd6561;
      27583:data<=16'd4484;
      27584:data<=16'd6501;
      27585:data<=16'd7441;
      27586:data<=16'd10320;
      27587:data<=16'd6754;
      27588:data<=16'd1122;
      27589:data<=16'd5856;
      27590:data<=16'd9882;
      27591:data<=16'd12266;
      27592:data<=16'd18442;
      27593:data<=16'd16584;
      27594:data<=16'd11778;
      27595:data<=16'd14205;
      27596:data<=16'd13224;
      27597:data<=16'd8514;
      27598:data<=16'd8432;
      27599:data<=16'd9053;
      27600:data<=16'd10079;
      27601:data<=16'd13982;
      27602:data<=16'd12598;
      27603:data<=16'd5330;
      27604:data<=16'd5159;
      27605:data<=16'd10498;
      27606:data<=16'd8493;
      27607:data<=16'd2792;
      27608:data<=16'd1830;
      27609:data<=16'd2849;
      27610:data<=16'd1271;
      27611:data<=-16'd1186;
      27612:data<=16'd3409;
      27613:data<=16'd8922;
      27614:data<=16'd728;
      27615:data<=-16'd8749;
      27616:data<=-16'd7662;
      27617:data<=-16'd5736;
      27618:data<=-16'd1739;
      27619:data<=16'd1636;
      27620:data<=-16'd3762;
      27621:data<=-16'd8346;
      27622:data<=-16'd10910;
      27623:data<=-16'd10272;
      27624:data<=-16'd1695;
      27625:data<=-16'd3345;
      27626:data<=-16'd10847;
      27627:data<=-16'd5313;
      27628:data<=-16'd3707;
      27629:data<=-16'd7051;
      27630:data<=-16'd3862;
      27631:data<=-16'd8194;
      27632:data<=-16'd10466;
      27633:data<=-16'd1785;
      27634:data<=-16'd5545;
      27635:data<=-16'd13300;
      27636:data<=-16'd7166;
      27637:data<=-16'd5761;
      27638:data<=-16'd11344;
      27639:data<=-16'd7112;
      27640:data<=-16'd4367;
      27641:data<=-16'd16146;
      27642:data<=-16'd24251;
      27643:data<=-16'd18730;
      27644:data<=-16'd17415;
      27645:data<=-16'd20967;
      27646:data<=-16'd17690;
      27647:data<=-16'd16308;
      27648:data<=-16'd17206;
      27649:data<=-16'd14302;
      27650:data<=-16'd16525;
      27651:data<=-16'd17511;
      27652:data<=-16'd10507;
      27653:data<=-16'd9841;
      27654:data<=-16'd14953;
      27655:data<=-16'd18536;
      27656:data<=-16'd19654;
      27657:data<=-16'd12619;
      27658:data<=-16'd9424;
      27659:data<=-16'd17643;
      27660:data<=-16'd19212;
      27661:data<=-16'd15471;
      27662:data<=-16'd13966;
      27663:data<=-16'd7953;
      27664:data<=-16'd5603;
      27665:data<=-16'd8094;
      27666:data<=-16'd6401;
      27667:data<=-16'd7808;
      27668:data<=-16'd10539;
      27669:data<=-16'd10188;
      27670:data<=-16'd12774;
      27671:data<=-16'd11223;
      27672:data<=-16'd7641;
      27673:data<=-16'd11952;
      27674:data<=-16'd11684;
      27675:data<=-16'd5471;
      27676:data<=-16'd7524;
      27677:data<=-16'd11646;
      27678:data<=-16'd8149;
      27679:data<=-16'd5271;
      27680:data<=-16'd9638;
      27681:data<=-16'd9066;
      27682:data<=-16'd1184;
      27683:data<=-16'd6504;
      27684:data<=-16'd16732;
      27685:data<=-16'd10002;
      27686:data<=-16'd5153;
      27687:data<=-16'd11471;
      27688:data<=-16'd10963;
      27689:data<=-16'd6912;
      27690:data<=-16'd2775;
      27691:data<=16'd6431;
      27692:data<=16'd11468;
      27693:data<=16'd9028;
      27694:data<=16'd5054;
      27695:data<=16'd4913;
      27696:data<=16'd8031;
      27697:data<=16'd3433;
      27698:data<=-16'd428;
      27699:data<=16'd7905;
      27700:data<=16'd8479;
      27701:data<=16'd1271;
      27702:data<=16'd5136;
      27703:data<=16'd7787;
      27704:data<=16'd5871;
      27705:data<=16'd11771;
      27706:data<=16'd13670;
      27707:data<=16'd7024;
      27708:data<=16'd5444;
      27709:data<=16'd10319;
      27710:data<=16'd14155;
      27711:data<=16'd11332;
      27712:data<=16'd8247;
      27713:data<=16'd11752;
      27714:data<=16'd10029;
      27715:data<=16'd4269;
      27716:data<=16'd8426;
      27717:data<=16'd12598;
      27718:data<=16'd9233;
      27719:data<=16'd8702;
      27720:data<=16'd12063;
      27721:data<=16'd13523;
      27722:data<=16'd11852;
      27723:data<=16'd11611;
      27724:data<=16'd12254;
      27725:data<=16'd5036;
      27726:data<=16'd610;
      27727:data<=16'd9374;
      27728:data<=16'd12510;
      27729:data<=16'd5645;
      27730:data<=16'd3116;
      27731:data<=16'd4796;
      27732:data<=16'd9197;
      27733:data<=16'd13547;
      27734:data<=16'd12947;
      27735:data<=16'd11426;
      27736:data<=16'd9694;
      27737:data<=16'd10458;
      27738:data<=16'd13679;
      27739:data<=16'd8727;
      27740:data<=16'd2601;
      27741:data<=16'd2951;
      27742:data<=16'd2722;
      27743:data<=16'd5280;
      27744:data<=16'd4804;
      27745:data<=-16'd3838;
      27746:data<=-16'd4079;
      27747:data<=-16'd235;
      27748:data<=-16'd2514;
      27749:data<=-16'd3256;
      27750:data<=-16'd2954;
      27751:data<=16'd1862;
      27752:data<=16'd5315;
      27753:data<=-16'd2557;
      27754:data<=16'd1715;
      27755:data<=16'd12102;
      27756:data<=16'd2517;
      27757:data<=-16'd2373;
      27758:data<=16'd2344;
      27759:data<=16'd412;
      27760:data<=16'd5589;
      27761:data<=16'd6764;
      27762:data<=-16'd572;
      27763:data<=16'd5630;
      27764:data<=16'd8607;
      27765:data<=16'd4081;
      27766:data<=16'd9444;
      27767:data<=16'd8718;
      27768:data<=16'd2504;
      27769:data<=16'd4041;
      27770:data<=16'd5254;
      27771:data<=16'd7383;
      27772:data<=16'd7131;
      27773:data<=16'd2968;
      27774:data<=16'd7924;
      27775:data<=16'd11185;
      27776:data<=16'd4999;
      27777:data<=16'd4899;
      27778:data<=16'd10052;
      27779:data<=16'd10627;
      27780:data<=16'd7203;
      27781:data<=16'd4951;
      27782:data<=16'd4302;
      27783:data<=16'd5116;
      27784:data<=16'd12839;
      27785:data<=16'd13204;
      27786:data<=16'd328;
      27787:data<=16'd2450;
      27788:data<=16'd11520;
      27789:data<=16'd7457;
      27790:data<=16'd11016;
      27791:data<=16'd18665;
      27792:data<=16'd17142;
      27793:data<=16'd16903;
      27794:data<=16'd13759;
      27795:data<=16'd12063;
      27796:data<=16'd13747;
      27797:data<=16'd6921;
      27798:data<=16'd9078;
      27799:data<=16'd14201;
      27800:data<=16'd2493;
      27801:data<=16'd3160;
      27802:data<=16'd13444;
      27803:data<=16'd5791;
      27804:data<=-16'd1266;
      27805:data<=-16'd795;
      27806:data<=16'd277;
      27807:data<=16'd4878;
      27808:data<=16'd4006;
      27809:data<=16'd2883;
      27810:data<=16'd2032;
      27811:data<=-16'd8079;
      27812:data<=-16'd6020;
      27813:data<=16'd5322;
      27814:data<=-16'd766;
      27815:data<=-16'd8589;
      27816:data<=-16'd5800;
      27817:data<=-16'd3877;
      27818:data<=-16'd3758;
      27819:data<=-16'd5846;
      27820:data<=-16'd6050;
      27821:data<=-16'd1222;
      27822:data<=-16'd1485;
      27823:data<=-16'd6795;
      27824:data<=-16'd8217;
      27825:data<=-16'd3717;
      27826:data<=-16'd2858;
      27827:data<=-16'd13327;
      27828:data<=-16'd17194;
      27829:data<=-16'd7785;
      27830:data<=-16'd6351;
      27831:data<=-16'd11420;
      27832:data<=-16'd10395;
      27833:data<=-16'd7533;
      27834:data<=-16'd6943;
      27835:data<=-16'd8792;
      27836:data<=-16'd7327;
      27837:data<=-16'd5683;
      27838:data<=-16'd11323;
      27839:data<=-16'd8771;
      27840:data<=-16'd6288;
      27841:data<=-16'd22522;
      27842:data<=-16'd26442;
      27843:data<=-16'd17108;
      27844:data<=-16'd23713;
      27845:data<=-16'd22732;
      27846:data<=-16'd14590;
      27847:data<=-16'd24115;
      27848:data<=-16'd22664;
      27849:data<=-16'd8772;
      27850:data<=-16'd11746;
      27851:data<=-16'd16636;
      27852:data<=-16'd17185;
      27853:data<=-16'd19781;
      27854:data<=-16'd12349;
      27855:data<=-16'd8075;
      27856:data<=-16'd16380;
      27857:data<=-16'd16125;
      27858:data<=-16'd10828;
      27859:data<=-16'd13449;
      27860:data<=-16'd13209;
      27861:data<=-16'd8943;
      27862:data<=-16'd11518;
      27863:data<=-16'd17541;
      27864:data<=-16'd16709;
      27865:data<=-16'd11314;
      27866:data<=-16'd11855;
      27867:data<=-16'd15350;
      27868:data<=-16'd12991;
      27869:data<=-16'd10753;
      27870:data<=-16'd11382;
      27871:data<=-16'd7761;
      27872:data<=-16'd5504;
      27873:data<=-16'd9985;
      27874:data<=-16'd12437;
      27875:data<=-16'd11377;
      27876:data<=-16'd11520;
      27877:data<=-16'd10800;
      27878:data<=-16'd8467;
      27879:data<=-16'd6868;
      27880:data<=-16'd8402;
      27881:data<=-16'd10463;
      27882:data<=-16'd6037;
      27883:data<=-16'd2687;
      27884:data<=-16'd8370;
      27885:data<=-16'd10316;
      27886:data<=-16'd6211;
      27887:data<=-16'd6214;
      27888:data<=-16'd5488;
      27889:data<=-16'd1760;
      27890:data<=16'd544;
      27891:data<=16'd3968;
      27892:data<=16'd6032;
      27893:data<=16'd4447;
      27894:data<=16'd3007;
      27895:data<=16'd949;
      27896:data<=16'd657;
      27897:data<=16'd4081;
      27898:data<=16'd4281;
      27899:data<=16'd2752;
      27900:data<=16'd5909;
      27901:data<=16'd8426;
      27902:data<=16'd7224;
      27903:data<=16'd7514;
      27904:data<=16'd8012;
      27905:data<=16'd6434;
      27906:data<=16'd6044;
      27907:data<=16'd4883;
      27908:data<=16'd2614;
      27909:data<=16'd5028;
      27910:data<=16'd9364;
      27911:data<=16'd10998;
      27912:data<=16'd9668;
      27913:data<=16'd4816;
      27914:data<=16'd3990;
      27915:data<=16'd9254;
      27916:data<=16'd10636;
      27917:data<=16'd10269;
      27918:data<=16'd11600;
      27919:data<=16'd7708;
      27920:data<=16'd1518;
      27921:data<=16'd2396;
      27922:data<=16'd7903;
      27923:data<=16'd6601;
      27924:data<=16'd3095;
      27925:data<=16'd9729;
      27926:data<=16'd12190;
      27927:data<=16'd6698;
      27928:data<=16'd10724;
      27929:data<=16'd12195;
      27930:data<=16'd8223;
      27931:data<=16'd13053;
      27932:data<=16'd10950;
      27933:data<=16'd6205;
      27934:data<=16'd12577;
      27935:data<=16'd10013;
      27936:data<=16'd5274;
      27937:data<=16'd10273;
      27938:data<=16'd7444;
      27939:data<=16'd3433;
      27940:data<=16'd4008;
      27941:data<=-16'd722;
      27942:data<=-16'd984;
      27943:data<=16'd2614;
      27944:data<=16'd886;
      27945:data<=16'd1460;
      27946:data<=16'd5538;
      27947:data<=16'd5958;
      27948:data<=16'd3121;
      27949:data<=16'd2772;
      27950:data<=16'd2675;
      27951:data<=16'd262;
      27952:data<=16'd4034;
      27953:data<=16'd5524;
      27954:data<=-16'd1209;
      27955:data<=16'd2801;
      27956:data<=16'd8839;
      27957:data<=16'd5033;
      27958:data<=16'd7326;
      27959:data<=16'd8525;
      27960:data<=16'd3547;
      27961:data<=16'd3917;
      27962:data<=16'd2799;
      27963:data<=16'd4197;
      27964:data<=16'd9430;
      27965:data<=16'd4238;
      27966:data<=16'd1679;
      27967:data<=16'd5968;
      27968:data<=16'd1591;
      27969:data<=16'd1204;
      27970:data<=16'd9767;
      27971:data<=16'd7824;
      27972:data<=16'd44;
      27973:data<=16'd1824;
      27974:data<=16'd5934;
      27975:data<=16'd6203;
      27976:data<=16'd6382;
      27977:data<=16'd3251;
      27978:data<=16'd3412;
      27979:data<=16'd10198;
      27980:data<=16'd6454;
      27981:data<=16'd1700;
      27982:data<=16'd7732;
      27983:data<=16'd6214;
      27984:data<=16'd5494;
      27985:data<=16'd9964;
      27986:data<=16'd3065;
      27987:data<=16'd3163;
      27988:data<=16'd9239;
      27989:data<=16'd4372;
      27990:data<=16'd10205;
      27991:data<=16'd19146;
      27992:data<=16'd13443;
      27993:data<=16'd13855;
      27994:data<=16'd17602;
      27995:data<=16'd12712;
      27996:data<=16'd10076;
      27997:data<=16'd12587;
      27998:data<=16'd13769;
      27999:data<=16'd8617;
      28000:data<=16'd6893;
      28001:data<=16'd11608;
      28002:data<=16'd6730;
      28003:data<=16'd3397;
      28004:data<=16'd7201;
      28005:data<=16'd1930;
      28006:data<=16'd3280;
      28007:data<=16'd10895;
      28008:data<=16'd4146;
      28009:data<=16'd282;
      28010:data<=16'd5430;
      28011:data<=16'd5802;
      28012:data<=16'd3356;
      28013:data<=-16'd669;
      28014:data<=-16'd479;
      28015:data<=16'd3348;
      28016:data<=-16'd453;
      28017:data<=-16'd3336;
      28018:data<=16'd23;
      28019:data<=-16'd993;
      28020:data<=-16'd6833;
      28021:data<=-16'd8067;
      28022:data<=-16'd2343;
      28023:data<=-16'd2593;
      28024:data<=-16'd6909;
      28025:data<=-16'd1519;
      28026:data<=-16'd1249;
      28027:data<=-16'd9221;
      28028:data<=-16'd7078;
      28029:data<=-16'd3920;
      28030:data<=-16'd7649;
      28031:data<=-16'd10806;
      28032:data<=-16'd10492;
      28033:data<=-16'd4040;
      28034:data<=-16'd2510;
      28035:data<=-16'd8432;
      28036:data<=-16'd6959;
      28037:data<=-16'd5177;
      28038:data<=-16'd6253;
      28039:data<=-16'd4185;
      28040:data<=-16'd11558;
      28041:data<=-16'd21077;
      28042:data<=-16'd16280;
      28043:data<=-16'd12692;
      28044:data<=-16'd19441;
      28045:data<=-16'd19895;
      28046:data<=-16'd11647;
      28047:data<=-16'd14637;
      28048:data<=-16'd25860;
      28049:data<=-16'd22588;
      28050:data<=-16'd14383;
      28051:data<=-16'd15606;
      28052:data<=-16'd17017;
      28053:data<=-16'd16305;
      28054:data<=-16'd11365;
      28055:data<=-16'd8161;
      28056:data<=-16'd17763;
      28057:data<=-16'd20310;
      28058:data<=-16'd13253;
      28059:data<=-16'd17276;
      28060:data<=-16'd20659;
      28061:data<=-16'd16732;
      28062:data<=-16'd14378;
      28063:data<=-16'd12563;
      28064:data<=-16'd13706;
      28065:data<=-16'd9791;
      28066:data<=-16'd3424;
      28067:data<=-16'd11135;
      28068:data<=-16'd14753;
      28069:data<=-16'd7517;
      28070:data<=-16'd7156;
      28071:data<=-16'd5213;
      28072:data<=-16'd3195;
      28073:data<=-16'd8331;
      28074:data<=-16'd6103;
      28075:data<=-16'd3368;
      28076:data<=-16'd9426;
      28077:data<=-16'd10477;
      28078:data<=-16'd7401;
      28079:data<=-16'd9706;
      28080:data<=-16'd12237;
      28081:data<=-16'd10334;
      28082:data<=-16'd9051;
      28083:data<=-16'd7932;
      28084:data<=-16'd5156;
      28085:data<=-16'd7806;
      28086:data<=-16'd8752;
      28087:data<=-16'd4502;
      28088:data<=-16'd9016;
      28089:data<=-16'd8995;
      28090:data<=16'd790;
      28091:data<=-16'd519;
      28092:data<=-16'd249;
      28093:data<=16'd7824;
      28094:data<=16'd7893;
      28095:data<=16'd6799;
      28096:data<=16'd4077;
      28097:data<=16'd1851;
      28098:data<=16'd9527;
      28099:data<=16'd11107;
      28100:data<=16'd5821;
      28101:data<=16'd3300;
      28102:data<=16'd2784;
      28103:data<=16'd10543;
      28104:data<=16'd12028;
      28105:data<=16'd3776;
      28106:data<=16'd6677;
      28107:data<=16'd9793;
      28108:data<=16'd9109;
      28109:data<=16'd11627;
      28110:data<=16'd7641;
      28111:data<=16'd8564;
      28112:data<=16'd12486;
      28113:data<=16'd6355;
      28114:data<=16'd7782;
      28115:data<=16'd13688;
      28116:data<=16'd13396;
      28117:data<=16'd13453;
      28118:data<=16'd9198;
      28119:data<=16'd8987;
      28120:data<=16'd13835;
      28121:data<=16'd9582;
      28122:data<=16'd10328;
      28123:data<=16'd15967;
      28124:data<=16'd10319;
      28125:data<=16'd8338;
      28126:data<=16'd17124;
      28127:data<=16'd17823;
      28128:data<=16'd7727;
      28129:data<=16'd6795;
      28130:data<=16'd14789;
      28131:data<=16'd13355;
      28132:data<=16'd10402;
      28133:data<=16'd11054;
      28134:data<=16'd8334;
      28135:data<=16'd11141;
      28136:data<=16'd13021;
      28137:data<=16'd11483;
      28138:data<=16'd14416;
      28139:data<=16'd7953;
      28140:data<=16'd3019;
      28141:data<=16'd5415;
      28142:data<=-16'd4839;
      28143:data<=-16'd5764;
      28144:data<=16'd4552;
      28145:data<=16'd913;
      28146:data<=-16'd1165;
      28147:data<=-16'd999;
      28148:data<=-16'd1036;
      28149:data<=16'd6364;
      28150:data<=16'd2375;
      28151:data<=-16'd714;
      28152:data<=16'd7908;
      28153:data<=16'd6860;
      28154:data<=16'd7154;
      28155:data<=16'd8407;
      28156:data<=16'd1246;
      28157:data<=16'd2229;
      28158:data<=16'd2863;
      28159:data<=16'd2631;
      28160:data<=16'd9638;
      28161:data<=16'd5855;
      28162:data<=16'd752;
      28163:data<=16'd4009;
      28164:data<=16'd2000;
      28165:data<=16'd1412;
      28166:data<=16'd5768;
      28167:data<=16'd10354;
      28168:data<=16'd10508;
      28169:data<=16'd2541;
      28170:data<=16'd1595;
      28171:data<=16'd5160;
      28172:data<=16'd1022;
      28173:data<=16'd604;
      28174:data<=16'd3673;
      28175:data<=16'd5140;
      28176:data<=16'd4777;
      28177:data<=16'd578;
      28178:data<=16'd3479;
      28179:data<=16'd8059;
      28180:data<=16'd6910;
      28181:data<=16'd11042;
      28182:data<=16'd10281;
      28183:data<=16'd4458;
      28184:data<=16'd7879;
      28185:data<=16'd9702;
      28186:data<=16'd9160;
      28187:data<=16'd9796;
      28188:data<=16'd5820;
      28189:data<=16'd7269;
      28190:data<=16'd13135;
      28191:data<=16'd14354;
      28192:data<=16'd13714;
      28193:data<=16'd10919;
      28194:data<=16'd11477;
      28195:data<=16'd17020;
      28196:data<=16'd18086;
      28197:data<=16'd12928;
      28198:data<=16'd5770;
      28199:data<=16'd7494;
      28200:data<=16'd12968;
      28201:data<=16'd3521;
      28202:data<=-16'd2598;
      28203:data<=16'd8331;
      28204:data<=16'd8981;
      28205:data<=-16'd3459;
      28206:data<=-16'd4889;
      28207:data<=16'd3935;
      28208:data<=16'd6237;
      28209:data<=16'd1237;
      28210:data<=-16'd872;
      28211:data<=-16'd1823;
      28212:data<=-16'd3964;
      28213:data<=-16'd1177;
      28214:data<=16'd2558;
      28215:data<=-16'd516;
      28216:data<=-16'd5618;
      28217:data<=-16'd3116;
      28218:data<=16'd1131;
      28219:data<=-16'd3566;
      28220:data<=-16'd6560;
      28221:data<=-16'd6149;
      28222:data<=-16'd10252;
      28223:data<=-16'd5676;
      28224:data<=-16'd1580;
      28225:data<=-16'd10843;
      28226:data<=-16'd10084;
      28227:data<=-16'd5658;
      28228:data<=-16'd11799;
      28229:data<=-16'd9944;
      28230:data<=-16'd8261;
      28231:data<=-16'd11600;
      28232:data<=-16'd4018;
      28233:data<=-16'd3049;
      28234:data<=-16'd11241;
      28235:data<=-16'd6830;
      28236:data<=-16'd3526;
      28237:data<=-16'd10545;
      28238:data<=-16'd10646;
      28239:data<=-16'd6704;
      28240:data<=-16'd11130;
      28241:data<=-16'd17896;
      28242:data<=-16'd18977;
      28243:data<=-16'd16286;
      28244:data<=-16'd14857;
      28245:data<=-16'd17594;
      28246:data<=-16'd18164;
      28247:data<=-16'd14942;
      28248:data<=-16'd19038;
      28249:data<=-16'd20594;
      28250:data<=-16'd10572;
      28251:data<=-16'd11699;
      28252:data<=-16'd18668;
      28253:data<=-16'd11468;
      28254:data<=-16'd10824;
      28255:data<=-16'd19949;
      28256:data<=-16'd17823;
      28257:data<=-16'd12301;
      28258:data<=-16'd11526;
      28259:data<=-16'd11315;
      28260:data<=-16'd13960;
      28261:data<=-16'd17875;
      28262:data<=-16'd19256;
      28263:data<=-16'd16055;
      28264:data<=-16'd9629;
      28265:data<=-16'd8442;
      28266:data<=-16'd12489;
      28267:data<=-16'd12037;
      28268:data<=-16'd8918;
      28269:data<=-16'd12145;
      28270:data<=-16'd13253;
      28271:data<=-16'd5551;
      28272:data<=-16'd5873;
      28273:data<=-16'd11586;
      28274:data<=-16'd6821;
      28275:data<=-16'd6211;
      28276:data<=-16'd12383;
      28277:data<=-16'd10716;
      28278:data<=-16'd8651;
      28279:data<=-16'd7482;
      28280:data<=-16'd6598;
      28281:data<=-16'd13876;
      28282:data<=-16'd16366;
      28283:data<=-16'd11121;
      28284:data<=-16'd12364;
      28285:data<=-16'd14213;
      28286:data<=-16'd10937;
      28287:data<=-16'd9159;
      28288:data<=-16'd10076;
      28289:data<=-16'd7923;
      28290:data<=-16'd1042;
      28291:data<=16'd164;
      28292:data<=-16'd1245;
      28293:data<=16'd5896;
      28294:data<=16'd7586;
      28295:data<=16'd1403;
      28296:data<=16'd3858;
      28297:data<=16'd7567;
      28298:data<=16'd5846;
      28299:data<=16'd8049;
      28300:data<=16'd13013;
      28301:data<=16'd15026;
      28302:data<=16'd14010;
      28303:data<=16'd13179;
      28304:data<=16'd14225;
      28305:data<=16'd14813;
      28306:data<=16'd15179;
      28307:data<=16'd14694;
      28308:data<=16'd12784;
      28309:data<=16'd12824;
      28310:data<=16'd13858;
      28311:data<=16'd14358;
      28312:data<=16'd14343;
      28313:data<=16'd13382;
      28314:data<=16'd13347;
      28315:data<=16'd12646;
      28316:data<=16'd12737;
      28317:data<=16'd15359;
      28318:data<=16'd13441;
      28319:data<=16'd11529;
      28320:data<=16'd14298;
      28321:data<=16'd12292;
      28322:data<=16'd10704;
      28323:data<=16'd14504;
      28324:data<=16'd14022;
      28325:data<=16'd11862;
      28326:data<=16'd12216;
      28327:data<=16'd11872;
      28328:data<=16'd11389;
      28329:data<=16'd10608;
      28330:data<=16'd11822;
      28331:data<=16'd13806;
      28332:data<=16'd11876;
      28333:data<=16'd11127;
      28334:data<=16'd11781;
      28335:data<=16'd11101;
      28336:data<=16'd12451;
      28337:data<=16'd11556;
      28338:data<=16'd9630;
      28339:data<=16'd11640;
      28340:data<=16'd8672;
      28341:data<=16'd1498;
      28342:data<=16'd408;
      28343:data<=16'd2091;
      28344:data<=16'd1066;
      28345:data<=-16'd388;
      28346:data<=16'd378;
      28347:data<=16'd355;
      28348:data<=-16'd1221;
      28349:data<=16'd834;
      28350:data<=16'd2231;
      28351:data<=16'd461;
      28352:data<=16'd2270;
      28353:data<=16'd2479;
      28354:data<=16'd52;
      28355:data<=16'd2628;
      28356:data<=16'd3632;
      28357:data<=16'd1571;
      28358:data<=16'd2093;
      28359:data<=16'd1756;
      28360:data<=16'd2214;
      28361:data<=16'd4140;
      28362:data<=16'd3694;
      28363:data<=16'd3456;
      28364:data<=16'd2379;
      28365:data<=16'd1310;
      28366:data<=16'd3457;
      28367:data<=16'd3770;
      28368:data<=16'd3823;
      28369:data<=16'd5465;
      28370:data<=16'd3507;
      28371:data<=16'd2218;
      28372:data<=16'd3394;
      28373:data<=16'd3266;
      28374:data<=16'd3912;
      28375:data<=16'd3826;
      28376:data<=16'd3544;
      28377:data<=16'd4725;
      28378:data<=16'd2805;
      28379:data<=16'd2258;
      28380:data<=16'd5147;
      28381:data<=16'd4438;
      28382:data<=16'd3565;
      28383:data<=16'd3527;
      28384:data<=16'd1574;
      28385:data<=16'd2943;
      28386:data<=16'd4356;
      28387:data<=16'd3325;
      28388:data<=16'd4610;
      28389:data<=16'd3823;
      28390:data<=16'd4363;
      28391:data<=16'd11705;
      28392:data<=16'd13509;
      28393:data<=16'd9853;
      28394:data<=16'd11298;
      28395:data<=16'd11831;
      28396:data<=16'd9512;
      28397:data<=16'd9547;
      28398:data<=16'd8025;
      28399:data<=16'd5324;
      28400:data<=16'd5521;
      28401:data<=16'd5360;
      28402:data<=16'd3906;
      28403:data<=16'd3701;
      28404:data<=16'd3200;
      28405:data<=16'd1407;
      28406:data<=16'd760;
      28407:data<=16'd1031;
      28408:data<=16'd490;
      28409:data<=16'd553;
      28410:data<=16'd769;
      28411:data<=-16'd789;
      28412:data<=-16'd2237;
      28413:data<=-16'd2596;
      28414:data<=-16'd2314;
      28415:data<=-16'd1574;
      28416:data<=-16'd2349;
      28417:data<=-16'd4000;
      28418:data<=-16'd5016;
      28419:data<=-16'd5630;
      28420:data<=-16'd4760;
      28421:data<=-16'd4596;
      28422:data<=-16'd5932;
      28423:data<=-16'd5465;
      28424:data<=-16'd5938;
      28425:data<=-16'd7611;
      28426:data<=-16'd6815;
      28427:data<=-16'd6636;
      28428:data<=-16'd7318;
      28429:data<=-16'd7520;
      28430:data<=-16'd8704;
      28431:data<=-16'd8302;
      28432:data<=-16'd8052;
      28433:data<=-16'd8872;
      28434:data<=-16'd6670;
      28435:data<=-16'd6495;
      28436:data<=-16'd9227;
      28437:data<=-16'd9344;
      28438:data<=-16'd9589;
      28439:data<=-16'd9162;
      28440:data<=-16'd9321;
      28441:data<=-16'd15697;
      28442:data<=-16'd20213;
      28443:data<=-16'd19029;
      28444:data<=-16'd19009;
      28445:data<=-16'd19359;
      28446:data<=-16'd18398;
      28447:data<=-16'd16689;
      28448:data<=-16'd15926;
      28449:data<=-16'd18292;
      28450:data<=-16'd18709;
      28451:data<=-16'd16475;
      28452:data<=-16'd15461;
      28453:data<=-16'd14099;
      28454:data<=-16'd14794;
      28455:data<=-16'd16254;
      28456:data<=-16'd13737;
      28457:data<=-16'd13145;
      28458:data<=-16'd14368;
      28459:data<=-16'd12536;
      28460:data<=-16'd12698;
      28461:data<=-16'd14835;
      28462:data<=-16'd14731;
      28463:data<=-16'd13979;
      28464:data<=-16'd13251;
      28465:data<=-16'd12484;
      28466:data<=-16'd12079;
      28467:data<=-16'd12049;
      28468:data<=-16'd12099;
      28469:data<=-16'd11162;
      28470:data<=-16'd10831;
      28471:data<=-16'd10994;
      28472:data<=-16'd9621;
      28473:data<=-16'd9209;
      28474:data<=-16'd9934;
      28475:data<=-16'd9871;
      28476:data<=-16'd10044;
      28477:data<=-16'd9690;
      28478:data<=-16'd8819;
      28479:data<=-16'd8827;
      28480:data<=-16'd9101;
      28481:data<=-16'd9216;
      28482:data<=-16'd8900;
      28483:data<=-16'd9160;
      28484:data<=-16'd9500;
      28485:data<=-16'd8533;
      28486:data<=-16'd9201;
      28487:data<=-16'd9130;
      28488:data<=-16'd6579;
      28489:data<=-16'd8012;
      28490:data<=-16'd7028;
      28491:data<=16'd1709;
      28492:data<=16'd5212;
      28493:data<=16'd3421;
      28494:data<=16'd4936;
      28495:data<=16'd5344;
      28496:data<=16'd4344;
      28497:data<=16'd4943;
      28498:data<=16'd5178;
      28499:data<=16'd5850;
      28500:data<=16'd6056;
      28501:data<=16'd5260;
      28502:data<=16'd6023;
      28503:data<=16'd6581;
      28504:data<=16'd6526;
      28505:data<=16'd7253;
      28506:data<=16'd7677;
      28507:data<=16'd9053;
      28508:data<=16'd10345;
      28509:data<=16'd9095;
      28510:data<=16'd8281;
      28511:data<=16'd8960;
      28512:data<=16'd9744;
      28513:data<=16'd10329;
      28514:data<=16'd9109;
      28515:data<=16'd7827;
      28516:data<=16'd8613;
      28517:data<=16'd9294;
      28518:data<=16'd9694;
      28519:data<=16'd9644;
      28520:data<=16'd8859;
      28521:data<=16'd9009;
      28522:data<=16'd8252;
      28523:data<=16'd8062;
      28524:data<=16'd11056;
      28525:data<=16'd11157;
      28526:data<=16'd9241;
      28527:data<=16'd10743;
      28528:data<=16'd10531;
      28529:data<=16'd8925;
      28530:data<=16'd10379;
      28531:data<=16'd10777;
      28532:data<=16'd10229;
      28533:data<=16'd10739;
      28534:data<=16'd9955;
      28535:data<=16'd9944;
      28536:data<=16'd11514;
      28537:data<=16'd11347;
      28538:data<=16'd9850;
      28539:data<=16'd9885;
      28540:data<=16'd10376;
      28541:data<=16'd6253;
      28542:data<=16'd773;
      28543:data<=16'd1371;
      28544:data<=16'd2843;
      28545:data<=16'd1560;
      28546:data<=16'd2018;
      28547:data<=16'd2367;
      28548:data<=16'd2551;
      28549:data<=16'd4366;
      28550:data<=16'd3929;
      28551:data<=16'd3027;
      28552:data<=16'd3914;
      28553:data<=16'd3448;
      28554:data<=16'd3751;
      28555:data<=16'd5871;
      28556:data<=16'd5843;
      28557:data<=16'd4687;
      28558:data<=16'd4924;
      28559:data<=16'd4884;
      28560:data<=16'd4516;
      28561:data<=16'd5651;
      28562:data<=16'd6131;
      28563:data<=16'd5236;
      28564:data<=16'd5820;
      28565:data<=16'd5557;
      28566:data<=16'd3932;
      28567:data<=16'd5221;
      28568:data<=16'd6719;
      28569:data<=16'd6135;
      28570:data<=16'd6405;
      28571:data<=16'd7033;
      28572:data<=16'd6965;
      28573:data<=16'd6446;
      28574:data<=16'd6927;
      28575:data<=16'd8614;
      28576:data<=16'd7814;
      28577:data<=16'd6784;
      28578:data<=16'd7241;
      28579:data<=16'd5674;
      28580:data<=16'd6332;
      28581:data<=16'd8294;
      28582:data<=16'd6460;
      28583:data<=16'd6620;
      28584:data<=16'd6874;
      28585:data<=16'd4478;
      28586:data<=16'd6096;
      28587:data<=16'd7271;
      28588:data<=16'd6352;
      28589:data<=16'd7483;
      28590:data<=16'd6276;
      28591:data<=16'd8689;
      28592:data<=16'd16258;
      28593:data<=16'd15872;
      28594:data<=16'd12833;
      28595:data<=16'd14302;
      28596:data<=16'd13236;
      28597:data<=16'd11603;
      28598:data<=16'd10850;
      28599:data<=16'd8064;
      28600:data<=16'd7465;
      28601:data<=16'd8247;
      28602:data<=16'd7482;
      28603:data<=16'd7432;
      28604:data<=16'd6542;
      28605:data<=16'd3997;
      28606:data<=16'd3209;
      28607:data<=16'd3717;
      28608:data<=16'd2892;
      28609:data<=16'd1777;
      28610:data<=16'd1973;
      28611:data<=16'd1456;
      28612:data<=-16'd499;
      28613:data<=-16'd1492;
      28614:data<=-16'd1563;
      28615:data<=-16'd1533;
      28616:data<=-16'd1240;
      28617:data<=-16'd1902;
      28618:data<=-16'd3388;
      28619:data<=-16'd4188;
      28620:data<=-16'd4660;
      28621:data<=-16'd5045;
      28622:data<=-16'd4246;
      28623:data<=-16'd3770;
      28624:data<=-16'd5896;
      28625:data<=-16'd7194;
      28626:data<=-16'd5850;
      28627:data<=-16'd5853;
      28628:data<=-16'd6103;
      28629:data<=-16'd5836;
      28630:data<=-16'd7971;
      28631:data<=-16'd8117;
      28632:data<=-16'd6454;
      28633:data<=-16'd8373;
      28634:data<=-16'd8326;
      28635:data<=-16'd6166;
      28636:data<=-16'd7862;
      28637:data<=-16'd8149;
      28638:data<=-16'd7139;
      28639:data<=-16'd8613;
      28640:data<=-16'd7410;
      28641:data<=-16'd8479;
      28642:data<=-16'd16681;
      28643:data<=-16'd20553;
      28644:data<=-16'd18383;
      28645:data<=-16'd18228;
      28646:data<=-16'd18161;
      28647:data<=-16'd16689;
      28648:data<=-16'd16477;
      28649:data<=-16'd16847;
      28650:data<=-16'd16857;
      28651:data<=-16'd16216;
      28652:data<=-16'd15787;
      28653:data<=-16'd16043;
      28654:data<=-16'd14756;
      28655:data<=-16'd13861;
      28656:data<=-16'd15628;
      28657:data<=-16'd15593;
      28658:data<=-16'd13315;
      28659:data<=-16'd12557;
      28660:data<=-16'd12302;
      28661:data<=-16'd12408;
      28662:data<=-16'd13497;
      28663:data<=-16'd12910;
      28664:data<=-16'd11526;
      28665:data<=-16'd11793;
      28666:data<=-16'd12066;
      28667:data<=-16'd11796;
      28668:data<=-16'd11873;
      28669:data<=-16'd11436;
      28670:data<=-16'd10722;
      28671:data<=-16'd10455;
      28672:data<=-16'd9926;
      28673:data<=-16'd9712;
      28674:data<=-16'd10572;
      28675:data<=-16'd10928;
      28676:data<=-16'd10248;
      28677:data<=-16'd9829;
      28678:data<=-16'd9506;
      28679:data<=-16'd9175;
      28680:data<=-16'd10055;
      28681:data<=-16'd11030;
      28682:data<=-16'd10078;
      28683:data<=-16'd9212;
      28684:data<=-16'd9711;
      28685:data<=-16'd8481;
      28686:data<=-16'd7072;
      28687:data<=-16'd8746;
      28688:data<=-16'd8813;
      28689:data<=-16'd7301;
      28690:data<=-16'd8645;
      28691:data<=-16'd5709;
      28692:data<=16'd2575;
      28693:data<=16'd5080;
      28694:data<=16'd3733;
      28695:data<=16'd4388;
      28696:data<=16'd3902;
      28697:data<=16'd3874;
      28698:data<=16'd5231;
      28699:data<=16'd4895;
      28700:data<=16'd5369;
      28701:data<=16'd6807;
      28702:data<=16'd6620;
      28703:data<=16'd6159;
      28704:data<=16'd5909;
      28705:data<=16'd6686;
      28706:data<=16'd8581;
      28707:data<=16'd8752;
      28708:data<=16'd8263;
      28709:data<=16'd8473;
      28710:data<=16'd8003;
      28711:data<=16'd8257;
      28712:data<=16'd9080;
      28713:data<=16'd8707;
      28714:data<=16'd8966;
      28715:data<=16'd9676;
      28716:data<=16'd8980;
      28717:data<=16'd9001;
      28718:data<=16'd10378;
      28719:data<=16'd10627;
      28720:data<=16'd10322;
      28721:data<=16'd10564;
      28722:data<=16'd10035;
      28723:data<=16'd9768;
      28724:data<=16'd11156;
      28725:data<=16'd11849;
      28726:data<=16'd11194;
      28727:data<=16'd11306;
      28728:data<=16'd11593;
      28729:data<=16'd10777;
      28730:data<=16'd10950;
      28731:data<=16'd12572;
      28732:data<=16'd12146;
      28733:data<=16'd10842;
      28734:data<=16'd11888;
      28735:data<=16'd11590;
      28736:data<=16'd10355;
      28737:data<=16'd12451;
      28738:data<=16'd12595;
      28739:data<=16'd10621;
      28740:data<=16'd12199;
      28741:data<=16'd9899;
      28742:data<=16'd2130;
      28743:data<=16'd249;
      28744:data<=16'd2626;
      28745:data<=16'd2408;
      28746:data<=16'd2024;
      28747:data<=16'd2135;
      28748:data<=16'd1833;
      28749:data<=16'd2913;
      28750:data<=16'd4400;
      28751:data<=16'd4329;
      28752:data<=16'd3885;
      28753:data<=16'd4002;
      28754:data<=16'd3735;
      28755:data<=16'd4258;
      28756:data<=16'd5771;
      28757:data<=16'd5338;
      28758:data<=16'd4723;
      28759:data<=16'd5592;
      28760:data<=16'd4860;
      28761:data<=16'd4554;
      28762:data<=16'd6061;
      28763:data<=16'd5927;
      28764:data<=16'd5600;
      28765:data<=16'd5700;
      28766:data<=16'd4763;
      28767:data<=16'd5137;
      28768:data<=16'd6031;
      28769:data<=16'd5944;
      28770:data<=16'd6234;
      28771:data<=16'd6146;
      28772:data<=16'd5764;
      28773:data<=16'd5412;
      28774:data<=16'd5303;
      28775:data<=16'd6633;
      28776:data<=16'd6678;
      28777:data<=16'd5424;
      28778:data<=16'd5659;
      28779:data<=16'd4939;
      28780:data<=16'd4549;
      28781:data<=16'd6308;
      28782:data<=16'd6024;
      28783:data<=16'd5159;
      28784:data<=16'd5817;
      28785:data<=16'd5536;
      28786:data<=16'd5306;
      28787:data<=16'd5624;
      28788:data<=16'd6131;
      28789:data<=16'd6040;
      28790:data<=16'd3814;
      28791:data<=16'd5535;
      28792:data<=16'd12416;
      28793:data<=16'd14795;
      28794:data<=16'd13317;
      28795:data<=16'd13344;
      28796:data<=16'd12331;
      28797:data<=16'd10789;
      28798:data<=16'd10707;
      28799:data<=16'd9955;
      28800:data<=16'd8272;
      28801:data<=16'd6990;
      28802:data<=16'd6299;
      28803:data<=16'd6053;
      28804:data<=16'd5856;
      28805:data<=16'd4570;
      28806:data<=16'd2460;
      28807:data<=16'd1729;
      28808:data<=16'd1527;
      28809:data<=16'd723;
      28810:data<=16'd792;
      28811:data<=16'd108;
      28812:data<=-16'd1536;
      28813:data<=-16'd1850;
      28814:data<=-16'd2531;
      28815:data<=-16'd3110;
      28816:data<=-16'd2394;
      28817:data<=-16'd2934;
      28818:data<=-16'd4021;
      28819:data<=-16'd4852;
      28820:data<=-16'd5927;
      28821:data<=-16'd5868;
      28822:data<=-16'd5718;
      28823:data<=-16'd5582;
      28824:data<=-16'd5670;
      28825:data<=-16'd7793;
      28826:data<=-16'd8246;
      28827:data<=-16'd7172;
      28828:data<=-16'd8204;
      28829:data<=-16'd7817;
      28830:data<=-16'd7332;
      28831:data<=-16'd9288;
      28832:data<=-16'd9112;
      28833:data<=-16'd8672;
      28834:data<=-16'd9903;
      28835:data<=-16'd9653;
      28836:data<=-16'd9620;
      28837:data<=-16'd9949;
      28838:data<=-16'd10119;
      28839:data<=-16'd11092;
      28840:data<=-16'd10232;
      28841:data<=-16'd11036;
      28842:data<=-16'd16724;
      28843:data<=-16'd20583;
      28844:data<=-16'd21315;
      28845:data<=-16'd21799;
      28846:data<=-16'd21291;
      28847:data<=-16'd20622;
      28848:data<=-16'd19667;
      28849:data<=-16'd19162;
      28850:data<=-16'd20202;
      28851:data<=-16'd19605;
      28852:data<=-16'd18642;
      28853:data<=-16'd18989;
      28854:data<=-16'd17379;
      28855:data<=-16'd16553;
      28856:data<=-16'd18130;
      28857:data<=-16'd17566;
      28858:data<=-16'd16166;
      28859:data<=-16'd16028;
      28860:data<=-16'd15188;
      28861:data<=-16'd14363;
      28862:data<=-16'd14624;
      28863:data<=-16'd15033;
      28864:data<=-16'd14616;
      28865:data<=-16'd13541;
      28866:data<=-16'd13076;
      28867:data<=-16'd12868;
      28868:data<=-16'd12844;
      28869:data<=-16'd13399;
      28870:data<=-16'd12692;
      28871:data<=-16'd11709;
      28872:data<=-16'd12051;
      28873:data<=-16'd11348;
      28874:data<=-16'd10586;
      28875:data<=-16'd11535;
      28876:data<=-16'd11461;
      28877:data<=-16'd10480;
      28878:data<=-16'd10108;
      28879:data<=-16'd9307;
      28880:data<=-16'd9197;
      28881:data<=-16'd10240;
      28882:data<=-16'd10120;
      28883:data<=-16'd9430;
      28884:data<=-16'd9424;
      28885:data<=-16'd8513;
      28886:data<=-16'd7553;
      28887:data<=-16'd8763;
      28888:data<=-16'd9418;
      28889:data<=-16'd8058;
      28890:data<=-16'd7870;
      28891:data<=-16'd6628;
      28892:data<=-16'd766;
      28893:data<=16'd4319;
      28894:data<=16'd4755;
      28895:data<=16'd4435;
      28896:data<=16'd5125;
      28897:data<=16'd5195;
      28898:data<=16'd4854;
      28899:data<=16'd5548;
      28900:data<=16'd6754;
      28901:data<=16'd6863;
      28902:data<=16'd6968;
      28903:data<=16'd7586;
      28904:data<=16'd6946;
      28905:data<=16'd6721;
      28906:data<=16'd8269;
      28907:data<=16'd8906;
      28908:data<=16'd8687;
      28909:data<=16'd8957;
      28910:data<=16'd8560;
      28911:data<=16'd8223;
      28912:data<=16'd9344;
      28913:data<=16'd10440;
      28914:data<=16'd10357;
      28915:data<=16'd10135;
      28916:data<=16'd10158;
      28917:data<=16'd9885;
      28918:data<=16'd10355;
      28919:data<=16'd11402;
      28920:data<=16'd11132;
      28921:data<=16'd11065;
      28922:data<=16'd11811;
      28923:data<=16'd10966;
      28924:data<=16'd10555;
      28925:data<=16'd11987;
      28926:data<=16'd12383;
      28927:data<=16'd12320;
      28928:data<=16'd12464;
      28929:data<=16'd11511;
      28930:data<=16'd11320;
      28931:data<=16'd12357;
      28932:data<=16'd12885;
      28933:data<=16'd12965;
      28934:data<=16'd12639;
      28935:data<=16'd12020;
      28936:data<=16'd11473;
      28937:data<=16'd11955;
      28938:data<=16'd13585;
      28939:data<=16'd13229;
      28940:data<=16'd12349;
      28941:data<=16'd12645;
      28942:data<=16'd7849;
      28943:data<=16'd1691;
      28944:data<=16'd2795;
      28945:data<=16'd4288;
      28946:data<=16'd3040;
      28947:data<=16'd3753;
      28948:data<=16'd3328;
      28949:data<=16'd2823;
      28950:data<=16'd4925;
      28951:data<=16'd5365;
      28952:data<=16'd5119;
      28953:data<=16'd5439;
      28954:data<=16'd4592;
      28955:data<=16'd5134;
      28956:data<=16'd6402;
      28957:data<=16'd6549;
      28958:data<=16'd6928;
      28959:data<=16'd6552;
      28960:data<=16'd5802;
      28961:data<=16'd5938;
      28962:data<=16'd6569;
      28963:data<=16'd7668;
      28964:data<=16'd7365;
      28965:data<=16'd6504;
      28966:data<=16'd6840;
      28967:data<=16'd6041;
      28968:data<=16'd6194;
      28969:data<=16'd8437;
      28970:data<=16'd8470;
      28971:data<=16'd7686;
      28972:data<=16'd7550;
      28973:data<=16'd6557;
      28974:data<=16'd6918;
      28975:data<=16'd8196;
      28976:data<=16'd8082;
      28977:data<=16'd7876;
      28978:data<=16'd8138;
      28979:data<=16'd7609;
      28980:data<=16'd6587;
      28981:data<=16'd7353;
      28982:data<=16'd8517;
      28983:data<=16'd7327;
      28984:data<=16'd6839;
      28985:data<=16'd7197;
      28986:data<=16'd6209;
      28987:data<=16'd6422;
      28988:data<=16'd6927;
      28989:data<=16'd7127;
      28990:data<=16'd7618;
      28991:data<=16'd5935;
      28992:data<=16'd8025;
      28993:data<=16'd15032;
      28994:data<=16'd16547;
      28995:data<=16'd14877;
      28996:data<=16'd14701;
      28997:data<=16'd13245;
      28998:data<=16'd13367;
      28999:data<=16'd13423;
      29000:data<=16'd10560;
      29001:data<=16'd9306;
      29002:data<=16'd8493;
      29003:data<=16'd7125;
      29004:data<=16'd7577;
      29005:data<=16'd7197;
      29006:data<=16'd5395;
      29007:data<=16'd3859;
      29008:data<=16'd3115;
      29009:data<=16'd3110;
      29010:data<=16'd2337;
      29011:data<=16'd2049;
      29012:data<=16'd1522;
      29013:data<=-16'd974;
      29014:data<=-16'd1240;
      29015:data<=-16'd566;
      29016:data<=-16'd1864;
      29017:data<=-16'd1515;
      29018:data<=-16'd1568;
      29019:data<=-16'd3802;
      29020:data<=-16'd4733;
      29021:data<=-16'd5253;
      29022:data<=-16'd5501;
      29023:data<=-16'd4737;
      29024:data<=-16'd4908;
      29025:data<=-16'd5911;
      29026:data<=-16'd6956;
      29027:data<=-16'd7227;
      29028:data<=-16'd7115;
      29029:data<=-16'd7327;
      29030:data<=-16'd6366;
      29031:data<=-16'd6683;
      29032:data<=-16'd8470;
      29033:data<=-16'd7788;
      29034:data<=-16'd7843;
      29035:data<=-16'd8660;
      29036:data<=-16'd7219;
      29037:data<=-16'd7779;
      29038:data<=-16'd9462;
      29039:data<=-16'd10006;
      29040:data<=-16'd10684;
      29041:data<=-16'd8980;
      29042:data<=-16'd10528;
      29043:data<=-16'd18750;
      29044:data<=-16'd22457;
      29045:data<=-16'd21171;
      29046:data<=-16'd21488;
      29047:data<=-16'd20648;
      29048:data<=-16'd19311;
      29049:data<=-16'd19666;
      29050:data<=-16'd19957;
      29051:data<=-16'd20296;
      29052:data<=-16'd19776;
      29053:data<=-16'd18527;
      29054:data<=-16'd17932;
      29055:data<=-16'd16892;
      29056:data<=-16'd16798;
      29057:data<=-16'd17917;
      29058:data<=-16'd17333;
      29059:data<=-16'd16477;
      29060:data<=-16'd16249;
      29061:data<=-16'd14854;
      29062:data<=-16'd14431;
      29063:data<=-16'd15743;
      29064:data<=-16'd15752;
      29065:data<=-16'd14966;
      29066:data<=-16'd14580;
      29067:data<=-16'd13302;
      29068:data<=-16'd12780;
      29069:data<=-16'd13964;
      29070:data<=-16'd13711;
      29071:data<=-16'd12627;
      29072:data<=-16'd12660;
      29073:data<=-16'd11876;
      29074:data<=-16'd11072;
      29075:data<=-16'd11973;
      29076:data<=-16'd12404;
      29077:data<=-16'd11740;
      29078:data<=-16'd11271;
      29079:data<=-16'd11022;
      29080:data<=-16'd10602;
      29081:data<=-16'd10426;
      29082:data<=-16'd11550;
      29083:data<=-16'd12276;
      29084:data<=-16'd11035;
      29085:data<=-16'd10275;
      29086:data<=-16'd9814;
      29087:data<=-16'd9206;
      29088:data<=-16'd10551;
      29089:data<=-16'd10354;
      29090:data<=-16'd8308;
      29091:data<=-16'd9072;
      29092:data<=-16'd6510;
      29093:data<=16'd1624;
      29094:data<=16'd4681;
      29095:data<=16'd3334;
      29096:data<=16'd4325;
      29097:data<=16'd4548;
      29098:data<=16'd3603;
      29099:data<=16'd4120;
      29100:data<=16'd4983;
      29101:data<=16'd6384;
      29102:data<=16'd7150;
      29103:data<=16'd6341;
      29104:data<=16'd6208;
      29105:data<=16'd5809;
      29106:data<=16'd5703;
      29107:data<=16'd7806;
      29108:data<=16'd8398;
      29109:data<=16'd7582;
      29110:data<=16'd8090;
      29111:data<=16'd7400;
      29112:data<=16'd6898;
      29113:data<=16'd8637;
      29114:data<=16'd9380;
      29115:data<=16'd9550;
      29116:data<=16'd9730;
      29117:data<=16'd8405;
      29118:data<=16'd8411;
      29119:data<=16'd10140;
      29120:data<=16'd10449;
      29121:data<=16'd9993;
      29122:data<=16'd9847;
      29123:data<=16'd9394;
      29124:data<=16'd8893;
      29125:data<=16'd9348;
      29126:data<=16'd10598;
      29127:data<=16'd10728;
      29128:data<=16'd10290;
      29129:data<=16'd10628;
      29130:data<=16'd9803;
      29131:data<=16'd9056;
      29132:data<=16'd10766;
      29133:data<=16'd11611;
      29134:data<=16'd10837;
      29135:data<=16'd10774;
      29136:data<=16'd9900;
      29137:data<=16'd9351;
      29138:data<=16'd11229;
      29139:data<=16'd11600;
      29140:data<=16'd10627;
      29141:data<=16'd11326;
      29142:data<=16'd8191;
      29143:data<=16'd1165;
      29144:data<=-16'd49;
      29145:data<=16'd2364;
      29146:data<=16'd1080;
      29147:data<=16'd326;
      29148:data<=16'd1691;
      29149:data<=16'd1259;
      29150:data<=16'd1475;
      29151:data<=16'd3251;
      29152:data<=16'd3480;
      29153:data<=16'd3325;
      29154:data<=16'd3482;
      29155:data<=16'd2719;
      29156:data<=16'd3058;
      29157:data<=16'd4874;
      29158:data<=16'd5275;
      29159:data<=16'd4596;
      29160:data<=16'd4432;
      29161:data<=16'd4140;
      29162:data<=16'd4632;
      29163:data<=16'd6419;
      29164:data<=16'd6717;
      29165:data<=16'd5636;
      29166:data<=16'd5671;
      29167:data<=16'd5829;
      29168:data<=16'd5218;
      29169:data<=16'd5597;
      29170:data<=16'd6645;
      29171:data<=16'd6431;
      29172:data<=16'd6156;
      29173:data<=16'd6628;
      29174:data<=16'd5665;
      29175:data<=16'd5382;
      29176:data<=16'd7514;
      29177:data<=16'd7238;
      29178:data<=16'd5776;
      29179:data<=16'd6549;
      29180:data<=16'd5877;
      29181:data<=16'd5909;
      29182:data<=16'd8452;
      29183:data<=16'd7708;
      29184:data<=16'd6161;
      29185:data<=16'd6830;
      29186:data<=16'd6338;
      29187:data<=16'd6516;
      29188:data<=16'd7427;
      29189:data<=16'd7221;
      29190:data<=16'd7362;
      29191:data<=16'd6596;
      29192:data<=16'd8226;
      29193:data<=16'd14413;
      29194:data<=16'd16824;
      29195:data<=16'd15355;
      29196:data<=16'd15465;
      29197:data<=16'd14521;
      29198:data<=16'd13019;
      29199:data<=16'd13124;
      29200:data<=16'd12135;
      29201:data<=16'd10205;
      29202:data<=16'd8933;
      29203:data<=16'd7720;
      29204:data<=16'd6846;
      29205:data<=16'd6940;
      29206:data<=16'd6407;
      29207:data<=16'd4156;
      29208:data<=16'd2705;
      29209:data<=16'd2523;
      29210:data<=16'd1989;
      29211:data<=16'd2259;
      29212:data<=16'd1800;
      29213:data<=-16'd670;
      29214:data<=-16'd1604;
      29215:data<=-16'd1347;
      29216:data<=-16'd1804;
      29217:data<=-16'd1768;
      29218:data<=-16'd1730;
      29219:data<=-16'd2676;
      29220:data<=-16'd4352;
      29221:data<=-16'd5215;
      29222:data<=-16'd4939;
      29223:data<=-16'd5571;
      29224:data<=-16'd5389;
      29225:data<=-16'd4763;
      29226:data<=-16'd6963;
      29227:data<=-16'd7826;
      29228:data<=-16'd6683;
      29229:data<=-16'd7144;
      29230:data<=-16'd6496;
      29231:data<=-16'd6608;
      29232:data<=-16'd9277;
      29233:data<=-16'd9580;
      29234:data<=-16'd9095;
      29235:data<=-16'd9350;
      29236:data<=-16'd8431;
      29237:data<=-16'd8815;
      29238:data<=-16'd9824;
      29239:data<=-16'd10043;
      29240:data<=-16'd10430;
      29241:data<=-16'd9659;
      29242:data<=-16'd10828;
      29243:data<=-16'd16101;
      29244:data<=-16'd20269;
      29245:data<=-16'd21514;
      29246:data<=-16'd21409;
      29247:data<=-16'd20387;
      29248:data<=-16'd18894;
      29249:data<=-16'd17355;
      29250:data<=-16'd17684;
      29251:data<=-16'd19297;
      29252:data<=-16'd19027;
      29253:data<=-16'd17720;
      29254:data<=-16'd16645;
      29255:data<=-16'd15631;
      29256:data<=-16'd15669;
      29257:data<=-16'd16278;
      29258:data<=-16'd16321;
      29259:data<=-16'd15675;
      29260:data<=-16'd14780;
      29261:data<=-16'd14272;
      29262:data<=-16'd13920;
      29263:data<=-16'd14172;
      29264:data<=-16'd14781;
      29265:data<=-16'd14327;
      29266:data<=-16'd13928;
      29267:data<=-16'd13405;
      29268:data<=-16'd11776;
      29269:data<=-16'd12096;
      29270:data<=-16'd13819;
      29271:data<=-16'd13106;
      29272:data<=-16'd11900;
      29273:data<=-16'd11975;
      29274:data<=-16'd11271;
      29275:data<=-16'd10830;
      29276:data<=-16'd12038;
      29277:data<=-16'd12369;
      29278:data<=-16'd11421;
      29279:data<=-16'd11276;
      29280:data<=-16'd11012;
      29281:data<=-16'd10194;
      29282:data<=-16'd10504;
      29283:data<=-16'd10843;
      29284:data<=-16'd10191;
      29285:data<=-16'd9899;
      29286:data<=-16'd9611;
      29287:data<=-16'd8877;
      29288:data<=-16'd9124;
      29289:data<=-16'd9906;
      29290:data<=-16'd9527;
      29291:data<=-16'd9101;
      29292:data<=-16'd8652;
      29293:data<=-16'd4605;
      29294:data<=16'd873;
      29295:data<=16'd2002;
      29296:data<=16'd1497;
      29297:data<=16'd2502;
      29298:data<=16'd2224;
      29299:data<=16'd1741;
      29300:data<=16'd3234;
      29301:data<=16'd4592;
      29302:data<=16'd4925;
      29303:data<=16'd5004;
      29304:data<=16'd4928;
      29305:data<=16'd4708;
      29306:data<=16'd4980;
      29307:data<=16'd6285;
      29308:data<=16'd7195;
      29309:data<=16'd6946;
      29310:data<=16'd6572;
      29311:data<=16'd6197;
      29312:data<=16'd6381;
      29313:data<=16'd7476;
      29314:data<=16'd8363;
      29315:data<=16'd8805;
      29316:data<=16'd8951;
      29317:data<=16'd8657;
      29318:data<=16'd8087;
      29319:data<=16'd8317;
      29320:data<=16'd9956;
      29321:data<=16'd10428;
      29322:data<=16'd9418;
      29323:data<=16'd9470;
      29324:data<=16'd9367;
      29325:data<=16'd9268;
      29326:data<=16'd10578;
      29327:data<=16'd10969;
      29328:data<=16'd10721;
      29329:data<=16'd10736;
      29330:data<=16'd10009;
      29331:data<=16'd10085;
      29332:data<=16'd10878;
      29333:data<=16'd11254;
      29334:data<=16'd11341;
      29335:data<=16'd10786;
      29336:data<=16'd10890;
      29337:data<=16'd10766;
      29338:data<=16'd10135;
      29339:data<=16'd11740;
      29340:data<=16'd11955;
      29341:data<=16'd10637;
      29342:data<=16'd11461;
      29343:data<=16'd8311;
      29344:data<=16'd3099;
      29345:data<=16'd3700;
      29346:data<=16'd4293;
      29347:data<=16'd3092;
      29348:data<=16'd3827;
      29349:data<=16'd3503;
      29350:data<=16'd3519;
      29351:data<=16'd5178;
      29352:data<=16'd5265;
      29353:data<=16'd5162;
      29354:data<=16'd5486;
      29355:data<=16'd5086;
      29356:data<=16'd4978;
      29357:data<=16'd5477;
      29358:data<=16'd6269;
      29359:data<=16'd6463;
      29360:data<=16'd6611;
      29361:data<=16'd6830;
      29362:data<=16'd5380;
      29363:data<=16'd5551;
      29364:data<=16'd7755;
      29365:data<=16'd7145;
      29366:data<=16'd6394;
      29367:data<=16'd6956;
      29368:data<=16'd5987;
      29369:data<=16'd6235;
      29370:data<=16'd7509;
      29371:data<=16'd7228;
      29372:data<=16'd7297;
      29373:data<=16'd7539;
      29374:data<=16'd7071;
      29375:data<=16'd6875;
      29376:data<=16'd7342;
      29377:data<=16'd8204;
      29378:data<=16'd8005;
      29379:data<=16'd7573;
      29380:data<=16'd7881;
      29381:data<=16'd7460;
      29382:data<=16'd7841;
      29383:data<=16'd8745;
      29384:data<=16'd8164;
      29385:data<=16'd8100;
      29386:data<=16'd7567;
      29387:data<=16'd6337;
      29388:data<=16'd7266;
      29389:data<=16'd7850;
      29390:data<=16'd7726;
      29391:data<=16'd8072;
      29392:data<=16'd6966;
      29393:data<=16'd8819;
      29394:data<=16'd14163;
      29395:data<=16'd15390;
      29396:data<=16'd14075;
      29397:data<=16'd14236;
      29398:data<=16'd13791;
      29399:data<=16'd12922;
      29400:data<=16'd11956;
      29401:data<=16'd10135;
      29402:data<=16'd8924;
      29403:data<=16'd8590;
      29404:data<=16'd7868;
      29405:data<=16'd7018;
      29406:data<=16'd6977;
      29407:data<=16'd6263;
      29408:data<=16'd4053;
      29409:data<=16'd3054;
      29410:data<=16'd2893;
      29411:data<=16'd2174;
      29412:data<=16'd2591;
      29413:data<=16'd1839;
      29414:data<=-16'd828;
      29415:data<=-16'd996;
      29416:data<=-16'd234;
      29417:data<=-16'd946;
      29418:data<=-16'd1074;
      29419:data<=-16'd1595;
      29420:data<=-16'd2998;
      29421:data<=-16'd3488;
      29422:data<=-16'd3541;
      29423:data<=-16'd3676;
      29424:data<=-16'd3952;
      29425:data<=-16'd4413;
      29426:data<=-16'd5039;
      29427:data<=-16'd6091;
      29428:data<=-16'd6326;
      29429:data<=-16'd5946;
      29430:data<=-16'd6197;
      29431:data<=-16'd6109;
      29432:data<=-16'd6686;
      29433:data<=-16'd8208;
      29434:data<=-16'd8373;
      29435:data<=-16'd8205;
      29436:data<=-16'd7888;
      29437:data<=-16'd7203;
      29438:data<=-16'd8563;
      29439:data<=-16'd9643;
      29440:data<=-16'd9000;
      29441:data<=-16'd9039;
      29442:data<=-16'd8281;
      29443:data<=-16'd9673;
      29444:data<=-16'd16207;
      29445:data<=-16'd19775;
      29446:data<=-16'd18457;
      29447:data<=-16'd18157;
      29448:data<=-16'd17858;
      29449:data<=-16'd16891;
      29450:data<=-16'd16985;
      29451:data<=-16'd17320;
      29452:data<=-16'd17670;
      29453:data<=-16'd16956;
      29454:data<=-16'd15602;
      29455:data<=-16'd15520;
      29456:data<=-16'd14854;
      29457:data<=-16'd14348;
      29458:data<=-16'd15361;
      29459:data<=-16'd14692;
      29460:data<=-16'd13709;
      29461:data<=-16'd14069;
      29462:data<=-16'd12881;
      29463:data<=-16'd12185;
      29464:data<=-16'd13288;
      29465:data<=-16'd12881;
      29466:data<=-16'd12179;
      29467:data<=-16'd12322;
      29468:data<=-16'd11253;
      29469:data<=-16'd10525;
      29470:data<=-16'd11682;
      29471:data<=-16'd12284;
      29472:data<=-16'd11489;
      29473:data<=-16'd10969;
      29474:data<=-16'd10392;
      29475:data<=-16'd9454;
      29476:data<=-16'd9972;
      29477:data<=-16'd10649;
      29478:data<=-16'd9632;
      29479:data<=-16'd9360;
      29480:data<=-16'd9524;
      29481:data<=-16'd8100;
      29482:data<=-16'd7958;
      29483:data<=-16'd9344;
      29484:data<=-16'd8813;
      29485:data<=-16'd7879;
      29486:data<=-16'd8164;
      29487:data<=-16'd7251;
      29488:data<=-16'd6501;
      29489:data<=-16'd7924;
      29490:data<=-16'd7746;
      29491:data<=-16'd6485;
      29492:data<=-16'd7527;
      29493:data<=-16'd5312;
      29494:data<=16'd1155;
      29495:data<=16'd3732;
      29496:data<=16'd3212;
      29497:data<=16'd3322;
      29498:data<=16'd2852;
      29499:data<=16'd3363;
      29500:data<=16'd4082;
      29501:data<=16'd3927;
      29502:data<=16'd5606;
      29503:data<=16'd6401;
      29504:data<=16'd5353;
      29505:data<=16'd5888;
      29506:data<=16'd5839;
      29507:data<=16'd5650;
      29508:data<=16'd7407;
      29509:data<=16'd7395;
      29510:data<=16'd6402;
      29511:data<=16'd6972;
      29512:data<=16'd6998;
      29513:data<=16'd7228;
      29514:data<=16'd8486;
      29515:data<=16'd8711;
      29516:data<=16'd8316;
      29517:data<=16'd8316;
      29518:data<=16'd8087;
      29519:data<=16'd7976;
      29520:data<=16'd9179;
      29521:data<=16'd10308;
      29522:data<=16'd9643;
      29523:data<=16'd9342;
      29524:data<=16'd9458;
      29525:data<=16'd8296;
      29526:data<=16'd8775;
      29527:data<=16'd10454;
      29528:data<=16'd9926;
      29529:data<=16'd9483;
      29530:data<=16'd9729;
      29531:data<=16'd8900;
      29532:data<=16'd9362;
      29533:data<=16'd10865;
      29534:data<=16'd10507;
      29535:data<=16'd9820;
      29536:data<=16'd10072;
      29537:data<=16'd9359;
      29538:data<=16'd8881;
      29539:data<=16'd10381;
      29540:data<=16'd10442;
      29541:data<=16'd9303;
      29542:data<=16'd10508;
      29543:data<=16'd8836;
      29544:data<=16'd2687;
      29545:data<=16'd895;
      29546:data<=16'd2783;
      29547:data<=16'd2532;
      29548:data<=16'd2613;
      29549:data<=16'd2921;
      29550:data<=16'd1676;
      29551:data<=16'd2220;
      29552:data<=16'd3802;
      29553:data<=16'd3494;
      29554:data<=16'd3483;
      29555:data<=16'd4179;
      29556:data<=16'd3368;
      29557:data<=16'd3024;
      29558:data<=16'd4520;
      29559:data<=16'd4983;
      29560:data<=16'd4684;
      29561:data<=16'd5241;
      29562:data<=16'd4555;
      29563:data<=16'd3489;
      29564:data<=16'd4610;
      29565:data<=16'd5823;
      29566:data<=16'd5727;
      29567:data<=16'd5319;
      29568:data<=16'd4664;
      29569:data<=16'd4314;
      29570:data<=16'd4939;
      29571:data<=16'd5988;
      29572:data<=16'd6125;
      29573:data<=16'd5312;
      29574:data<=16'd5101;
      29575:data<=16'd4902;
      29576:data<=16'd4711;
      29577:data<=16'd5880;
      29578:data<=16'd6205;
      29579:data<=16'd5715;
      29580:data<=16'd6223;
      29581:data<=16'd5335;
      29582:data<=16'd4628;
      29583:data<=16'd6360;
      29584:data<=16'd6786;
      29585:data<=16'd6382;
      29586:data<=16'd6423;
      29587:data<=16'd4907;
      29588:data<=16'd4719;
      29589:data<=16'd6351;
      29590:data<=16'd6640;
      29591:data<=16'd6498;
      29592:data<=16'd5444;
      29593:data<=16'd5333;
      29594:data<=16'd9966;
      29595:data<=16'd13415;
      29596:data<=16'd12198;
      29597:data<=16'd11506;
      29598:data<=16'd11215;
      29599:data<=16'd10323;
      29600:data<=16'd10401;
      29601:data<=16'd9042;
      29602:data<=16'd6849;
      29603:data<=16'd6687;
      29604:data<=16'd6169;
      29605:data<=16'd4707;
      29606:data<=16'd4576;
      29607:data<=16'd4284;
      29608:data<=16'd2648;
      29609:data<=16'd1644;
      29610:data<=16'd1619;
      29611:data<=16'd1248;
      29612:data<=16'd782;
      29613:data<=16'd611;
      29614:data<=-16'd284;
      29615:data<=-16'd1797;
      29616:data<=-16'd2529;
      29617:data<=-16'd2463;
      29618:data<=-16'd2291;
      29619:data<=-16'd2217;
      29620:data<=-16'd3080;
      29621:data<=-16'd4702;
      29622:data<=-16'd4989;
      29623:data<=-16'd4541;
      29624:data<=-16'd5204;
      29625:data<=-16'd5360;
      29626:data<=-16'd5470;
      29627:data<=-16'd7279;
      29628:data<=-16'd7649;
      29629:data<=-16'd6716;
      29630:data<=-16'd7342;
      29631:data<=-16'd6977;
      29632:data<=-16'd6422;
      29633:data<=-16'd8202;
      29634:data<=-16'd8822;
      29635:data<=-16'd8580;
      29636:data<=-16'd9224;
      29637:data<=-16'd8316;
      29638:data<=-16'd7908;
      29639:data<=-16'd9467;
      29640:data<=-16'd10125;
      29641:data<=-16'd10378;
      29642:data<=-16'd10270;
      29643:data<=-16'd9922;
      29644:data<=-16'd12994;
      29645:data<=-16'd18078;
      29646:data<=-16'd20137;
      29647:data<=-16'd19246;
      29648:data<=-16'd18374;
      29649:data<=-16'd18218;
      29650:data<=-16'd17585;
      29651:data<=-16'd17252;
      29652:data<=-16'd18058;
      29653:data<=-16'd18008;
      29654:data<=-16'd17186;
      29655:data<=-16'd16913;
      29656:data<=-16'd16122;
      29657:data<=-16'd15377;
      29658:data<=-16'd15966;
      29659:data<=-16'd16595;
      29660:data<=-16'd16269;
      29661:data<=-16'd15464;
      29662:data<=-16'd14556;
      29663:data<=-16'd13866;
      29664:data<=-16'd14393;
      29665:data<=-16'd15493;
      29666:data<=-16'd14792;
      29667:data<=-16'd13565;
      29668:data<=-16'd13540;
      29669:data<=-16'd12918;
      29670:data<=-16'd12686;
      29671:data<=-16'd13802;
      29672:data<=-16'd13532;
      29673:data<=-16'd12662;
      29674:data<=-16'd12375;
      29675:data<=-16'd11154;
      29676:data<=-16'd10743;
      29677:data<=-16'd11826;
      29678:data<=-16'd11873;
      29679:data<=-16'd11283;
      29680:data<=-16'd10883;
      29681:data<=-16'd10073;
      29682:data<=-16'd9785;
      29683:data<=-16'd10642;
      29684:data<=-16'd11298;
      29685:data<=-16'd10437;
      29686:data<=-16'd9169;
      29687:data<=-16'd8925;
      29688:data<=-16'd8499;
      29689:data<=-16'd8311;
      29690:data<=-16'd9283;
      29691:data<=-16'd8663;
      29692:data<=-16'd7606;
      29693:data<=-16'd8167;
      29694:data<=-16'd4877;
      29695:data<=16'd1494;
      29696:data<=16'd3024;
      29697:data<=16'd1657;
      29698:data<=16'd1820;
      29699:data<=16'd1952;
      29700:data<=16'd2208;
      29701:data<=16'd3015;
      29702:data<=16'd3845;
      29703:data<=16'd4848;
      29704:data<=16'd4733;
      29705:data<=16'd4513;
      29706:data<=16'd5245;
      29707:data<=16'd5086;
      29708:data<=16'd5604;
      29709:data<=16'd7365;
      29710:data<=16'd7441;
      29711:data<=16'd6959;
      29712:data<=16'd6963;
      29713:data<=16'd6617;
      29714:data<=16'd7451;
      29715:data<=16'd8672;
      29716:data<=16'd8367;
      29717:data<=16'd8029;
      29718:data<=16'd8023;
      29719:data<=16'd7558;
      29720:data<=16'd8191;
      29721:data<=16'd9897;
      29722:data<=16'd10044;
      29723:data<=16'd9407;
      29724:data<=16'd9585;
      29725:data<=16'd8681;
      29726:data<=16'd8067;
      29727:data<=16'd9768;
      29728:data<=16'd10320;
      29729:data<=16'd9688;
      29730:data<=16'd10087;
      29731:data<=16'd9500;
      29732:data<=16'd8796;
      29733:data<=16'd10073;
      29734:data<=16'd11173;
      29735:data<=16'd10548;
      29736:data<=16'd9614;
      29737:data<=16'd9793;
      29738:data<=16'd9527;
      29739:data<=16'd9118;
      29740:data<=16'd10810;
      29741:data<=16'd10730;
      29742:data<=16'd9317;
      29743:data<=16'd10683;
      29744:data<=16'd7820;
      29745:data<=16'd1469;
      29746:data<=16'd1659;
      29747:data<=16'd3721;
      29748:data<=16'd3344;
      29749:data<=16'd3858;
      29750:data<=16'd2940;
      29751:data<=16'd2205;
      29752:data<=16'd4428;
      29753:data<=16'd5570;
      29754:data<=16'd5248;
      29755:data<=16'd4927;
      29756:data<=16'd4168;
      29757:data<=16'd4065;
      29758:data<=16'd5086;
      29759:data<=16'd6357;
      29760:data<=16'd6316;
      29761:data<=16'd5688;
      29762:data<=16'd5899;
      29763:data<=16'd4995;
      29764:data<=16'd4645;
      29765:data<=16'd6630;
      29766:data<=16'd7145;
      29767:data<=16'd6616;
      29768:data<=16'd6493;
      29769:data<=16'd5432;
      29770:data<=16'd5500;
      29771:data<=16'd6833;
      29772:data<=16'd7406;
      29773:data<=16'd7341;
      29774:data<=16'd6719;
      29775:data<=16'd6746;
      29776:data<=16'd7356;
      29777:data<=16'd7800;
      29778:data<=16'd8631;
      29779:data<=16'd8102;
      29780:data<=16'd7233;
      29781:data<=16'd7409;
      29782:data<=16'd6320;
      29783:data<=16'd6626;
      29784:data<=16'd8504;
      29785:data<=16'd8119;
      29786:data<=16'd8082;
      29787:data<=16'd7856;
      29788:data<=16'd6422;
      29789:data<=16'd7771;
      29790:data<=16'd8990;
      29791:data<=16'd8622;
      29792:data<=16'd8868;
      29793:data<=16'd7436;
      29794:data<=16'd8862;
      29795:data<=16'd14963;
      29796:data<=16'd16395;
      29797:data<=16'd13993;
      29798:data<=16'd13759;
      29799:data<=16'd13273;
      29800:data<=16'd12354;
      29801:data<=16'd12314;
      29802:data<=16'd10771;
      29803:data<=16'd8387;
      29804:data<=16'd7861;
      29805:data<=16'd7979;
      29806:data<=16'd7233;
      29807:data<=16'd6877;
      29808:data<=16'd5893;
      29809:data<=16'd3751;
      29810:data<=16'd3513;
      29811:data<=16'd3697;
      29812:data<=16'd2588;
      29813:data<=16'd2875;
      29814:data<=16'd2569;
      29815:data<=16'd490;
      29816:data<=-16'd118;
      29817:data<=-16'd314;
      29818:data<=-16'd550;
      29819:data<=16'd218;
      29820:data<=-16'd382;
      29821:data<=-16'd2080;
      29822:data<=-16'd2899;
      29823:data<=-16'd3240;
      29824:data<=-16'd3410;
      29825:data<=-16'd3503;
      29826:data<=-16'd3662;
      29827:data<=-16'd4843;
      29828:data<=-16'd6443;
      29829:data<=-16'd5868;
      29830:data<=-16'd5234;
      29831:data<=-16'd5882;
      29832:data<=-16'd5210;
      29833:data<=-16'd5489;
      29834:data<=-16'd7294;
      29835:data<=-16'd7336;
      29836:data<=-16'd7288;
      29837:data<=-16'd7348;
      29838:data<=-16'd6496;
      29839:data<=-16'd7277;
      29840:data<=-16'd8525;
      29841:data<=-16'd9063;
      29842:data<=-16'd9512;
      29843:data<=-16'd8102;
      29844:data<=-16'd8997;
      29845:data<=-16'd15217;
      29846:data<=-16'd19082;
      29847:data<=-16'd18436;
      29848:data<=-16'd17940;
      29849:data<=-16'd17194;
      29850:data<=-16'd16140;
      29851:data<=-16'd16236;
      29852:data<=-16'd16759;
      29853:data<=-16'd17227;
      29854:data<=-16'd16810;
      29855:data<=-16'd16037;
      29856:data<=-16'd15849;
      29857:data<=-16'd14684;
      29858:data<=-16'd14287;
      29859:data<=-16'd15945;
      29860:data<=-16'd15822;
      29861:data<=-16'd14739;
      29862:data<=-16'd14621;
      29863:data<=-16'd13189;
      29864:data<=-16'd12789;
      29865:data<=-16'd14650;
      29866:data<=-16'd14600;
      29867:data<=-16'd13436;
      29868:data<=-16'd12995;
      29869:data<=-16'd11925;
      29870:data<=-16'd11671;
      29871:data<=-16'd12795;
      29872:data<=-16'd13097;
      29873:data<=-16'd12481;
      29874:data<=-16'd11664;
      29875:data<=-16'd10537;
      29876:data<=-16'd9577;
      29877:data<=-16'd9838;
      29878:data<=-16'd10839;
      29879:data<=-16'd10748;
      29880:data<=-16'd10043;
      29881:data<=-16'd9541;
      29882:data<=-16'd8683;
      29883:data<=-16'd9021;
      29884:data<=-16'd10361;
      29885:data<=-16'd9847;
      29886:data<=-16'd8883;
      29887:data<=-16'd8802;
      29888:data<=-16'd7699;
      29889:data<=-16'd7385;
      29890:data<=-16'd8906;
      29891:data<=-16'd8429;
      29892:data<=-16'd7212;
      29893:data<=-16'd8103;
      29894:data<=-16'd5982;
      29895:data<=16'd82;
      29896:data<=16'd3015;
      29897:data<=16'd2660;
      29898:data<=16'd2675;
      29899:data<=16'd2599;
      29900:data<=16'd2861;
      29901:data<=16'd3457;
      29902:data<=16'd3818;
      29903:data<=16'd4977;
      29904:data<=16'd5391;
      29905:data<=16'd4898;
      29906:data<=16'd5453;
      29907:data<=16'd5611;
      29908:data<=16'd5638;
      29909:data<=16'd6714;
      29910:data<=16'd7203;
      29911:data<=16'd7512;
      29912:data<=16'd7618;
      29913:data<=16'd6786;
      29914:data<=16'd7156;
      29915:data<=16'd8487;
      29916:data<=16'd8909;
      29917:data<=16'd8819;
      29918:data<=16'd8580;
      29919:data<=16'd8170;
      29920:data<=16'd7934;
      29921:data<=16'd9051;
      29922:data<=16'd10587;
      29923:data<=16'd9799;
      29924:data<=16'd8921;
      29925:data<=16'd9265;
      29926:data<=16'd8419;
      29927:data<=16'd8483;
      29928:data<=16'd9667;
      29929:data<=16'd9426;
      29930:data<=16'd9564;
      29931:data<=16'd9453;
      29932:data<=16'd8263;
      29933:data<=16'd8801;
      29934:data<=16'd10022;
      29935:data<=16'd10290;
      29936:data<=16'd10140;
      29937:data<=16'd9338;
      29938:data<=16'd8595;
      29939:data<=16'd8663;
      29940:data<=16'd9896;
      29941:data<=16'd10481;
      29942:data<=16'd9045;
      29943:data<=16'd9421;
      29944:data<=16'd8978;
      29945:data<=16'd3175;
      29946:data<=16'd287;
      29947:data<=16'd2508;
      29948:data<=16'd2710;
      29949:data<=16'd2655;
      29950:data<=16'd3002;
      29951:data<=16'd1541;
      29952:data<=16'd2369;
      29953:data<=16'd4708;
      29954:data<=16'd4543;
      29955:data<=16'd4241;
      29956:data<=16'd4614;
      29957:data<=16'd3703;
      29958:data<=16'd3630;
      29959:data<=16'd5620;
      29960:data<=16'd6061;
      29961:data<=16'd4781;
      29962:data<=16'd4945;
      29963:data<=16'd5080;
      29964:data<=16'd4795;
      29965:data<=16'd6123;
      29966:data<=16'd6670;
      29967:data<=16'd6087;
      29968:data<=16'd6284;
      29969:data<=16'd5618;
      29970:data<=16'd4981;
      29971:data<=16'd6023;
      29972:data<=16'd6769;
      29973:data<=16'd6807;
      29974:data<=16'd6672;
      29975:data<=16'd6197;
      29976:data<=16'd5941;
      29977:data<=16'd6488;
      29978:data<=16'd7706;
      29979:data<=16'd7962;
      29980:data<=16'd7288;
      29981:data<=16'd7341;
      29982:data<=16'd7063;
      29983:data<=16'd6893;
      29984:data<=16'd7949;
      29985:data<=16'd7900;
      29986:data<=16'd7329;
      29987:data<=16'd7588;
      29988:data<=16'd7028;
      29989:data<=16'd6804;
      29990:data<=16'd7529;
      29991:data<=16'd7794;
      29992:data<=16'd8228;
      29993:data<=16'd7617;
      29994:data<=16'd6843;
      29995:data<=16'd10361;
      29996:data<=16'd14504;
      29997:data<=16'd14108;
      29998:data<=16'd12972;
      29999:data<=16'd12731;
      30000:data<=16'd11627;
      30001:data<=16'd11359;
      30002:data<=16'd10668;
      30003:data<=16'd8232;
      30004:data<=16'd7253;
      30005:data<=16'd6921;
      30006:data<=16'd5979;
      30007:data<=16'd6249;
      30008:data<=16'd5406;
      30009:data<=16'd3087;
      30010:data<=16'd2628;
      30011:data<=16'd2790;
      30012:data<=16'd2446;
      30013:data<=16'd2258;
      30014:data<=16'd1160;
      30015:data<=-16'd312;
      30016:data<=-16'd1121;
      30017:data<=-16'd1468;
      30018:data<=-16'd1651;
      30019:data<=-16'd1915;
      30020:data<=-16'd1853;
      30021:data<=-16'd2701;
      30022:data<=-16'd4645;
      30023:data<=-16'd4871;
      30024:data<=-16'd4437;
      30025:data<=-16'd4757;
      30026:data<=-16'd4419;
      30027:data<=-16'd5053;
      30028:data<=-16'd6689;
      30029:data<=-16'd7025;
      30030:data<=-16'd6974;
      30031:data<=-16'd6802;
      30032:data<=-16'd6326;
      30033:data<=-16'd6904;
      30034:data<=-16'd8193;
      30035:data<=-16'd8710;
      30036:data<=-16'd8237;
      30037:data<=-16'd8267;
      30038:data<=-16'd8713;
      30039:data<=-16'd8422;
      30040:data<=-16'd9039;
      30041:data<=-16'd10228;
      30042:data<=-16'd10384;
      30043:data<=-16'd10158;
      30044:data<=-16'd9179;
      30045:data<=-16'd10983;
      30046:data<=-16'd17273;
      30047:data<=-16'd20058;
      30048:data<=-16'd18801;
      30049:data<=-16'd19089;
      30050:data<=-16'd18516;
      30051:data<=-16'd16977;
      30052:data<=-16'd17420;
      30053:data<=-16'd18271;
      30054:data<=-16'd18210;
      30055:data<=-16'd17347;
      30056:data<=-16'd16838;
      30057:data<=-16'd16735;
      30058:data<=-16'd15799;
      30059:data<=-16'd15984;
      30060:data<=-16'd16842;
      30061:data<=-16'd16271;
      30062:data<=-16'd16130;
      30063:data<=-16'd15625;
      30064:data<=-16'd14016;
      30065:data<=-16'd14252;
      30066:data<=-16'd15374;
      30067:data<=-16'd15112;
      30068:data<=-16'd14374;
      30069:data<=-16'd14002;
      30070:data<=-16'd13588;
      30071:data<=-16'd13305;
      30072:data<=-16'd14032;
      30073:data<=-16'd13993;
      30074:data<=-16'd12756;
      30075:data<=-16'd12847;
      30076:data<=-16'd12389;
      30077:data<=-16'd11402;
      30078:data<=-16'd12498;
      30079:data<=-16'd12387;
      30080:data<=-16'd11259;
      30081:data<=-16'd11485;
      30082:data<=-16'd10580;
      30083:data<=-16'd10097;
      30084:data<=-16'd11001;
      30085:data<=-16'd10901;
      30086:data<=-16'd10869;
      30087:data<=-16'd10358;
      30088:data<=-16'd9113;
      30089:data<=-16'd8627;
      30090:data<=-16'd8520;
      30091:data<=-16'd9542;
      30092:data<=-16'd9451;
      30093:data<=-16'd8125;
      30094:data<=-16'd9276;
      30095:data<=-16'd6636;
      30096:data<=16'd472;
      30097:data<=16'd1959;
      30098:data<=16'd1011;
      30099:data<=16'd2396;
      30100:data<=16'd2106;
      30101:data<=16'd1630;
      30102:data<=16'd2663;
      30103:data<=16'd4002;
      30104:data<=16'd5109;
      30105:data<=16'd4517;
      30106:data<=16'd4223;
      30107:data<=16'd4962;
      30108:data<=16'd4763;
      30109:data<=16'd5559;
      30110:data<=16'd6872;
      30111:data<=16'd6831;
      30112:data<=16'd6957;
      30113:data<=16'd6646;
      30114:data<=16'd5868;
      30115:data<=16'd6677;
      30116:data<=16'd8187;
      30117:data<=16'd8404;
      30118:data<=16'd7659;
      30119:data<=16'd7708;
      30120:data<=16'd7929;
      30121:data<=16'd7821;
      30122:data<=16'd9121;
      30123:data<=16'd9670;
      30124:data<=16'd8564;
      30125:data<=16'd8889;
      30126:data<=16'd8893;
      30127:data<=16'd8258;
      30128:data<=16'd9385;
      30129:data<=16'd9673;
      30130:data<=16'd9007;
      30131:data<=16'd9262;
      30132:data<=16'd8836;
      30133:data<=16'd8478;
      30134:data<=16'd9367;
      30135:data<=16'd10034;
      30136:data<=16'd9679;
      30137:data<=16'd9075;
      30138:data<=16'd9003;
      30139:data<=16'd8254;
      30140:data<=16'd8284;
      30141:data<=16'd10313;
      30142:data<=16'd9492;
      30143:data<=16'd8237;
      30144:data<=16'd10378;
      30145:data<=16'd7602;
      30146:data<=16'd1454;
      30147:data<=16'd1516;
      30148:data<=16'd2872;
      30149:data<=16'd1851;
      30150:data<=16'd2162;
      30151:data<=16'd2228;
      30152:data<=16'd2003;
      30153:data<=16'd3189;
      30154:data<=16'd3874;
      30155:data<=16'd3858;
      30156:data<=16'd3953;
      30157:data<=16'd3782;
      30158:data<=16'd3598;
      30159:data<=16'd4296;
      30160:data<=16'd5498;
      30161:data<=16'd5342;
      30162:data<=16'd4839;
      30163:data<=16'd5327;
      30164:data<=16'd5048;
      30165:data<=16'd5189;
      30166:data<=16'd6522;
      30167:data<=16'd6484;
      30168:data<=16'd6164;
      30169:data<=16'd6213;
      30170:data<=16'd5551;
      30171:data<=16'd6059;
      30172:data<=16'd7089;
      30173:data<=16'd7004;
      30174:data<=16'd7053;
      30175:data<=16'd6910;
      30176:data<=16'd6425;
      30177:data<=16'd6555;
      30178:data<=16'd7241;
      30179:data<=16'd8078;
      30180:data<=16'd7847;
      30181:data<=16'd7275;
      30182:data<=16'd7354;
      30183:data<=16'd6699;
      30184:data<=16'd6937;
      30185:data<=16'd8244;
      30186:data<=16'd7796;
      30187:data<=16'd7517;
      30188:data<=16'd7689;
      30189:data<=16'd6949;
      30190:data<=16'd7597;
      30191:data<=16'd8172;
      30192:data<=16'd7937;
      30193:data<=16'd8263;
      30194:data<=16'd6833;
      30195:data<=16'd7908;
      30196:data<=16'd13825;
      30197:data<=16'd15402;
      30198:data<=16'd13226;
      30199:data<=16'd13602;
      30200:data<=16'd13191;
      30201:data<=16'd12032;
      30202:data<=16'd12217;
      30203:data<=16'd10584;
      30204:data<=16'd8241;
      30205:data<=16'd7803;
      30206:data<=16'd7667;
      30207:data<=16'd7210;
      30208:data<=16'd6889;
      30209:data<=16'd5736;
      30210:data<=16'd3738;
      30211:data<=16'd2971;
      30212:data<=16'd3275;
      30213:data<=16'd2795;
      30214:data<=16'd2617;
      30215:data<=16'd2328;
      30216:data<=16'd561;
      30217:data<=-16'd196;
      30218:data<=-16'd74;
      30219:data<=-16'd591;
      30220:data<=-16'd305;
      30221:data<=-16'd605;
      30222:data<=-16'd2259;
      30223:data<=-16'd3001;
      30224:data<=-16'd3312;
      30225:data<=-16'd3595;
      30226:data<=-16'd3201;
      30227:data<=-16'd3127;
      30228:data<=-16'd4062;
      30229:data<=-16'd5395;
      30230:data<=-16'd5650;
      30231:data<=-16'd5274;
      30232:data<=-16'd5407;
      30233:data<=-16'd5112;
      30234:data<=-16'd5887;
      30235:data<=-16'd7605;
      30236:data<=-16'd6948;
      30237:data<=-16'd6344;
      30238:data<=-16'd7024;
      30239:data<=-16'd6734;
      30240:data<=-16'd7486;
      30241:data<=-16'd8507;
      30242:data<=-16'd8341;
      30243:data<=-16'd8601;
      30244:data<=-16'd7483;
      30245:data<=-16'd8167;
      30246:data<=-16'd14063;
      30247:data<=-16'd17529;
      30248:data<=-16'd16874;
      30249:data<=-16'd17120;
      30250:data<=-16'd16733;
      30251:data<=-16'd15462;
      30252:data<=-16'd15344;
      30253:data<=-16'd15951;
      30254:data<=-16'd16624;
      30255:data<=-16'd16070;
      30256:data<=-16'd15238;
      30257:data<=-16'd15159;
      30258:data<=-16'd14216;
      30259:data<=-16'd14013;
      30260:data<=-16'd14922;
      30261:data<=-16'd14352;
      30262:data<=-16'd13758;
      30263:data<=-16'd13718;
      30264:data<=-16'd12869;
      30265:data<=-16'd12747;
      30266:data<=-16'd13579;
      30267:data<=-16'd13767;
      30268:data<=-16'd13223;
      30269:data<=-16'd12622;
      30270:data<=-16'd11982;
      30271:data<=-16'd11147;
      30272:data<=-16'd11473;
      30273:data<=-16'd12399;
      30274:data<=-16'd11682;
      30275:data<=-16'd11035;
      30276:data<=-16'd10988;
      30277:data<=-16'd9962;
      30278:data<=-16'd10058;
      30279:data<=-16'd11006;
      30280:data<=-16'd10407;
      30281:data<=-16'd9752;
      30282:data<=-16'd9371;
      30283:data<=-16'd8636;
      30284:data<=-16'd8968;
      30285:data<=-16'd9759;
      30286:data<=-16'd9488;
      30287:data<=-16'd8883;
      30288:data<=-16'd8528;
      30289:data<=-16'd7479;
      30290:data<=-16'd6751;
      30291:data<=-16'd8085;
      30292:data<=-16'd8423;
      30293:data<=-16'd7125;
      30294:data<=-16'd7796;
      30295:data<=-16'd6314;
      30296:data<=-16'd282;
      30297:data<=16'd2866;
      30298:data<=16'd2259;
      30299:data<=16'd2369;
      30300:data<=16'd2798;
      30301:data<=16'd3092;
      30302:data<=16'd3366;
      30303:data<=16'd4179;
      30304:data<=16'd5773;
      30305:data<=16'd5721;
      30306:data<=16'd5256;
      30307:data<=16'd6140;
      30308:data<=16'd6037;
      30309:data<=16'd6097;
      30310:data<=16'd7321;
      30311:data<=16'd7524;
      30312:data<=16'd7595;
      30313:data<=16'd7870;
      30314:data<=16'd7656;
      30315:data<=16'd8240;
      30316:data<=16'd9183;
      30317:data<=16'd9586;
      30318:data<=16'd9559;
      30319:data<=16'd9266;
      30320:data<=16'd9116;
      30321:data<=16'd8669;
      30322:data<=16'd9024;
      30323:data<=16'd10442;
      30324:data<=16'd10161;
      30325:data<=16'd9539;
      30326:data<=16'd9876;
      30327:data<=16'd9177;
      30328:data<=16'd9508;
      30329:data<=16'd10684;
      30330:data<=16'd9832;
      30331:data<=16'd9424;
      30332:data<=16'd9639;
      30333:data<=16'd8974;
      30334:data<=16'd9741;
      30335:data<=16'd10869;
      30336:data<=16'd10477;
      30337:data<=16'd10063;
      30338:data<=16'd9823;
      30339:data<=16'd9283;
      30340:data<=16'd8824;
      30341:data<=16'd9667;
      30342:data<=16'd11010;
      30343:data<=16'd10255;
      30344:data<=16'd10069;
      30345:data<=16'd9949;
      30346:data<=16'd4821;
      30347:data<=16'd1249;
      30348:data<=16'd3553;
      30349:data<=16'd3811;
      30350:data<=16'd2672;
      30351:data<=16'd3389;
      30352:data<=16'd2649;
      30353:data<=16'd2942;
      30354:data<=16'd4833;
      30355:data<=16'd4473;
      30356:data<=16'd4472;
      30357:data<=16'd5172;
      30358:data<=16'd4249;
      30359:data<=16'd4520;
      30360:data<=16'd6012;
      30361:data<=16'd6131;
      30362:data<=16'd5941;
      30363:data<=16'd6073;
      30364:data<=16'd5421;
      30365:data<=16'd4675;
      30366:data<=16'd5658;
      30367:data<=16'd7103;
      30368:data<=16'd6648;
      30369:data<=16'd5970;
      30370:data<=16'd6043;
      30371:data<=16'd5579;
      30372:data<=16'd5971;
      30373:data<=16'd7186;
      30374:data<=16'd7181;
      30375:data<=16'd6737;
      30376:data<=16'd6366;
      30377:data<=16'd5868;
      30378:data<=16'd6331;
      30379:data<=16'd7389;
      30380:data<=16'd7762;
      30381:data<=16'd7605;
      30382:data<=16'd7471;
      30383:data<=16'd7025;
      30384:data<=16'd6693;
      30385:data<=16'd7645;
      30386:data<=16'd8310;
      30387:data<=16'd7691;
      30388:data<=16'd7602;
      30389:data<=16'd7353;
      30390:data<=16'd6877;
      30391:data<=16'd7627;
      30392:data<=16'd7864;
      30393:data<=16'd7670;
      30394:data<=16'd7344;
      30395:data<=16'd6117;
      30396:data<=16'd8649;
      30397:data<=16'd13644;
      30398:data<=16'd13773;
      30399:data<=16'd12419;
      30400:data<=16'd12680;
      30401:data<=16'd11217;
      30402:data<=16'd10163;
      30403:data<=16'd9958;
      30404:data<=16'd8196;
      30405:data<=16'd7066;
      30406:data<=16'd6370;
      30407:data<=16'd5069;
      30408:data<=16'd4816;
      30409:data<=16'd4323;
      30410:data<=16'd2860;
      30411:data<=16'd1962;
      30412:data<=16'd1354;
      30413:data<=16'd845;
      30414:data<=16'd930;
      30415:data<=16'd977;
      30416:data<=-16'd173;
      30417:data<=-16'd1800;
      30418:data<=-16'd1971;
      30419:data<=-16'd1821;
      30420:data<=-16'd2531;
      30421:data<=-16'd2851;
      30422:data<=-16'd3570;
      30423:data<=-16'd4861;
      30424:data<=-16'd5092;
      30425:data<=-16'd5096;
      30426:data<=-16'd5313;
      30427:data<=-16'd5263;
      30428:data<=-16'd5755;
      30429:data<=-16'd6522;
      30430:data<=-16'd6886;
      30431:data<=-16'd7012;
      30432:data<=-16'd7204;
      30433:data<=-16'd7347;
      30434:data<=-16'd7003;
      30435:data<=-16'd7473;
      30436:data<=-16'd8763;
      30437:data<=-16'd8692;
      30438:data<=-16'd8519;
      30439:data<=-16'd8981;
      30440:data<=-16'd8693;
      30441:data<=-16'd9174;
      30442:data<=-16'd10164;
      30443:data<=-16'd10284;
      30444:data<=-16'd10255;
      30445:data<=-16'd9461;
      30446:data<=-16'd11016;
      30447:data<=-16'd16986;
      30448:data<=-16'd20028;
      30449:data<=-16'd18668;
      30450:data<=-16'd18697;
      30451:data<=-16'd18675;
      30452:data<=-16'd17171;
      30453:data<=-16'd17291;
      30454:data<=-16'd18483;
      30455:data<=-16'd18406;
      30456:data<=-16'd17337;
      30457:data<=-16'd16782;
      30458:data<=-16'd16427;
      30459:data<=-16'd15609;
      30460:data<=-16'd16137;
      30461:data<=-16'd16983;
      30462:data<=-16'd15773;
      30463:data<=-16'd15135;
      30464:data<=-16'd15403;
      30465:data<=-16'd14254;
      30466:data<=-16'd14167;
      30467:data<=-16'd15546;
      30468:data<=-16'd15226;
      30469:data<=-16'd14245;
      30470:data<=-16'd13782;
      30471:data<=-16'd12842;
      30472:data<=-16'd12833;
      30473:data<=-16'd13805;
      30474:data<=-16'd13420;
      30475:data<=-16'd12757;
      30476:data<=-16'd12604;
      30477:data<=-16'd11242;
      30478:data<=-16'd10740;
      30479:data<=-16'd12289;
      30480:data<=-16'd12404;
      30481:data<=-16'd11386;
      30482:data<=-16'd11028;
      30483:data<=-16'd9988;
      30484:data<=-16'd9427;
      30485:data<=-16'd10498;
      30486:data<=-16'd11054;
      30487:data<=-16'd10572;
      30488:data<=-16'd10061;
      30489:data<=-16'd9491;
      30490:data<=-16'd8517;
      30491:data<=-16'd8463;
      30492:data<=-16'd9899;
      30493:data<=-16'd9647;
      30494:data<=-16'd8487;
      30495:data<=-16'd9010;
      30496:data<=-16'd6029;
      30497:data<=16'd250;
      30498:data<=16'd2062;
      30499:data<=16'd1268;
      30500:data<=16'd1979;
      30501:data<=16'd2378;
      30502:data<=16'd2538;
      30503:data<=16'd2924;
      30504:data<=16'd3644;
      30505:data<=16'd4816;
      30506:data<=16'd4833;
      30507:data<=16'd4861;
      30508:data<=16'd5388;
      30509:data<=16'd4855;
      30510:data<=16'd5551;
      30511:data<=16'd7071;
      30512:data<=16'd6663;
      30513:data<=16'd6557;
      30514:data<=16'd7024;
      30515:data<=16'd6443;
      30516:data<=16'd7003;
      30517:data<=16'd8578;
      30518:data<=16'd8540;
      30519:data<=16'd7774;
      30520:data<=16'd7794;
      30521:data<=16'd7841;
      30522:data<=16'd8076;
      30523:data<=16'd8963;
      30524:data<=16'd9024;
      30525:data<=16'd8561;
      30526:data<=16'd8724;
      30527:data<=16'd8222;
      30528:data<=16'd7975;
      30529:data<=16'd9300;
      30530:data<=16'd9826;
      30531:data<=16'd9198;
      30532:data<=16'd8884;
      30533:data<=16'd8595;
      30534:data<=16'd8337;
      30535:data<=16'd8624;
      30536:data<=16'd9474;
      30537:data<=16'd9632;
      30538:data<=16'd9045;
      30539:data<=16'd9233;
      30540:data<=16'd8523;
      30541:data<=16'd7859;
      30542:data<=16'd9849;
      30543:data<=16'd9956;
      30544:data<=16'd8842;
      30545:data<=16'd10332;
      30546:data<=16'd7506;
      30547:data<=16'd1221;
      30548:data<=16'd978;
      30549:data<=16'd3034;
      30550:data<=16'd2325;
      30551:data<=16'd2052;
      30552:data<=16'd2218;
      30553:data<=16'd2015;
      30554:data<=16'd3107;
      30555:data<=16'd4438;
      30556:data<=16'd3944;
      30557:data<=16'd3178;
      30558:data<=16'd3682;
      30559:data<=16'd3494;
      30560:data<=16'd3544;
      30561:data<=16'd5256;
      30562:data<=16'd5228;
      30563:data<=16'd4470;
      30564:data<=16'd5197;
      30565:data<=16'd4634;
      30566:data<=16'd4593;
      30567:data<=16'd6269;
      30568:data<=16'd6228;
      30569:data<=16'd5955;
      30570:data<=16'd6031;
      30571:data<=16'd4864;
      30572:data<=16'd5140;
      30573:data<=16'd6790;
      30574:data<=16'd7248;
      30575:data<=16'd6884;
      30576:data<=16'd6366;
      30577:data<=16'd5962;
      30578:data<=16'd5695;
      30579:data<=16'd6200;
      30580:data<=16'd7391;
      30581:data<=16'd7177;
      30582:data<=16'd6575;
      30583:data<=16'd6536;
      30584:data<=16'd5711;
      30585:data<=16'd6249;
      30586:data<=16'd7779;
      30587:data<=16'd7404;
      30588:data<=16'd6992;
      30589:data<=16'd6590;
      30590:data<=16'd5723;
      30591:data<=16'd6728;
      30592:data<=16'd7665;
      30593:data<=16'd7477;
      30594:data<=16'd7301;
      30595:data<=16'd5732;
      30596:data<=16'd6887;
      30597:data<=16'd12932;
      30598:data<=16'd15249;
      30599:data<=16'd12751;
      30600:data<=16'd12213;
      30601:data<=16'd12128;
      30602:data<=16'd10783;
      30603:data<=16'd10651;
      30604:data<=16'd9834;
      30605:data<=16'd7696;
      30606:data<=16'd6974;
      30607:data<=16'd6558;
      30608:data<=16'd5723;
      30609:data<=16'd5850;
      30610:data<=16'd5325;
      30611:data<=16'd3700;
      30612:data<=16'd2870;
      30613:data<=16'd2150;
      30614:data<=16'd1333;
      30615:data<=16'd1569;
      30616:data<=16'd1286;
      30617:data<=-16'd375;
      30618:data<=-16'd1328;
      30619:data<=-16'd1357;
      30620:data<=-16'd1700;
      30621:data<=-16'd1698;
      30622:data<=-16'd1595;
      30623:data<=-16'd2968;
      30624:data<=-16'd4444;
      30625:data<=-16'd4435;
      30626:data<=-16'd4407;
      30627:data<=-16'd4510;
      30628:data<=-16'd4153;
      30629:data<=-16'd4966;
      30630:data<=-16'd6270;
      30631:data<=-16'd6111;
      30632:data<=-16'd6100;
      30633:data<=-16'd6549;
      30634:data<=-16'd5924;
      30635:data<=-16'd6140;
      30636:data<=-16'd7562;
      30637:data<=-16'd7802;
      30638:data<=-16'd7765;
      30639:data<=-16'd7803;
      30640:data<=-16'd6996;
      30641:data<=-16'd7370;
      30642:data<=-16'd8654;
      30643:data<=-16'd9091;
      30644:data<=-16'd9085;
      30645:data<=-16'd8038;
      30646:data<=-16'd8722;
      30647:data<=-16'd13941;
      30648:data<=-16'd17890;
      30649:data<=-16'd17676;
      30650:data<=-16'd17311;
      30651:data<=-16'd17344;
      30652:data<=-16'd16656;
      30653:data<=-16'd15558;
      30654:data<=-16'd15515;
      30655:data<=-16'd16991;
      30656:data<=-16'd16691;
      30657:data<=-16'd15317;
      30658:data<=-16'd15411;
      30659:data<=-16'd14495;
      30660:data<=-16'd14170;
      30661:data<=-16'd15987;
      30662:data<=-16'd15534;
      30663:data<=-16'd13860;
      30664:data<=-16'd13430;
      30665:data<=-16'd12707;
      30666:data<=-16'd12797;
      30667:data<=-16'd13720;
      30668:data<=-16'd13665;
      30669:data<=-16'd12892;
      30670:data<=-16'd11947;
      30671:data<=-16'd11603;
      30672:data<=-16'd11445;
      30673:data<=-16'd11388;
      30674:data<=-16'd12148;
      30675:data<=-16'd11676;
      30676:data<=-16'd10621;
      30677:data<=-16'd10575;
      30678:data<=-16'd9403;
      30679:data<=-16'd9072;
      30680:data<=-16'd10693;
      30681:data<=-16'd10496;
      30682:data<=-16'd9523;
      30683:data<=-16'd8971;
      30684:data<=-16'd7771;
      30685:data<=-16'd8125;
      30686:data<=-16'd9558;
      30687:data<=-16'd9260;
      30688:data<=-16'd8081;
      30689:data<=-16'd7624;
      30690:data<=-16'd7365;
      30691:data<=-16'd6816;
      30692:data<=-16'd7497;
      30693:data<=-16'd8204;
      30694:data<=-16'd6834;
      30695:data<=-16'd6664;
      30696:data<=-16'd6129;
      30697:data<=-16'd789;
      30698:data<=16'd3395;
      30699:data<=16'd3162;
      30700:data<=16'd3327;
      30701:data<=16'd4146;
      30702:data<=16'd4244;
      30703:data<=16'd3902;
      30704:data<=16'd3892;
      30705:data<=16'd5350;
      30706:data<=16'd6194;
      30707:data<=16'd6085;
      30708:data<=16'd6501;
      30709:data<=16'd5820;
      30710:data<=16'd5753;
      30711:data<=16'd7861;
      30712:data<=16'd8660;
      30713:data<=16'd8211;
      30714:data<=16'd8144;
      30715:data<=16'd7700;
      30716:data<=16'd7738;
      30717:data<=16'd8892;
      30718:data<=16'd9884;
      30719:data<=16'd9454;
      30720:data<=16'd8546;
      30721:data<=16'd8766;
      30722:data<=16'd8687;
      30723:data<=16'd8634;
      30724:data<=16'd10169;
      30725:data<=16'd10577;
      30726:data<=16'd9905;
      30727:data<=16'd9969;
      30728:data<=16'd9047;
      30729:data<=16'd8969;
      30730:data<=16'd10790;
      30731:data<=16'd10860;
      30732:data<=16'd10279;
      30733:data<=16'd10423;
      30734:data<=16'd9474;
      30735:data<=16'd9652;
      30736:data<=16'd11470;
      30737:data<=16'd11570;
      30738:data<=16'd10633;
      30739:data<=16'd10417;
      30740:data<=16'd9987;
      30741:data<=16'd9376;
      30742:data<=16'd10066;
      30743:data<=16'd11306;
      30744:data<=16'd10789;
      30745:data<=16'd10396;
      30746:data<=16'd10636;
      30747:data<=16'd6246;
      30748:data<=16'd1036;
      30749:data<=16'd2519;
      30750:data<=16'd4337;
      30751:data<=16'd2729;
      30752:data<=16'd2748;
      30753:data<=16'd2772;
      30754:data<=16'd2736;
      30755:data<=16'd5053;
      30756:data<=16'd5633;
      30757:data<=16'd4717;
      30758:data<=16'd4881;
      30759:data<=16'd4429;
      30760:data<=16'd4772;
      30761:data<=16'd5935;
      30762:data<=16'd5694;
      30763:data<=16'd5495;
      30764:data<=16'd5524;
      30765:data<=16'd5257;
      30766:data<=16'd5254;
      30767:data<=16'd5651;
      30768:data<=16'd7025;
      30769:data<=16'd7457;
      30770:data<=16'd6496;
      30771:data<=16'd6311;
      30772:data<=16'd5692;
      30773:data<=16'd5944;
      30774:data<=16'd7990;
      30775:data<=16'd7732;
      30776:data<=16'd6689;
      30777:data<=16'd6734;
      30778:data<=16'd5817;
      30779:data<=16'd6197;
      30780:data<=16'd7699;
      30781:data<=16'd7585;
      30782:data<=16'd7227;
      30783:data<=16'd6918;
      30784:data<=16'd6504;
      30785:data<=16'd6608;
      30786:data<=16'd6924;
      30787:data<=16'd7647;
      30788:data<=16'd7805;
      30789:data<=16'd7254;
      30790:data<=16'd6834;
      30791:data<=16'd6448;
      30792:data<=16'd7109;
      30793:data<=16'd7702;
      30794:data<=16'd7460;
      30795:data<=16'd7183;
      30796:data<=16'd5689;
      30797:data<=16'd7890;
      30798:data<=16'd14487;
      30799:data<=16'd15123;
      30800:data<=16'd12225;
      30801:data<=16'd12498;
      30802:data<=16'd11917;
      30803:data<=16'd11530;
      30804:data<=16'd11541;
      30805:data<=16'd8904;
      30806:data<=16'd7539;
      30807:data<=16'd7009;
      30808:data<=16'd5777;
      30809:data<=16'd6375;
      30810:data<=16'd6028;
      30811:data<=16'd4331;
      30812:data<=16'd3580;
      30813:data<=16'd2669;
      30814:data<=16'd2287;
      30815:data<=16'd2205;
      30816:data<=16'd1879;
      30817:data<=16'd1421;
      30818:data<=-16'd811;
      30819:data<=-16'd2184;
      30820:data<=-16'd1480;
      30821:data<=-16'd1418;
      30822:data<=-16'd977;
      30823:data<=-16'd1704;
      30824:data<=-16'd4360;
      30825:data<=-16'd4755;
      30826:data<=-16'd4353;
      30827:data<=-16'd4614;
      30828:data<=-16'd3889;
      30829:data<=-16'd4353;
      30830:data<=-16'd5926;
      30831:data<=-16'd6420;
      30832:data<=-16'd6270;
      30833:data<=-16'd6111;
      30834:data<=-16'd6325;
      30835:data<=-16'd6449;
      30836:data<=-16'd6927;
      30837:data<=-16'd8217;
      30838:data<=-16'd8616;
      30839:data<=-16'd8552;
      30840:data<=-16'd8219;
      30841:data<=-16'd7507;
      30842:data<=-16'd8552;
      30843:data<=-16'd9514;
      30844:data<=-16'd9461;
      30845:data<=-16'd9661;
      30846:data<=-16'd8225;
      30847:data<=-16'd9835;
      30848:data<=-16'd16788;
      30849:data<=-16'd19613;
      30850:data<=-16'd18046;
      30851:data<=-16'd18048;
      30852:data<=-16'd17637;
      30853:data<=-16'd16822;
      30854:data<=-16'd17045;
      30855:data<=-16'd17191;
      30856:data<=-16'd17437;
      30857:data<=-16'd16848;
      30858:data<=-16'd15850;
      30859:data<=-16'd15641;
      30860:data<=-16'd14957;
      30861:data<=-16'd15241;
      30862:data<=-16'd16660;
      30863:data<=-16'd15949;
      30864:data<=-16'd14598;
      30865:data<=-16'd14398;
      30866:data<=-16'd13643;
      30867:data<=-16'd13599;
      30868:data<=-16'd14882;
      30869:data<=-16'd14443;
      30870:data<=-16'd13016;
      30871:data<=-16'd13048;
      30872:data<=-16'd12938;
      30873:data<=-16'd12510;
      30874:data<=-16'd13080;
      30875:data<=-16'd12834;
      30876:data<=-16'd11923;
      30877:data<=-16'd11841;
      30878:data<=-16'd11156;
      30879:data<=-16'd10430;
      30880:data<=-16'd10992;
      30881:data<=-16'd11207;
      30882:data<=-16'd10704;
      30883:data<=-16'd10257;
      30884:data<=-16'd9594;
      30885:data<=-16'd8915;
      30886:data<=-16'd9233;
      30887:data<=-16'd10337;
      30888:data<=-16'd9961;
      30889:data<=-16'd8718;
      30890:data<=-16'd8833;
      30891:data<=-16'd8329;
      30892:data<=-16'd7777;
      30893:data<=-16'd9271;
      30894:data<=-16'd9122;
      30895:data<=-16'd8117;
      30896:data<=-16'd9165;
      30897:data<=-16'd6329;
      30898:data<=16'd534;
      30899:data<=16'd2977;
      30900:data<=16'd1780;
      30901:data<=16'd2171;
      30902:data<=16'd2837;
      30903:data<=16'd2432;
      30904:data<=16'd2634;
      30905:data<=16'd3621;
      30906:data<=16'd4376;
      30907:data<=16'd4799;
      30908:data<=16'd5016;
      30909:data<=16'd4687;
      30910:data<=16'd4117;
      30911:data<=16'd4963;
      30912:data<=16'd7156;
      30913:data<=16'd7685;
      30914:data<=16'd6458;
      30915:data<=16'd5988;
      30916:data<=16'd5844;
      30917:data<=16'd6381;
      30918:data<=16'd8432;
      30919:data<=16'd8928;
      30920:data<=16'd7674;
      30921:data<=16'd7385;
      30922:data<=16'd7459;
      30923:data<=16'd7985;
      30924:data<=16'd9259;
      30925:data<=16'd9426;
      30926:data<=16'd8968;
      30927:data<=16'd8866;
      30928:data<=16'd8520;
      30929:data<=16'd8352;
      30930:data<=16'd8927;
      30931:data<=16'd9928;
      30932:data<=16'd10017;
      30933:data<=16'd8965;
      30934:data<=16'd8617;
      30935:data<=16'd8570;
      30936:data<=16'd8633;
      30937:data<=16'd10202;
      30938:data<=16'd10619;
      30939:data<=16'd9245;
      30940:data<=16'd9283;
      30941:data<=16'd9003;
      30942:data<=16'd8416;
      30943:data<=16'd10398;
      30944:data<=16'd11157;
      30945:data<=16'd10241;
      30946:data<=16'd11251;
      30947:data<=16'd8919;
      30948:data<=16'd2605;
      30949:data<=16'd1287;
      30950:data<=16'd3566;
      30951:data<=16'd3425;
      30952:data<=16'd3086;
      30953:data<=16'd3131;
      30954:data<=16'd2447;
      30955:data<=16'd3362;
      30956:data<=16'd4798;
      30957:data<=16'd4491;
      30958:data<=16'd4225;
      30959:data<=16'd4485;
      30960:data<=16'd4047;
      30961:data<=16'd4068;
      30962:data<=16'd5130;
      30963:data<=16'd5459;
      30964:data<=16'd5162;
      30965:data<=16'd5321;
      30966:data<=16'd5046;
      30967:data<=16'd5084;
      30968:data<=16'd6300;
      30969:data<=16'd6596;
      30970:data<=16'd6311;
      30971:data<=16'd6431;
      30972:data<=16'd5504;
      30973:data<=16'd5124;
      30974:data<=16'd6425;
      30975:data<=16'd7001;
      30976:data<=16'd6821;
      30977:data<=16'd6721;
      30978:data<=16'd6222;
      30979:data<=16'd5809;
      30980:data<=16'd6229;
      30981:data<=16'd7248;
      30982:data<=16'd7332;
      30983:data<=16'd6755;
      30984:data<=16'd6959;
      30985:data<=16'd6505;
      30986:data<=16'd6231;
      30987:data<=16'd7477;
      30988:data<=16'd7294;
      30989:data<=16'd6604;
      30990:data<=16'd6965;
      30991:data<=16'd6169;
      30992:data<=16'd6005;
      30993:data<=16'd7004;
      30994:data<=16'd7054;
      30995:data<=16'd6948;
      30996:data<=16'd5782;
      30997:data<=16'd6173;
      30998:data<=16'd11555;
      30999:data<=16'd14812;
      31000:data<=16'd13113;
      31001:data<=16'd12093;
      31002:data<=16'd11473;
      31003:data<=16'd10707;
      31004:data<=16'd11022;
      31005:data<=16'd9740;
      31006:data<=16'd7194;
      31007:data<=16'd6240;
      31008:data<=16'd6015;
      31009:data<=16'd5474;
      31010:data<=16'd5341;
      31011:data<=16'd4673;
      31012:data<=16'd2702;
      31013:data<=16'd1891;
      31014:data<=16'd2223;
      31015:data<=16'd1466;
      31016:data<=16'd1133;
      31017:data<=16'd587;
      31018:data<=-16'd1539;
      31019:data<=-16'd2030;
      31020:data<=-16'd1850;
      31021:data<=-16'd2746;
      31022:data<=-16'd2162;
      31023:data<=-16'd2038;
      31024:data<=-16'd3868;
      31025:data<=-16'd4945;
      31026:data<=-16'd5310;
      31027:data<=-16'd5209;
      31028:data<=-16'd4733;
      31029:data<=-16'd4998;
      31030:data<=-16'd6040;
      31031:data<=-16'd7662;
      31032:data<=-16'd7821;
      31033:data<=-16'd6725;
      31034:data<=-16'd7338;
      31035:data<=-16'd7768;
      31036:data<=-16'd7888;
      31037:data<=-16'd9436;
      31038:data<=-16'd9288;
      31039:data<=-16'd8442;
      31040:data<=-16'd8972;
      31041:data<=-16'd8664;
      31042:data<=-16'd8804;
      31043:data<=-16'd9612;
      31044:data<=-16'd9782;
      31045:data<=-16'd10281;
      31046:data<=-16'd9330;
      31047:data<=-16'd9206;
      31048:data<=-16'd14001;
      31049:data<=-16'd18701;
      31050:data<=-16'd19714;
      31051:data<=-16'd19155;
      31052:data<=-16'd18243;
      31053:data<=-16'd17910;
      31054:data<=-16'd17431;
      31055:data<=-16'd17065;
      31056:data<=-16'd17916;
      31057:data<=-16'd17541;
      31058:data<=-16'd16430;
      31059:data<=-16'd16371;
      31060:data<=-16'd15481;
      31061:data<=-16'd15018;
      31062:data<=-16'd16172;
      31063:data<=-16'd16167;
      31064:data<=-16'd14992;
      31065:data<=-16'd14219;
      31066:data<=-16'd13652;
      31067:data<=-16'd13315;
      31068:data<=-16'd13755;
      31069:data<=-16'd14280;
      31070:data<=-16'd13474;
      31071:data<=-16'd12718;
      31072:data<=-16'd12892;
      31073:data<=-16'd12041;
      31074:data<=-16'd11623;
      31075:data<=-16'd12560;
      31076:data<=-16'd12225;
      31077:data<=-16'd11740;
      31078:data<=-16'd11611;
      31079:data<=-16'd10167;
      31080:data<=-16'd9729;
      31081:data<=-16'd10557;
      31082:data<=-16'd10510;
      31083:data<=-16'd10379;
      31084:data<=-16'd9687;
      31085:data<=-16'd8305;
      31086:data<=-16'd8223;
      31087:data<=-16'd8966;
      31088:data<=-16'd9544;
      31089:data<=-16'd9608;
      31090:data<=-16'd8683;
      31091:data<=-16'd7691;
      31092:data<=-16'd7138;
      31093:data<=-16'd7571;
      31094:data<=-16'd8887;
      31095:data<=-16'd8461;
      31096:data<=-16'd7527;
      31097:data<=-16'd7808;
      31098:data<=-16'd4303;
      31099:data<=16'd2232;
      31100:data<=16'd4071;
      31101:data<=16'd2684;
      31102:data<=16'd3045;
      31103:data<=16'd3250;
      31104:data<=16'd2846;
      31105:data<=16'd4103;
      31106:data<=16'd5488;
      31107:data<=16'd5486;
      31108:data<=16'd5562;
      31109:data<=16'd5721;
      31110:data<=16'd5222;
      31111:data<=16'd5800;
      31112:data<=16'd7598;
      31113:data<=16'd8202;
      31114:data<=16'd7921;
      31115:data<=16'd7862;
      31116:data<=16'd7403;
      31117:data<=16'd7409;
      31118:data<=16'd8573;
      31119:data<=16'd9450;
      31120:data<=16'd9253;
      31121:data<=16'd8740;
      31122:data<=16'd8731;
      31123:data<=16'd8696;
      31124:data<=16'd8895;
      31125:data<=16'd10302;
      31126:data<=16'd10818;
      31127:data<=16'd10052;
      31128:data<=16'd10202;
      31129:data<=16'd9873;
      31130:data<=16'd9500;
      31131:data<=16'd10787;
      31132:data<=16'd11025;
      31133:data<=16'd10577;
      31134:data<=16'd10998;
      31135:data<=16'd10369;
      31136:data<=16'd9774;
      31137:data<=16'd10358;
      31138:data<=16'd11036;
      31139:data<=16'd11576;
      31140:data<=16'd11145;
      31141:data<=16'd10561;
      31142:data<=16'd10278;
      31143:data<=16'd10166;
      31144:data<=16'd11956;
      31145:data<=16'd12263;
      31146:data<=16'd10792;
      31147:data<=16'd12132;
      31148:data<=16'd9545;
      31149:data<=16'd2399;
      31150:data<=16'd1847;
      31151:data<=16'd4250;
      31152:data<=16'd3817;
      31153:data<=16'd4253;
      31154:data<=16'd3888;
      31155:data<=16'd3228;
      31156:data<=16'd4898;
      31157:data<=16'd5503;
      31158:data<=16'd5247;
      31159:data<=16'd5419;
      31160:data<=16'd4845;
      31161:data<=16'd4719;
      31162:data<=16'd5180;
      31163:data<=16'd5712;
      31164:data<=16'd5946;
      31165:data<=16'd5529;
      31166:data<=16'd5674;
      31167:data<=16'd5335;
      31168:data<=16'd5051;
      31169:data<=16'd6764;
      31170:data<=16'd7203;
      31171:data<=16'd6319;
      31172:data<=16'd6516;
      31173:data<=16'd5973;
      31174:data<=16'd6067;
      31175:data<=16'd7764;
      31176:data<=16'd8105;
      31177:data<=16'd7500;
      31178:data<=16'd6936;
      31179:data<=16'd6461;
      31180:data<=16'd6852;
      31181:data<=16'd7670;
      31182:data<=16'd8281;
      31183:data<=16'd7765;
      31184:data<=16'd6781;
      31185:data<=16'd6795;
      31186:data<=16'd6811;
      31187:data<=16'd7702;
      31188:data<=16'd8872;
      31189:data<=16'd7756;
      31190:data<=16'd7203;
      31191:data<=16'd7194;
      31192:data<=16'd5902;
      31193:data<=16'd6742;
      31194:data<=16'd8059;
      31195:data<=16'd7800;
      31196:data<=16'd7805;
      31197:data<=16'd6206;
      31198:data<=16'd6862;
      31199:data<=16'd12821;
      31200:data<=16'd15644;
      31201:data<=16'd14207;
      31202:data<=16'd13435;
      31203:data<=16'd12090;
      31204:data<=16'd11174;
      31205:data<=16'd11166;
      31206:data<=16'd9539;
      31207:data<=16'd7906;
      31208:data<=16'd7274;
      31209:data<=16'd6584;
      31210:data<=16'd6314;
      31211:data<=16'd6170;
      31212:data<=16'd5169;
      31213:data<=16'd3491;
      31214:data<=16'd2575;
      31215:data<=16'd2579;
      31216:data<=16'd2231;
      31217:data<=16'd1961;
      31218:data<=16'd1116;
      31219:data<=-16'd763;
      31220:data<=-16'd1119;
      31221:data<=-16'd869;
      31222:data<=-16'd1554;
      31223:data<=-16'd1485;
      31224:data<=-16'd2065;
      31225:data<=-16'd3803;
      31226:data<=-16'd4320;
      31227:data<=-16'd4358;
      31228:data<=-16'd4356;
      31229:data<=-16'd4070;
      31230:data<=-16'd4611;
      31231:data<=-16'd5436;
      31232:data<=-16'd6220;
      31233:data<=-16'd6642;
      31234:data<=-16'd6150;
      31235:data<=-16'd6319;
      31236:data<=-16'd6869;
      31237:data<=-16'd7297;
      31238:data<=-16'd8454;
      31239:data<=-16'd8376;
      31240:data<=-16'd7820;
      31241:data<=-16'd8520;
      31242:data<=-16'd7846;
      31243:data<=-16'd7638;
      31244:data<=-16'd9541;
      31245:data<=-16'd9714;
      31246:data<=-16'd9473;
      31247:data<=-16'd9462;
      31248:data<=-16'd8392;
      31249:data<=-16'd12184;
      31250:data<=-16'd19215;
      31251:data<=-16'd20510;
      31252:data<=-16'd18729;
      31253:data<=-16'd18114;
      31254:data<=-16'd16962;
      31255:data<=-16'd16801;
      31256:data<=-16'd17817;
      31257:data<=-16'd17546;
      31258:data<=-16'd16851;
      31259:data<=-16'd16600;
      31260:data<=-16'd16010;
      31261:data<=-16'd15247;
      31262:data<=-16'd15435;
      31263:data<=-16'd16392;
      31264:data<=-16'd16258;
      31265:data<=-16'd15379;
      31266:data<=-16'd14897;
      31267:data<=-16'd13994;
      31268:data<=-16'd13682;
      31269:data<=-16'd14886;
      31270:data<=-16'd15262;
      31271:data<=-16'd14184;
      31272:data<=-16'd13311;
      31273:data<=-16'd12790;
      31274:data<=-16'd12417;
      31275:data<=-16'd12907;
      31276:data<=-16'd13497;
      31277:data<=-16'd12672;
      31278:data<=-16'd11759;
      31279:data<=-16'd11530;
      31280:data<=-16'd10736;
      31281:data<=-16'd11071;
      31282:data<=-16'd12439;
      31283:data<=-16'd11734;
      31284:data<=-16'd10774;
      31285:data<=-16'd10637;
      31286:data<=-16'd9320;
      31287:data<=-16'd9142;
      31288:data<=-16'd10627;
      31289:data<=-16'd10709;
      31290:data<=-16'd9820;
      31291:data<=-16'd8839;
      31292:data<=-16'd8059;
      31293:data<=-16'd8478;
      31294:data<=-16'd9364;
      31295:data<=-16'd9596;
      31296:data<=-16'd8499;
      31297:data<=-16'd7567;
      31298:data<=-16'd8116;
      31299:data<=-16'd5301;
      31300:data<=16'd1215;
      31301:data<=16'd3598;
      31302:data<=16'd2299;
      31303:data<=16'd2470;
      31304:data<=16'd2720;
      31305:data<=16'd2499;
      31306:data<=16'd3516;
      31307:data<=16'd4837;
      31308:data<=16'd5436;
      31309:data<=16'd5521;
      31310:data<=16'd5322;
      31311:data<=16'd4857;
      31312:data<=16'd5195;
      31313:data<=16'd6904;
      31314:data<=16'd7623;
      31315:data<=16'd7263;
      31316:data<=16'd7523;
      31317:data<=16'd6933;
      31318:data<=16'd6667;
      31319:data<=16'd8492;
      31320:data<=16'd9207;
      31321:data<=16'd8793;
      31322:data<=16'd9009;
      31323:data<=16'd8179;
      31324:data<=16'd7658;
      31325:data<=16'd9085;
      31326:data<=16'd10056;
      31327:data<=16'd9849;
      31328:data<=16'd9411;
      31329:data<=16'd8737;
      31330:data<=16'd8113;
      31331:data<=16'd8504;
      31332:data<=16'd9767;
      31333:data<=16'd9962;
      31334:data<=16'd9483;
      31335:data<=16'd9632;
      31336:data<=16'd8846;
      31337:data<=16'd8204;
      31338:data<=16'd9445;
      31339:data<=16'd10158;
      31340:data<=16'd9950;
      31341:data<=16'd9544;
      31342:data<=16'd8546;
      31343:data<=16'd8689;
      31344:data<=16'd9955;
      31345:data<=16'd10492;
      31346:data<=16'd10056;
      31347:data<=16'd9521;
      31348:data<=16'd9823;
      31349:data<=16'd7856;
      31350:data<=16'd2934;
      31351:data<=16'd1336;
      31352:data<=16'd2306;
      31353:data<=16'd1786;
      31354:data<=16'd2002;
      31355:data<=16'd2083;
      31356:data<=16'd1806;
      31357:data<=16'd3475;
      31358:data<=16'd3803;
      31359:data<=16'd3011;
      31360:data<=16'd3741;
      31361:data<=16'd3377;
      31362:data<=16'd3001;
      31363:data<=16'd4432;
      31364:data<=16'd4884;
      31365:data<=16'd4291;
      31366:data<=16'd3962;
      31367:data<=16'd3767;
      31368:data<=16'd4008;
      31369:data<=16'd4916;
      31370:data<=16'd5818;
      31371:data<=16'd5301;
      31372:data<=16'd4666;
      31373:data<=16'd5301;
      31374:data<=16'd5136;
      31375:data<=16'd5187;
      31376:data<=16'd6385;
      31377:data<=16'd6129;
      31378:data<=16'd5786;
      31379:data<=16'd5941;
      31380:data<=16'd5075;
      31381:data<=16'd5717;
      31382:data<=16'd7347;
      31383:data<=16'd7269;
      31384:data<=16'd6639;
      31385:data<=16'd5805;
      31386:data<=16'd5303;
      31387:data<=16'd6346;
      31388:data<=16'd7392;
      31389:data<=16'd7450;
      31390:data<=16'd7106;
      31391:data<=16'd6751;
      31392:data<=16'd6355;
      31393:data<=16'd6296;
      31394:data<=16'd7410;
      31395:data<=16'd7911;
      31396:data<=16'd7136;
      31397:data<=16'd7083;
      31398:data<=16'd6211;
      31399:data<=16'd5764;
      31400:data<=16'd9882;
      31401:data<=16'd14090;
      31402:data<=16'd13964;
      31403:data<=16'd12502;
      31404:data<=16'd11597;
      31405:data<=16'd11312;
      31406:data<=16'd10619;
      31407:data<=16'd8457;
      31408:data<=16'd6977;
      31409:data<=16'd6485;
      31410:data<=16'd5839;
      31411:data<=16'd5993;
      31412:data<=16'd5556;
      31413:data<=16'd3462;
      31414:data<=16'd2161;
      31415:data<=16'd2076;
      31416:data<=16'd2090;
      31417:data<=16'd2202;
      31418:data<=16'd1657;
      31419:data<=16'd152;
      31420:data<=-16'd980;
      31421:data<=-16'd1231;
      31422:data<=-16'd1545;
      31423:data<=-16'd2005;
      31424:data<=-16'd2108;
      31425:data<=-16'd2729;
      31426:data<=-16'd3982;
      31427:data<=-16'd4637;
      31428:data<=-16'd4989;
      31429:data<=-16'd4930;
      31430:data<=-16'd4082;
      31431:data<=-16'd4670;
      31432:data<=-16'd6628;
      31433:data<=-16'd7275;
      31434:data<=-16'd7188;
      31435:data<=-16'd7036;
      31436:data<=-16'd6498;
      31437:data<=-16'd7122;
      31438:data<=-16'd8428;
      31439:data<=-16'd8837;
      31440:data<=-16'd8922;
      31441:data<=-16'd8790;
      31442:data<=-16'd8461;
      31443:data<=-16'd8419;
      31444:data<=-16'd9133;
      31445:data<=-16'd10302;
      31446:data<=-16'd10146;
      31447:data<=-16'd10087;
      31448:data<=-16'd10346;
      31449:data<=-16'd8338;
      31450:data<=-16'd10887;
      31451:data<=-16'd19420;
      31452:data<=-16'd21265;
      31453:data<=-16'd18193;
      31454:data<=-16'd18600;
      31455:data<=-16'd17928;
      31456:data<=-16'd17009;
      31457:data<=-16'd18653;
      31458:data<=-16'd18409;
      31459:data<=-16'd17582;
      31460:data<=-16'd17308;
      31461:data<=-16'd15863;
      31462:data<=-16'd15750;
      31463:data<=-16'd16675;
      31464:data<=-16'd16772;
      31465:data<=-16'd16130;
      31466:data<=-16'd15064;
      31467:data<=-16'd15039;
      31468:data<=-16'd14892;
      31469:data<=-16'd14551;
      31470:data<=-16'd15679;
      31471:data<=-16'd15268;
      31472:data<=-16'd13957;
      31473:data<=-16'd13979;
      31474:data<=-16'd12747;
      31475:data<=-16'd12437;
      31476:data<=-16'd14152;
      31477:data<=-16'd13879;
      31478:data<=-16'd12871;
      31479:data<=-16'd12405;
      31480:data<=-16'd11473;
      31481:data<=-16'd11515;
      31482:data<=-16'd12323;
      31483:data<=-16'd12475;
      31484:data<=-16'd11688;
      31485:data<=-16'd10727;
      31486:data<=-16'd10305;
      31487:data<=-16'd9929;
      31488:data<=-16'd10426;
      31489:data<=-16'd10810;
      31490:data<=-16'd9580;
      31491:data<=-16'd9339;
      31492:data<=-16'd9171;
      31493:data<=-16'd8113;
      31494:data<=-16'd9075;
      31495:data<=-16'd9820;
      31496:data<=-16'd9078;
      31497:data<=-16'd8366;
      31498:data<=-16'd7465;
      31499:data<=-16'd8144;
      31500:data<=-16'd6061;
      31501:data<=16'd1081;
      31502:data<=16'd3645;
      31503:data<=16'd2453;
      31504:data<=16'd3480;
      31505:data<=16'd3025;
      31506:data<=16'd3112;
      31507:data<=16'd5453;
      31508:data<=16'd5768;
      31509:data<=16'd5937;
      31510:data<=16'd6279;
      31511:data<=16'd5307;
      31512:data<=16'd5883;
      31513:data<=16'd7403;
      31514:data<=16'd8046;
      31515:data<=16'd8137;
      31516:data<=16'd7938;
      31517:data<=16'd7988;
      31518:data<=16'd7594;
      31519:data<=16'd7917;
      31520:data<=16'd9667;
      31521:data<=16'd9837;
      31522:data<=16'd9444;
      31523:data<=16'd9608;
      31524:data<=16'd8507;
      31525:data<=16'd8736;
      31526:data<=16'd10662;
      31527:data<=16'd10915;
      31528:data<=16'd10519;
      31529:data<=16'd10478;
      31530:data<=16'd9931;
      31531:data<=16'd9838;
      31532:data<=16'd10824;
      31533:data<=16'd11656;
      31534:data<=16'd11439;
      31535:data<=16'd11144;
      31536:data<=16'd10701;
      31537:data<=16'd9696;
      31538:data<=16'd10290;
      31539:data<=16'd11570;
      31540:data<=16'd11109;
      31541:data<=16'd10768;
      31542:data<=16'd10560;
      31543:data<=16'd9677;
      31544:data<=16'd10387;
      31545:data<=16'd11717;
      31546:data<=16'd11753;
      31547:data<=16'd11456;
      31548:data<=16'd10934;
      31549:data<=16'd10684;
      31550:data<=16'd10199;
      31551:data<=16'd7040;
      31552:data<=16'd3677;
      31553:data<=16'd3424;
      31554:data<=16'd3592;
      31555:data<=16'd2964;
      31556:data<=16'd3657;
      31557:data<=16'd4896;
      31558:data<=16'd5354;
      31559:data<=16'd5209;
      31560:data<=16'd4798;
      31561:data<=16'd4769;
      31562:data<=16'd4522;
      31563:data<=16'd4636;
      31564:data<=16'd6379;
      31565:data<=16'd6752;
      31566:data<=16'd5542;
      31567:data<=16'd5791;
      31568:data<=16'd5674;
      31569:data<=16'd5658;
      31570:data<=16'd7447;
      31571:data<=16'd7433;
      31572:data<=16'd6414;
      31573:data<=16'd6754;
      31574:data<=16'd6337;
      31575:data<=16'd6560;
      31576:data<=16'd7940;
      31577:data<=16'd7850;
      31578:data<=16'd7580;
      31579:data<=16'd7706;
      31580:data<=16'd7121;
      31581:data<=16'd7059;
      31582:data<=16'd7903;
      31583:data<=16'd8376;
      31584:data<=16'd7893;
      31585:data<=16'd7470;
      31586:data<=16'd7424;
      31587:data<=16'd7101;
      31588:data<=16'd7838;
      31589:data<=16'd8857;
      31590:data<=16'd8137;
      31591:data<=16'd7783;
      31592:data<=16'd8043;
      31593:data<=16'd7410;
      31594:data<=16'd7602;
      31595:data<=16'd8802;
      31596:data<=16'd8886;
      31597:data<=16'd7626;
      31598:data<=16'd7471;
      31599:data<=16'd8096;
      31600:data<=16'd6652;
      31601:data<=16'd8020;
      31602:data<=16'd13954;
      31603:data<=16'd15164;
      31604:data<=16'd12756;
      31605:data<=16'd13110;
      31606:data<=16'd12275;
      31607:data<=16'd9903;
      31608:data<=16'd8939;
      31609:data<=16'd8069;
      31610:data<=16'd7562;
      31611:data<=16'd7374;
      31612:data<=16'd7115;
      31613:data<=16'd6222;
      31614:data<=16'd3659;
      31615:data<=16'd2475;
      31616:data<=16'd2737;
      31617:data<=16'd2350;
      31618:data<=16'd3049;
      31619:data<=16'd2258;
      31620:data<=-16'd517;
      31621:data<=-16'd578;
      31622:data<=-16'd149;
      31623:data<=-16'd811;
      31624:data<=-16'd479;
      31625:data<=-16'd1107;
      31626:data<=-16'd2711;
      31627:data<=-16'd3450;
      31628:data<=-16'd3618;
      31629:data<=-16'd3562;
      31630:data<=-16'd3651;
      31631:data<=-16'd3644;
      31632:data<=-16'd4472;
      31633:data<=-16'd6206;
      31634:data<=-16'd6275;
      31635:data<=-16'd5923;
      31636:data<=-16'd5991;
      31637:data<=-16'd5206;
      31638:data<=-16'd6264;
      31639:data<=-16'd8290;
      31640:data<=-16'd8100;
      31641:data<=-16'd7705;
      31642:data<=-16'd7617;
      31643:data<=-16'd7188;
      31644:data<=-16'd7692;
      31645:data<=-16'd9019;
      31646:data<=-16'd9737;
      31647:data<=-16'd8711;
      31648:data<=-16'd8251;
      31649:data<=-16'd8971;
      31650:data<=-16'd8210;
      31651:data<=-16'd10798;
      31652:data<=-16'd17656;
      31653:data<=-16'd19458;
      31654:data<=-16'd17437;
      31655:data<=-16'd17142;
      31656:data<=-16'd16401;
      31657:data<=-16'd16478;
      31658:data<=-16'd17863;
      31659:data<=-16'd17233;
      31660:data<=-16'd16337;
      31661:data<=-16'd16092;
      31662:data<=-16'd15095;
      31663:data<=-16'd15197;
      31664:data<=-16'd16151;
      31665:data<=-16'd15503;
      31666:data<=-16'd14472;
      31667:data<=-16'd14413;
      31668:data<=-16'd13964;
      31669:data<=-16'd13744;
      31670:data<=-16'd14697;
      31671:data<=-16'd14671;
      31672:data<=-16'd13835;
      31673:data<=-16'd13590;
      31674:data<=-16'd12672;
      31675:data<=-16'd12099;
      31676:data<=-16'd13024;
      31677:data<=-16'd13362;
      31678:data<=-16'd12633;
      31679:data<=-16'd11728;
      31680:data<=-16'd11156;
      31681:data<=-16'd11065;
      31682:data<=-16'd11116;
      31683:data<=-16'd11599;
      31684:data<=-16'd11341;
      31685:data<=-16'd10125;
      31686:data<=-16'd10016;
      31687:data<=-16'd9797;
      31688:data<=-16'd9373;
      31689:data<=-16'd10220;
      31690:data<=-16'd9882;
      31691:data<=-16'd9013;
      31692:data<=-16'd9012;
      31693:data<=-16'd7779;
      31694:data<=-16'd7653;
      31695:data<=-16'd8934;
      31696:data<=-16'd8214;
      31697:data<=-16'd7712;
      31698:data<=-16'd7609;
      31699:data<=-16'd6481;
      31700:data<=-16'd6871;
      31701:data<=-16'd5383;
      31702:data<=16'd566;
      31703:data<=16'd4135;
      31704:data<=16'd3623;
      31705:data<=16'd3318;
      31706:data<=16'd3336;
      31707:data<=16'd3953;
      31708:data<=16'd5858;
      31709:data<=16'd6667;
      31710:data<=16'd6285;
      31711:data<=16'd6006;
      31712:data<=16'd5374;
      31713:data<=16'd6020;
      31714:data<=16'd7982;
      31715:data<=16'd8155;
      31716:data<=16'd7706;
      31717:data<=16'd7855;
      31718:data<=16'd7059;
      31719:data<=16'd7448;
      31720:data<=16'd9438;
      31721:data<=16'd9829;
      31722:data<=16'd9362;
      31723:data<=16'd9373;
      31724:data<=16'd9065;
      31725:data<=16'd8859;
      31726:data<=16'd9541;
      31727:data<=16'd10751;
      31728:data<=16'd10777;
      31729:data<=16'd9571;
      31730:data<=16'd9125;
      31731:data<=16'd9148;
      31732:data<=16'd9730;
      31733:data<=16'd11194;
      31734:data<=16'd11075;
      31735:data<=16'd10075;
      31736:data<=16'd10093;
      31737:data<=16'd9726;
      31738:data<=16'd9870;
      31739:data<=16'd11132;
      31740:data<=16'd11159;
      31741:data<=16'd10557;
      31742:data<=16'd10311;
      31743:data<=16'd9517;
      31744:data<=16'd9555;
      31745:data<=16'd10903;
      31746:data<=16'd10950;
      31747:data<=16'd10181;
      31748:data<=16'd10490;
      31749:data<=16'd9741;
      31750:data<=16'd8872;
      31751:data<=16'd10408;
      31752:data<=16'd8519;
      31753:data<=16'd2535;
      31754:data<=16'd1198;
      31755:data<=16'd2500;
      31756:data<=16'd1516;
      31757:data<=16'd2575;
      31758:data<=16'd4479;
      31759:data<=16'd3577;
      31760:data<=16'd3307;
      31761:data<=16'd3958;
      31762:data<=16'd3557;
      31763:data<=16'd3832;
      31764:data<=16'd4807;
      31765:data<=16'd5153;
      31766:data<=16'd5222;
      31767:data<=16'd5071;
      31768:data<=16'd4491;
      31769:data<=16'd4464;
      31770:data<=16'd5691;
      31771:data<=16'd6543;
      31772:data<=16'd5850;
      31773:data<=16'd5194;
      31774:data<=16'd5175;
      31775:data<=16'd4969;
      31776:data<=16'd5357;
      31777:data<=16'd6514;
      31778:data<=16'd6777;
      31779:data<=16'd6297;
      31780:data<=16'd6235;
      31781:data<=16'd5915;
      31782:data<=16'd5846;
      31783:data<=16'd6843;
      31784:data<=16'd6989;
      31785:data<=16'd6476;
      31786:data<=16'd6438;
      31787:data<=16'd5695;
      31788:data<=16'd5988;
      31789:data<=16'd7591;
      31790:data<=16'd7232;
      31791:data<=16'd6695;
      31792:data<=16'd6905;
      31793:data<=16'd5726;
      31794:data<=16'd5532;
      31795:data<=16'd6626;
      31796:data<=16'd6886;
      31797:data<=16'd6866;
      31798:data<=16'd6028;
      31799:data<=16'd5791;
      31800:data<=16'd6454;
      31801:data<=16'd5031;
      31802:data<=16'd6393;
      31803:data<=16'd12091;
      31804:data<=16'd13356;
      31805:data<=16'd11417;
      31806:data<=16'd11658;
      31807:data<=16'd10387;
      31808:data<=16'd7688;
      31809:data<=16'd6963;
      31810:data<=16'd6686;
      31811:data<=16'd6172;
      31812:data<=16'd5962;
      31813:data<=16'd4939;
      31814:data<=16'd3057;
      31815:data<=16'd1965;
      31816:data<=16'd1991;
      31817:data<=16'd1653;
      31818:data<=16'd1257;
      31819:data<=16'd1168;
      31820:data<=-16'd364;
      31821:data<=-16'd2020;
      31822:data<=-16'd1911;
      31823:data<=-16'd1942;
      31824:data<=-16'd2243;
      31825:data<=-16'd1977;
      31826:data<=-16'd2884;
      31827:data<=-16'd4510;
      31828:data<=-16'd4861;
      31829:data<=-16'd4731;
      31830:data<=-16'd4874;
      31831:data<=-16'd4698;
      31832:data<=-16'd5257;
      31833:data<=-16'd6836;
      31834:data<=-16'd7165;
      31835:data<=-16'd6783;
      31836:data<=-16'd7300;
      31837:data<=-16'd7094;
      31838:data<=-16'd6752;
      31839:data<=-16'd7853;
      31840:data<=-16'd8523;
      31841:data<=-16'd8495;
      31842:data<=-16'd8481;
      31843:data<=-16'd7941;
      31844:data<=-16'd7837;
      31845:data<=-16'd8583;
      31846:data<=-16'd9630;
      31847:data<=-16'd10044;
      31848:data<=-16'd9206;
      31849:data<=-16'd9315;
      31850:data<=-16'd9682;
      31851:data<=-16'd9254;
      31852:data<=-16'd12886;
      31853:data<=-16'd18660;
      31854:data<=-16'd19792;
      31855:data<=-16'd18636;
      31856:data<=-16'd18130;
      31857:data<=-16'd17887;
      31858:data<=-16'd18548;
      31859:data<=-16'd18569;
      31860:data<=-16'd17898;
      31861:data<=-16'd17531;
      31862:data<=-16'd16345;
      31863:data<=-16'd15922;
      31864:data<=-16'd16815;
      31865:data<=-16'd16876;
      31866:data<=-16'd16493;
      31867:data<=-16'd16031;
      31868:data<=-16'd15273;
      31869:data<=-16'd14731;
      31870:data<=-16'd14901;
      31871:data<=-16'd15937;
      31872:data<=-16'd15779;
      31873:data<=-16'd14577;
      31874:data<=-16'd14389;
      31875:data<=-16'd13635;
      31876:data<=-16'd13292;
      31877:data<=-16'd14654;
      31878:data<=-16'd14521;
      31879:data<=-16'd13764;
      31880:data<=-16'd13458;
      31881:data<=-16'd12157;
      31882:data<=-16'd12316;
      31883:data<=-16'd13494;
      31884:data<=-16'd13294;
      31885:data<=-16'd12959;
      31886:data<=-16'd12008;
      31887:data<=-16'd10854;
      31888:data<=-16'd11204;
      31889:data<=-16'd11822;
      31890:data<=-16'd11999;
      31891:data<=-16'd11562;
      31892:data<=-16'd11004;
      31893:data<=-16'd10621;
      31894:data<=-16'd9274;
      31895:data<=-16'd9435;
      31896:data<=-16'd10959;
      31897:data<=-16'd10169;
      31898:data<=-16'd9550;
      31899:data<=-16'd9301;
      31900:data<=-16'd7746;
      31901:data<=-16'd7987;
      31902:data<=-16'd6279;
      31903:data<=-16'd217;
      31904:data<=16'd2804;
      31905:data<=16'd2499;
      31906:data<=16'd2798;
      31907:data<=16'd3075;
      31908:data<=16'd4011;
      31909:data<=16'd4925;
      31910:data<=16'd4767;
      31911:data<=16'd5054;
      31912:data<=16'd5046;
      31913:data<=16'd4780;
      31914:data<=16'd5821;
      31915:data<=16'd6740;
      31916:data<=16'd6602;
      31917:data<=16'd6584;
      31918:data<=16'd6702;
      31919:data<=16'd6583;
      31920:data<=16'd7251;
      31921:data<=16'd8499;
      31922:data<=16'd8526;
      31923:data<=16'd8237;
      31924:data<=16'd8454;
      31925:data<=16'd8044;
      31926:data<=16'd8408;
      31927:data<=16'd9526;
      31928:data<=16'd9498;
      31929:data<=16'd9706;
      31930:data<=16'd9967;
      31931:data<=16'd9213;
      31932:data<=16'd9312;
      31933:data<=16'd10208;
      31934:data<=16'd10871;
      31935:data<=16'd10934;
      31936:data<=16'd10102;
      31937:data<=16'd9876;
      31938:data<=16'd9999;
      31939:data<=16'd9944;
      31940:data<=16'd10950;
      31941:data<=16'd11159;
      31942:data<=16'd10452;
      31943:data<=16'd10596;
      31944:data<=16'd9984;
      31945:data<=16'd10082;
      31946:data<=16'd11496;
      31947:data<=16'd10857;
      31948:data<=16'd10470;
      31949:data<=16'd10904;
      31950:data<=16'd9464;
      31951:data<=16'd9997;
      31952:data<=16'd10945;
      31953:data<=16'd6661;
      31954:data<=16'd2675;
      31955:data<=16'd2593;
      31956:data<=16'd2103;
      31957:data<=16'd1992;
      31958:data<=16'd3761;
      31959:data<=16'd4552;
      31960:data<=16'd4073;
      31961:data<=16'd4264;
      31962:data<=16'd4678;
      31963:data<=16'd4211;
      31964:data<=16'd4579;
      31965:data<=16'd6173;
      31966:data<=16'd6238;
      31967:data<=16'd5902;
      31968:data<=16'd6448;
      31969:data<=16'd5495;
      31970:data<=16'd5291;
      31971:data<=16'd7232;
      31972:data<=16'd7298;
      31973:data<=16'd6622;
      31974:data<=16'd6931;
      31975:data<=16'd6064;
      31976:data<=16'd6018;
      31977:data<=16'd7617;
      31978:data<=16'd8011;
      31979:data<=16'd7752;
      31980:data<=16'd7518;
      31981:data<=16'd6795;
      31982:data<=16'd6581;
      31983:data<=16'd7178;
      31984:data<=16'd7826;
      31985:data<=16'd7821;
      31986:data<=16'd7714;
      31987:data<=16'd7793;
      31988:data<=16'd7003;
      31989:data<=16'd7068;
      31990:data<=16'd8578;
      31991:data<=16'd8624;
      31992:data<=16'd7987;
      31993:data<=16'd7585;
      31994:data<=16'd6499;
      31995:data<=16'd6761;
      31996:data<=16'd8067;
      31997:data<=16'd8370;
      31998:data<=16'd8076;
      31999:data<=16'd7224;
      32000:data<=16'd6898;
      32001:data<=16'd7019;
      32002:data<=16'd6910;
      32003:data<=16'd9891;
      32004:data<=16'd13843;
      32005:data<=16'd13602;
      32006:data<=16'd12657;
      32007:data<=16'd12833;
      32008:data<=16'd11144;
      32009:data<=16'd9286;
      32010:data<=16'd8746;
      32011:data<=16'd7940;
      32012:data<=16'd7059;
      32013:data<=16'd6645;
      32014:data<=16'd5615;
      32015:data<=16'd3936;
      32016:data<=16'd3245;
      32017:data<=16'd2878;
      32018:data<=16'd1947;
      32019:data<=16'd2115;
      32020:data<=16'd1924;
      32021:data<=16'd50;
      32022:data<=-16'd678;
      32023:data<=-16'd651;
      32024:data<=-16'd1063;
      32025:data<=-16'd716;
      32026:data<=-16'd922;
      32027:data<=-16'd2231;
      32028:data<=-16'd3245;
      32029:data<=-16'd3824;
      32030:data<=-16'd3891;
      32031:data<=-16'd3723;
      32032:data<=-16'd3545;
      32033:data<=-16'd4027;
      32034:data<=-16'd5394;
      32035:data<=-16'd5441;
      32036:data<=-16'd5401;
      32037:data<=-16'd6558;
      32038:data<=-16'd5864;
      32039:data<=-16'd5588;
      32040:data<=-16'd7418;
      32041:data<=-16'd7500;
      32042:data<=-16'd7441;
      32043:data<=-16'd7928;
      32044:data<=-16'd6754;
      32045:data<=-16'd6959;
      32046:data<=-16'd8307;
      32047:data<=-16'd8584;
      32048:data<=-16'd9065;
      32049:data<=-16'd8630;
      32050:data<=-16'd7905;
      32051:data<=-16'd8243;
      32052:data<=-16'd8668;
      32053:data<=-16'd11708;
      32054:data<=-16'd15872;
      32055:data<=-16'd16431;
      32056:data<=-16'd15719;
      32057:data<=-16'd15267;
      32058:data<=-16'd14922;
      32059:data<=-16'd15925;
      32060:data<=-16'd15869;
      32061:data<=-16'd15095;
      32062:data<=-16'd15194;
      32063:data<=-16'd13673;
      32064:data<=-16'd12872;
      32065:data<=-16'd14574;
      32066:data<=-16'd14640;
      32067:data<=-16'd13620;
      32068:data<=-16'd13241;
      32069:data<=-16'd12176;
      32070:data<=-16'd11949;
      32071:data<=-16'd13103;
      32072:data<=-16'd13549;
      32073:data<=-16'd13212;
      32074:data<=-16'd12678;
      32075:data<=-16'd11856;
      32076:data<=-16'd11341;
      32077:data<=-16'd12005;
      32078:data<=-16'd12842;
      32079:data<=-16'd12392;
      32080:data<=-16'd11844;
      32081:data<=-16'd11383;
      32082:data<=-16'd10038;
      32083:data<=-16'd10076;
      32084:data<=-16'd11788;
      32085:data<=-16'd12158;
      32086:data<=-16'd11197;
      32087:data<=-16'd9999;
      32088:data<=-16'd8995;
      32089:data<=-16'd9371;
      32090:data<=-16'd10311;
      32091:data<=-16'd10151;
      32092:data<=-16'd9439;
      32093:data<=-16'd8821;
      32094:data<=-16'd8114;
      32095:data<=-16'd8167;
      32096:data<=-16'd9251;
      32097:data<=-16'd9320;
      32098:data<=-16'd8410;
      32099:data<=-16'd8199;
      32100:data<=-16'd7232;
      32101:data<=-16'd6255;
      32102:data<=-16'd6836;
      32103:data<=-16'd4566;
      32104:data<=16'd179;
      32105:data<=16'd1668;
      32106:data<=16'd1535;
      32107:data<=16'd2176;
      32108:data<=16'd2604;
      32109:data<=16'd3656;
      32110:data<=16'd4396;
      32111:data<=16'd4399;
      32112:data<=16'd4808;
      32113:data<=16'd4246;
      32114:data<=16'd4126;
      32115:data<=16'd5882;
      32116:data<=16'd6569;
      32117:data<=16'd6376;
      32118:data<=16'd6516;
      32119:data<=16'd6034;
      32120:data<=16'd6169;
      32121:data<=16'd7338;
      32122:data<=16'd8084;
      32123:data<=16'd8264;
      32124:data<=16'd8287;
      32125:data<=16'd8208;
      32126:data<=16'd7855;
      32127:data<=16'd8381;
      32128:data<=16'd9806;
      32129:data<=16'd9735;
      32130:data<=16'd9359;
      32131:data<=16'd9552;
      32132:data<=16'd8420;
      32133:data<=16'd8640;
      32134:data<=16'd10683;
      32135:data<=16'd10871;
      32136:data<=16'd10583;
      32137:data<=16'd10422;
      32138:data<=16'd9218;
      32139:data<=16'd9320;
      32140:data<=16'd10487;
      32141:data<=16'd10781;
      32142:data<=16'd10551;
      32143:data<=16'd10006;
      32144:data<=16'd9582;
      32145:data<=16'd9697;
      32146:data<=16'd10689;
      32147:data<=16'd11579;
      32148:data<=16'd10646;
      32149:data<=16'd10075;
      32150:data<=16'd9976;
      32151:data<=16'd8763;
      32152:data<=16'd9831;
      32153:data<=16'd10340;
      32154:data<=16'd6162;
      32155:data<=16'd4073;
      32156:data<=16'd4649;
      32157:data<=16'd3224;
      32158:data<=16'd3774;
      32159:data<=16'd6187;
      32160:data<=16'd6128;
      32161:data<=16'd5412;
      32162:data<=16'd5100;
      32163:data<=16'd4614;
      32164:data<=16'd5269;
      32165:data<=16'd6949;
      32166:data<=16'd7717;
      32167:data<=16'd6774;
      32168:data<=16'd6155;
      32169:data<=16'd6297;
      32170:data<=16'd5677;
      32171:data<=16'd6216;
      32172:data<=16'd7834;
      32173:data<=16'd7558;
      32174:data<=16'd6816;
      32175:data<=16'd6384;
      32176:data<=16'd5298;
      32177:data<=16'd5868;
      32178:data<=16'd7752;
      32179:data<=16'd7824;
      32180:data<=16'd6984;
      32181:data<=16'd6764;
      32182:data<=16'd6328;
      32183:data<=16'd6481;
      32184:data<=16'd7926;
      32185:data<=16'd8081;
      32186:data<=16'd6898;
      32187:data<=16'd6863;
      32188:data<=16'd6796;
      32189:data<=16'd6602;
      32190:data<=16'd7826;
      32191:data<=16'd8345;
      32192:data<=16'd7838;
      32193:data<=16'd7529;
      32194:data<=16'd6466;
      32195:data<=16'd5912;
      32196:data<=16'd6590;
      32197:data<=16'd7215;
      32198:data<=16'd7667;
      32199:data<=16'd6974;
      32200:data<=16'd6091;
      32201:data<=16'd6138;
      32202:data<=16'd5265;
      32203:data<=16'd6270;
      32204:data<=16'd10234;
      32205:data<=16'd11194;
      32206:data<=16'd9911;
      32207:data<=16'd10254;
      32208:data<=16'd9526;
      32209:data<=16'd7215;
      32210:data<=16'd6068;
      32211:data<=16'd5703;
      32212:data<=16'd5009;
      32213:data<=16'd4613;
      32214:data<=16'd4264;
      32215:data<=16'd2408;
      32216:data<=16'd723;
      32217:data<=16'd1045;
      32218:data<=16'd581;
      32219:data<=-16'd415;
      32220:data<=16'd187;
      32221:data<=-16'd576;
      32222:data<=-16'd2543;
      32223:data<=-16'd2695;
      32224:data<=-16'd2875;
      32225:data<=-16'd3274;
      32226:data<=-16'd2397;
      32227:data<=-16'd2895;
      32228:data<=-16'd4930;
      32229:data<=-16'd5479;
      32230:data<=-16'd5341;
      32231:data<=-16'd5639;
      32232:data<=-16'd5171;
      32233:data<=-16'd5292;
      32234:data<=-16'd7095;
      32235:data<=-16'd7914;
      32236:data<=-16'd7374;
      32237:data<=-16'd7341;
      32238:data<=-16'd7282;
      32239:data<=-16'd7301;
      32240:data<=-16'd8352;
      32241:data<=-16'd9359;
      32242:data<=-16'd9564;
      32243:data<=-16'd9454;
      32244:data<=-16'd9128;
      32245:data<=-16'd8511;
      32246:data<=-16'd8704;
      32247:data<=-16'd10398;
      32248:data<=-16'd11124;
      32249:data<=-16'd10119;
      32250:data<=-16'd9908;
      32251:data<=-16'd9703;
      32252:data<=-16'd9414;
      32253:data<=-16'd12342;
      32254:data<=-16'd16568;
      32255:data<=-16'd17954;
      32256:data<=-16'd17182;
      32257:data<=-16'd16342;
      32258:data<=-16'd16645;
      32259:data<=-16'd17608;
      32260:data<=-16'd17438;
      32261:data<=-16'd16413;
      32262:data<=-16'd15807;
      32263:data<=-16'd15547;
      32264:data<=-16'd15270;
      32265:data<=-16'd15465;
      32266:data<=-16'd16022;
      32267:data<=-16'd15421;
      32268:data<=-16'd14351;
      32269:data<=-16'd14217;
      32270:data<=-16'd13584;
      32271:data<=-16'd13261;
      32272:data<=-16'd14642;
      32273:data<=-16'd14833;
      32274:data<=-16'd13693;
      32275:data<=-16'd13409;
      32276:data<=-16'd12948;
      32277:data<=-16'd12912;
      32278:data<=-16'd14210;
      32279:data<=-16'd14216;
      32280:data<=-16'd12784;
      32281:data<=-16'd12047;
      32282:data<=-16'd11670;
      32283:data<=-16'd11562;
      32284:data<=-16'd12427;
      32285:data<=-16'd12825;
      32286:data<=-16'd11882;
      32287:data<=-16'd11142;
      32288:data<=-16'd10722;
      32289:data<=-16'd9868;
      32290:data<=-16'd10058;
      32291:data<=-16'd11127;
      32292:data<=-16'd10787;
      32293:data<=-16'd9812;
      32294:data<=-16'd9433;
      32295:data<=-16'd8909;
      32296:data<=-16'd9145;
      32297:data<=-16'd10060;
      32298:data<=-16'd9508;
      32299:data<=-16'd8552;
      32300:data<=-16'd8369;
      32301:data<=-16'd7934;
      32302:data<=-16'd7908;
      32303:data<=-16'd6672;
      32304:data<=-16'd2097;
      32305:data<=16'd1174;
      32306:data<=16'd822;
      32307:data<=16'd682;
      32308:data<=16'd1518;
      32309:data<=16'd2717;
      32310:data<=16'd3847;
      32311:data<=16'd3501;
      32312:data<=16'd3444;
      32313:data<=16'd3958;
      32314:data<=16'd3327;
      32315:data<=16'd3973;
      32316:data<=16'd5647;
      32317:data<=16'd5624;
      32318:data<=16'd5683;
      32319:data<=16'd5952;
      32320:data<=16'd5238;
      32321:data<=16'd5732;
      32322:data<=16'd7272;
      32323:data<=16'd7741;
      32324:data<=16'd7571;
      32325:data<=16'd7392;
      32326:data<=16'd7175;
      32327:data<=16'd7686;
      32328:data<=16'd9089;
      32329:data<=16'd9770;
      32330:data<=16'd9203;
      32331:data<=16'd8790;
      32332:data<=16'd8470;
      32333:data<=16'd8147;
      32334:data<=16'd8960;
      32335:data<=16'd9915;
      32336:data<=16'd9849;
      32337:data<=16'd9726;
      32338:data<=16'd9542;
      32339:data<=16'd8693;
      32340:data<=16'd8698;
      32341:data<=16'd10295;
      32342:data<=16'd10887;
      32343:data<=16'd10052;
      32344:data<=16'd9914;
      32345:data<=16'd9480;
      32346:data<=16'd9285;
      32347:data<=16'd10828;
      32348:data<=16'd10871;
      32349:data<=16'd9871;
      32350:data<=16'd10144;
      32351:data<=16'd9362;
      32352:data<=16'd9629;
      32353:data<=16'd11215;
      32354:data<=16'd8207;
      32355:data<=16'd4038;
      32356:data<=16'd4018;
      32357:data<=16'd4187;
      32358:data<=16'd3354;
      32359:data<=16'd4167;
      32360:data<=16'd5647;
      32361:data<=16'd5809;
      32362:data<=16'd5369;
      32363:data<=16'd5510;
      32364:data<=16'd4998;
      32365:data<=16'd4999;
      32366:data<=16'd7066;
      32367:data<=16'd7365;
      32368:data<=16'd6243;
      32369:data<=16'd6728;
      32370:data<=16'd6266;
      32371:data<=16'd5999;
      32372:data<=16'd7774;
      32373:data<=16'd7844;
      32374:data<=16'd6948;
      32375:data<=16'd7154;
      32376:data<=16'd6702;
      32377:data<=16'd6275;
      32378:data<=16'd6910;
      32379:data<=16'd7532;
      32380:data<=16'd7451;
      32381:data<=16'd7048;
      32382:data<=16'd6892;
      32383:data<=16'd6458;
      32384:data<=16'd6813;
      32385:data<=16'd8240;
      32386:data<=16'd7902;
      32387:data<=16'd7090;
      32388:data<=16'd7283;
      32389:data<=16'd6596;
      32390:data<=16'd7124;
      32391:data<=16'd8580;
      32392:data<=16'd7746;
      32393:data<=16'd7183;
      32394:data<=16'd7500;
      32395:data<=16'd6871;
      32396:data<=16'd7018;
      32397:data<=16'd7492;
      32398:data<=16'd7338;
      32399:data<=16'd7319;
      32400:data<=16'd6933;
      32401:data<=16'd6819;
      32402:data<=16'd6426;
      32403:data<=16'd5354;
      32404:data<=16'd7467;
      32405:data<=16'd11371;
      32406:data<=16'd11621;
      32407:data<=16'd10608;
      32408:data<=16'd11069;
      32409:data<=16'd9794;
      32410:data<=16'd7330;
      32411:data<=16'd6717;
      32412:data<=16'd6340;
      32413:data<=16'd5633;
      32414:data<=16'd5932;
      32415:data<=16'd4893;
      32416:data<=16'd2560;
      32417:data<=16'd2144;
      32418:data<=16'd2206;
      32419:data<=16'd1686;
      32420:data<=16'd2177;
      32421:data<=16'd1695;
      32422:data<=-16'd352;
      32423:data<=-16'd1099;
      32424:data<=-16'd813;
      32425:data<=-16'd905;
      32426:data<=-16'd945;
      32427:data<=-16'd1098;
      32428:data<=-16'd2109;
      32429:data<=-16'd3348;
      32430:data<=-16'd3468;
      32431:data<=-16'd3224;
      32432:data<=-16'd3442;
      32433:data<=-16'd3046;
      32434:data<=-16'd3386;
      32435:data<=-16'd5256;
      32436:data<=-16'd5579;
      32437:data<=-16'd4931;
      32438:data<=-16'd5169;
      32439:data<=-16'd4681;
      32440:data<=-16'd5072;
      32441:data<=-16'd7138;
      32442:data<=-16'd7310;
      32443:data<=-16'd6652;
      32444:data<=-16'd6878;
      32445:data<=-16'd6351;
      32446:data<=-16'd6639;
      32447:data<=-16'd8049;
      32448:data<=-16'd8263;
      32449:data<=-16'd7976;
      32450:data<=-16'd7670;
      32451:data<=-16'd7559;
      32452:data<=-16'd7770;
      32453:data<=-16'd7699;
      32454:data<=-16'd10490;
      32455:data<=-16'd15162;
      32456:data<=-16'd15749;
      32457:data<=-16'd14607;
      32458:data<=-16'd14810;
      32459:data<=-16'd14722;
      32460:data<=-16'd15538;
      32461:data<=-16'd15747;
      32462:data<=-16'd14293;
      32463:data<=-16'd14389;
      32464:data<=-16'd14154;
      32465:data<=-16'd13306;
      32466:data<=-16'd14471;
      32467:data<=-16'd14317;
      32468:data<=-16'd12771;
      32469:data<=-16'd12786;
      32470:data<=-16'd12639;
      32471:data<=-16'd12333;
      32472:data<=-16'd12818;
      32473:data<=-16'd12998;
      32474:data<=-16'd12790;
      32475:data<=-16'd12330;
      32476:data<=-16'd11859;
      32477:data<=-16'd11303;
      32478:data<=-16'd11342;
      32479:data<=-16'd12715;
      32480:data<=-16'd12612;
      32481:data<=-16'd11229;
      32482:data<=-16'd11057;
      32483:data<=-16'd10281;
      32484:data<=-16'd10063;
      32485:data<=-16'd11620;
      32486:data<=-16'd11395;
      32487:data<=-16'd10307;
      32488:data<=-16'd10029;
      32489:data<=-16'd9312;
      32490:data<=-16'd9351;
      32491:data<=-16'd9919;
      32492:data<=-16'd9765;
      32493:data<=-16'd9527;
      32494:data<=-16'd9025;
      32495:data<=-16'd8307;
      32496:data<=-16'd7829;
      32497:data<=-16'd8131;
      32498:data<=-16'd8652;
      32499:data<=-16'd8011;
      32500:data<=-16'd7803;
      32501:data<=-16'd7712;
      32502:data<=-16'd6667;
      32503:data<=-16'd6990;
      32504:data<=-16'd5069;
      32505:data<=16'd526;
      32506:data<=16'd2358;
      32507:data<=16'd1240;
      32508:data<=16'd1695;
      32509:data<=16'd2608;
      32510:data<=16'd4211;
      32511:data<=16'd4858;
      32512:data<=16'd3987;
      32513:data<=16'd4373;
      32514:data<=16'd4313;
      32515:data<=16'd4350;
      32516:data<=16'd6331;
      32517:data<=16'd6839;
      32518:data<=16'd6056;
      32519:data<=16'd5918;
      32520:data<=16'd5689;
      32521:data<=16'd6167;
      32522:data<=16'd7235;
      32523:data<=16'd8093;
      32524:data<=16'd8539;
      32525:data<=16'd8234;
      32526:data<=16'd7968;
      32527:data<=16'd7611;
      32528:data<=16'd8214;
      32529:data<=16'd10292;
      32530:data<=16'd10305;
      32531:data<=16'd9377;
      32532:data<=16'd9809;
      32533:data<=16'd9212;
      32534:data<=16'd9283;
      32535:data<=16'd10863;
      32536:data<=16'd10881;
      32537:data<=16'd10455;
      32538:data<=16'd10228;
      32539:data<=16'd9611;
      32540:data<=16'd9919;
      32541:data<=16'd10593;
      32542:data<=16'd10972;
      32543:data<=16'd10866;
      32544:data<=16'd10329;
      32545:data<=16'd10120;
      32546:data<=16'd9614;
      32547:data<=16'd10060;
      32548:data<=16'd11253;
      32549:data<=16'd10425;
      32550:data<=16'd10182;
      32551:data<=16'd10502;
      32552:data<=16'd9219;
      32553:data<=16'd10464;
      32554:data<=16'd10812;
      32555:data<=16'd5782;
      32556:data<=16'd3450;
      32557:data<=16'd4775;
      32558:data<=16'd4044;
      32559:data<=16'd4037;
      32560:data<=16'd5609;
      32561:data<=16'd5956;
      32562:data<=16'd5791;
      32563:data<=16'd5709;
      32564:data<=16'd5553;
      32565:data<=16'd5536;
      32566:data<=16'd6255;
      32567:data<=16'd7313;
      32568:data<=16'd6978;
      32569:data<=16'd6727;
      32570:data<=16'd7213;
      32571:data<=16'd6294;
      32572:data<=16'd6332;
      32573:data<=16'd7952;
      32574:data<=16'd7429;
      32575:data<=16'd6605;
      32576:data<=16'd7113;
      32577:data<=16'd6357;
      32578:data<=16'd6032;
      32579:data<=16'd7500;
      32580:data<=16'd7783;
      32581:data<=16'd7094;
      32582:data<=16'd6975;
      32583:data<=16'd6435;
      32584:data<=16'd6304;
      32585:data<=16'd7460;
      32586:data<=16'd7806;
      32587:data<=16'd7313;
      32588:data<=16'd7363;
      32589:data<=16'd6761;
      32590:data<=16'd6097;
      32591:data<=16'd7227;
      32592:data<=16'd8193;
      32593:data<=16'd7655;
      32594:data<=16'd7141;
      32595:data<=16'd6875;
      32596:data<=16'd6593;
      32597:data<=16'd6821;
      32598:data<=16'd7388;
      32599:data<=16'd7316;
      32600:data<=16'd6492;
      32601:data<=16'd6546;
      32602:data<=16'd6802;
      32603:data<=16'd5357;
      32604:data<=16'd5856;
      32605:data<=16'd9861;
      32606:data<=16'd11582;
      32607:data<=16'd10381;
      32608:data<=16'd10060;
      32609:data<=16'd9312;
      32610:data<=16'd7471;
      32611:data<=16'd6464;
      32612:data<=16'd5849;
      32613:data<=16'd5218;
      32614:data<=16'd4945;
      32615:data<=16'd4379;
      32616:data<=16'd3030;
      32617:data<=16'd1542;
      32618:data<=16'd1043;
      32619:data<=16'd870;
      32620:data<=16'd334;
      32621:data<=16'd470;
      32622:data<=-16'd153;
      32623:data<=-16'd2127;
      32624:data<=-16'd2391;
      32625:data<=-16'd2002;
      32626:data<=-16'd2875;
      32627:data<=-16'd2776;
      32628:data<=-16'd2801;
      32629:data<=-16'd4449;
      32630:data<=-16'd5031;
      32631:data<=-16'd4804;
      32632:data<=-16'd5136;
      32633:data<=-16'd4766;
      32634:data<=-16'd4723;
      32635:data<=-16'd6167;
      32636:data<=-16'd7110;
      32637:data<=-16'd6930;
      32638:data<=-16'd6925;
      32639:data<=-16'd6940;
      32640:data<=-16'd6760;
      32641:data<=-16'd7791;
      32642:data<=-16'd9480;
      32643:data<=-16'd9433;
      32644:data<=-16'd8630;
      32645:data<=-16'd8674;
      32646:data<=-16'd8431;
      32647:data<=-16'd8701;
      32648:data<=-16'd10308;
      32649:data<=-16'd10666;
      32650:data<=-16'd9752;
      32651:data<=-16'd9718;
      32652:data<=-16'd9538;
      32653:data<=-16'd9169;
      32654:data<=-16'd11417;
      32655:data<=-16'd15587;
      32656:data<=-16'd17647;
      32657:data<=-16'd16979;
      32658:data<=-16'd16210;
      32659:data<=-16'd16311;
      32660:data<=-16'd16985;
      32661:data<=-16'd17675;
      32662:data<=-16'd17085;
      32663:data<=-16'd15934;
      32664:data<=-16'd15587;
      32665:data<=-16'd15185;
      32666:data<=-16'd15238;
      32667:data<=-16'd16126;
      32668:data<=-16'd15634;
      32669:data<=-16'd14530;
      32670:data<=-16'd14442;
      32671:data<=-16'd13966;
      32672:data<=-16'd13870;
      32673:data<=-16'd14875;
      32674:data<=-16'd14781;
      32675:data<=-16'd14104;
      32676:data<=-16'd13872;
      32677:data<=-16'd13029;
      32678:data<=-16'd12824;
      32679:data<=-16'd13923;
      32680:data<=-16'd14129;
      32681:data<=-16'd13391;
      32682:data<=-16'd12856;
      32683:data<=-16'd11963;
      32684:data<=-16'd11342;
      32685:data<=-16'd12416;
      32686:data<=-16'd13511;
      32687:data<=-16'd12769;
      32688:data<=-16'd11765;
      32689:data<=-16'd11157;
      32690:data<=-16'd10075;
      32691:data<=-16'd10103;
      32692:data<=-16'd11306;
      32693:data<=-16'd11050;
      32694:data<=-16'd10113;
      32695:data<=-16'd9867;
      32696:data<=-16'd9094;
      32697:data<=-16'd8869;
      32698:data<=-16'd10091;
      32699:data<=-16'd10246;
      32700:data<=-16'd9385;
      32701:data<=-16'd8995;
      32702:data<=-16'd8069;
      32703:data<=-16'd7415;
      32704:data<=-16'd6983;
      32705:data<=-16'd3597;
      32706:data<=16'd277;
      32707:data<=16'd649;
      32708:data<=16'd429;
      32709:data<=16'd1406;
      32710:data<=16'd2314;
      32711:data<=16'd3422;
      32712:data<=16'd3765;
      32713:data<=16'd3356;
      32714:data<=16'd3629;
      32715:data<=16'd3727;
      32716:data<=16'd4352;
      32717:data<=16'd5946;
      32718:data<=16'd6006;
      32719:data<=16'd5336;
      32720:data<=16'd5530;
      32721:data<=16'd5435;
      32722:data<=16'd5791;
      32723:data<=16'd7056;
      32724:data<=16'd7562;
      32725:data<=16'd7448;
      32726:data<=16'd7479;
      32727:data<=16'd7268;
      32728:data<=16'd7233;
      32729:data<=16'd8305;
      32730:data<=16'd9380;
      32731:data<=16'd9033;
      32732:data<=16'd8634;
      32733:data<=16'd8675;
      32734:data<=16'd8244;
      32735:data<=16'd9050;
      32736:data<=16'd10625;
      32737:data<=16'd10102;
      32738:data<=16'd9250;
      32739:data<=16'd9520;
      32740:data<=16'd8987;
      32741:data<=16'd8815;
      32742:data<=16'd10123;
      32743:data<=16'd10516;
      32744:data<=16'd10028;
      32745:data<=16'd10113;
      32746:data<=16'd9556;
      32747:data<=16'd8939;
      32748:data<=16'd10143;
      32749:data<=16'd11030;
      32750:data<=16'd10480;
      32751:data<=16'd10378;
      32752:data<=16'd9800;
      32753:data<=16'd9210;
      32754:data<=16'd10446;
      32755:data<=16'd9315;
      32756:data<=16'd4945;
      32757:data<=16'd3538;
      32758:data<=16'd4438;
      32759:data<=16'd3909;
      32760:data<=16'd4331;
      32761:data<=16'd5702;
      32762:data<=16'd5436;
      32763:data<=16'd5131;
      32764:data<=16'd5213;
      32765:data<=16'd4467;
      32766:data<=16'd4798;
      32767:data<=16'd6156;
      32768:data<=16'd6305;
      32769:data<=16'd6326;
      32770:data<=16'd6602;
      32771:data<=16'd5971;
      32772:data<=16'd6131;
      32773:data<=16'd7439;
      32774:data<=16'd7815;
      32775:data<=16'd7377;
      32776:data<=16'd6834;
      32777:data<=16'd6351;
      32778:data<=16'd6490;
      32779:data<=16'd7186;
      32780:data<=16'd7814;
      32781:data<=16'd7559;
      32782:data<=16'd6883;
      32783:data<=16'd6702;
      32784:data<=16'd6096;
      32785:data<=16'd6059;
      32786:data<=16'd7524;
      32787:data<=16'd7653;
      32788:data<=16'd6959;
      32789:data<=16'd7047;
      32790:data<=16'd6158;
      32791:data<=16'd6255;
      32792:data<=16'd8119;
      32793:data<=16'd8106;
      32794:data<=16'd7301;
      32795:data<=16'd7039;
      32796:data<=16'd6297;
      32797:data<=16'd6807;
      32798:data<=16'd7814;
      32799:data<=16'd7683;
      32800:data<=16'd7556;
      32801:data<=16'd6854;
      32802:data<=16'd6411;
      32803:data<=16'd6716;
      32804:data<=16'd5689;
      32805:data<=16'd6795;
      32806:data<=16'd10950;
      32807:data<=16'd11668;
      32808:data<=16'd10032;
      32809:data<=16'd9959;
      32810:data<=16'd8842;
      32811:data<=16'd7072;
      32812:data<=16'd6520;
      32813:data<=16'd5665;
      32814:data<=16'd5160;
      32815:data<=16'd5238;
      32816:data<=16'd4182;
      32817:data<=16'd2933;
      32818:data<=16'd2270;
      32819:data<=16'd1515;
      32820:data<=16'd1122;
      32821:data<=16'd1071;
      32822:data<=16'd563;
      32823:data<=-16'd541;
      32824:data<=-16'd1673;
      32825:data<=-16'd2035;
      32826:data<=-16'd2137;
      32827:data<=-16'd2637;
      32828:data<=-16'd2902;
      32829:data<=-16'd3503;
      32830:data<=-16'd4681;
      32831:data<=-16'd4778;
      32832:data<=-16'd4645;
      32833:data<=-16'd5263;
      32834:data<=-16'd4872;
      32835:data<=-16'd4884;
      32836:data<=-16'd6587;
      32837:data<=-16'd6899;
      32838:data<=-16'd6514;
      32839:data<=-16'd7210;
      32840:data<=-16'd6646;
      32841:data<=-16'd6411;
      32842:data<=-16'd8304;
      32843:data<=-16'd8950;
      32844:data<=-16'd8570;
      32845:data<=-16'd8686;
      32846:data<=-16'd7947;
      32847:data<=-16'd7920;
      32848:data<=-16'd9427;
      32849:data<=-16'd10263;
      32850:data<=-16'd10060;
      32851:data<=-16'd9415;
      32852:data<=-16'd9332;
      32853:data<=-16'd9535;
      32854:data<=-16'd9362;
      32855:data<=-16'd12017;
      32856:data<=-16'd16449;
      32857:data<=-16'd17247;
      32858:data<=-16'd16151;
      32859:data<=-16'd15894;
      32860:data<=-16'd15793;
      32861:data<=-16'd16566;
      32862:data<=-16'd16751;
      32863:data<=-16'd15820;
      32864:data<=-16'd15588;
      32865:data<=-16'd14518;
      32866:data<=-16'd13878;
      32867:data<=-16'd15599;
      32868:data<=-16'd15766;
      32869:data<=-16'd14266;
      32870:data<=-16'd13759;
      32871:data<=-16'd13110;
      32872:data<=-16'd12897;
      32873:data<=-16'd13828;
      32874:data<=-16'd14164;
      32875:data<=-16'd13628;
      32876:data<=-16'd12759;
      32877:data<=-16'd11970;
      32878:data<=-16'd11347;
      32879:data<=-16'd11285;
      32880:data<=-16'd12422;
      32881:data<=-16'd12734;
      32882:data<=-16'd11599;
      32883:data<=-16'd10933;
      32884:data<=-16'd10160;
      32885:data<=-16'd10035;
      32886:data<=-16'd11476;
      32887:data<=-16'd11582;
      32888:data<=-16'd10551;
      32889:data<=-16'd10170;
      32890:data<=-16'd9448;
      32891:data<=-16'd9241;
      32892:data<=-16'd10064;
      32893:data<=-16'd10035;
      32894:data<=-16'd9216;
      32895:data<=-16'd8801;
      32896:data<=-16'd8460;
      32897:data<=-16'd7645;
      32898:data<=-16'd7644;
      32899:data<=-16'd8602;
      32900:data<=-16'd8325;
      32901:data<=-16'd7451;
      32902:data<=-16'd6884;
      32903:data<=-16'd5952;
      32904:data<=-16'd5946;
      32905:data<=-16'd4508;
      32906:data<=16'd271;
      32907:data<=16'd2716;
      32908:data<=16'd2043;
      32909:data<=16'd2532;
      32910:data<=16'd3488;
      32911:data<=16'd4238;
      32912:data<=16'd4995;
      32913:data<=16'd5159;
      32914:data<=16'd5266;
      32915:data<=16'd4846;
      32916:data<=16'd4902;
      32917:data<=16'd6502;
      32918:data<=16'd7301;
      32919:data<=16'd7241;
      32920:data<=16'd7250;
      32921:data<=16'd6666;
      32922:data<=16'd6610;
      32923:data<=16'd7491;
      32924:data<=16'd8542;
      32925:data<=16'd9145;
      32926:data<=16'd8736;
      32927:data<=16'd8417;
      32928:data<=16'd8398;
      32929:data<=16'd8836;
      32930:data<=16'd10463;
      32931:data<=16'd10851;
      32932:data<=16'd10093;
      32933:data<=16'd10238;
      32934:data<=16'd9777;
      32935:data<=16'd9909;
      32936:data<=16'd11552;
      32937:data<=16'd11767;
      32938:data<=16'd11236;
      32939:data<=16'd11065;
      32940:data<=16'd10508;
      32941:data<=16'd10672;
      32942:data<=16'd11582;
      32943:data<=16'd12116;
      32944:data<=16'd11758;
      32945:data<=16'd11348;
      32946:data<=16'd11505;
      32947:data<=16'd10508;
      32948:data<=16'd10235;
      32949:data<=16'd12044;
      32950:data<=16'd11934;
      32951:data<=16'd11217;
      32952:data<=16'd11341;
      32953:data<=16'd10025;
      32954:data<=16'd10625;
      32955:data<=16'd11242;
      32956:data<=16'd7203;
      32957:data<=16'd4793;
      32958:data<=16'd5460;
      32959:data<=16'd4760;
      32960:data<=16'd5145;
      32961:data<=16'd6663;
      32962:data<=16'd6743;
      32963:data<=16'd6416;
      32964:data<=16'd6199;
      32965:data<=16'd6293;
      32966:data<=16'd6492;
      32967:data<=16'd6839;
      32968:data<=16'd7912;
      32969:data<=16'd8026;
      32970:data<=16'd7521;
      32971:data<=16'd7453;
      32972:data<=16'd6614;
      32973:data<=16'd7127;
      32974:data<=16'd9124;
      32975:data<=16'd9022;
      32976:data<=16'd8331;
      32977:data<=16'd8213;
      32978:data<=16'd7303;
      32979:data<=16'd7712;
      32980:data<=16'd9138;
      32981:data<=16'd8846;
      32982:data<=16'd8307;
      32983:data<=16'd8294;
      32984:data<=16'd7491;
      32985:data<=16'd7397;
      32986:data<=16'd8637;
      32987:data<=16'd8859;
      32988:data<=16'd8193;
      32989:data<=16'd8123;
      32990:data<=16'd7739;
      32991:data<=16'd7197;
      32992:data<=16'd7899;
      32993:data<=16'd8869;
      32994:data<=16'd8760;
      32995:data<=16'd8002;
      32996:data<=16'd7394;
      32997:data<=16'd7250;
      32998:data<=16'd7726;
      32999:data<=16'd8668;
      33000:data<=16'd8781;
      33001:data<=16'd7832;
      33002:data<=16'd7676;
      33003:data<=16'd7714;
      33004:data<=16'd6616;
      33005:data<=16'd7189;
      33006:data<=16'd10398;
      33007:data<=16'd12266;
      33008:data<=16'd11721;
      33009:data<=16'd11176;
      33010:data<=16'd10319;
      33011:data<=16'd8316;
      33012:data<=16'd6948;
      33013:data<=16'd6649;
      33014:data<=16'd6264;
      33015:data<=16'd5894;
      33016:data<=16'd5280;
      33017:data<=16'd3894;
      33018:data<=16'd2596;
      33019:data<=16'd1900;
      33020:data<=16'd1416;
      33021:data<=16'd1251;
      33022:data<=16'd1336;
      33023:data<=16'd326;
      33024:data<=-16'd1621;
      33025:data<=-16'd2364;
      33026:data<=-16'd2496;
      33027:data<=-16'd2849;
      33028:data<=-16'd2188;
      33029:data<=-16'd2549;
      33030:data<=-16'd4631;
      33031:data<=-16'd5103;
      33032:data<=-16'd4837;
      33033:data<=-16'd5198;
      33034:data<=-16'd4784;
      33035:data<=-16'd5036;
      33036:data<=-16'd6481;
      33037:data<=-16'd7245;
      33038:data<=-16'd7286;
      33039:data<=-16'd7283;
      33040:data<=-16'd7401;
      33041:data<=-16'd7116;
      33042:data<=-16'd7291;
      33043:data<=-16'd9010;
      33044:data<=-16'd9677;
      33045:data<=-16'd9119;
      33046:data<=-16'd9262;
      33047:data<=-16'd8605;
      33048:data<=-16'd8599;
      33049:data<=-16'd10568;
      33050:data<=-16'd11106;
      33051:data<=-16'd10546;
      33052:data<=-16'd10537;
      33053:data<=-16'd10132;
      33054:data<=-16'd10184;
      33055:data<=-16'd12087;
      33056:data<=-16'd15719;
      33057:data<=-16'd18175;
      33058:data<=-16'd17567;
      33059:data<=-16'd16918;
      33060:data<=-16'd16935;
      33061:data<=-16'd16965;
      33062:data<=-16'd17901;
      33063:data<=-16'd17452;
      33064:data<=-16'd16284;
      33065:data<=-16'd16316;
      33066:data<=-16'd15080;
      33067:data<=-16'd14772;
      33068:data<=-16'd16647;
      33069:data<=-16'd16304;
      33070:data<=-16'd15141;
      33071:data<=-16'd14894;
      33072:data<=-16'd13835;
      33073:data<=-16'd13954;
      33074:data<=-16'd15329;
      33075:data<=-16'd15244;
      33076:data<=-16'd14186;
      33077:data<=-16'd13385;
      33078:data<=-16'd12980;
      33079:data<=-16'd13050;
      33080:data<=-16'd13894;
      33081:data<=-16'd14439;
      33082:data<=-16'd13323;
      33083:data<=-16'd12377;
      33084:data<=-16'd12172;
      33085:data<=-16'd11465;
      33086:data<=-16'd11844;
      33087:data<=-16'd12730;
      33088:data<=-16'd12037;
      33089:data<=-16'd11236;
      33090:data<=-16'd10786;
      33091:data<=-16'd10122;
      33092:data<=-16'd10320;
      33093:data<=-16'd11019;
      33094:data<=-16'd10798;
      33095:data<=-16'd10009;
      33096:data<=-16'd9749;
      33097:data<=-16'd9320;
      33098:data<=-16'd8790;
      33099:data<=-16'd9549;
      33100:data<=-16'd9565;
      33101:data<=-16'd8454;
      33102:data<=-16'd8684;
      33103:data<=-16'd8155;
      33104:data<=-16'd6986;
      33105:data<=-16'd7013;
      33106:data<=-16'd4225;
      33107:data<=16'd2;
      33108:data<=16'd726;
      33109:data<=16'd405;
      33110:data<=16'd798;
      33111:data<=16'd1676;
      33112:data<=16'd3200;
      33113:data<=16'd3338;
      33114:data<=16'd3247;
      33115:data<=16'd3762;
      33116:data<=16'd2966;
      33117:data<=16'd3321;
      33118:data<=16'd5145;
      33119:data<=16'd5442;
      33120:data<=16'd5557;
      33121:data<=16'd5582;
      33122:data<=16'd4626;
      33123:data<=16'd5295;
      33124:data<=16'd7228;
      33125:data<=16'd7662;
      33126:data<=16'd7156;
      33127:data<=16'd7156;
      33128:data<=16'd7221;
      33129:data<=16'd7147;
      33130:data<=16'd8106;
      33131:data<=16'd9253;
      33132:data<=16'd9006;
      33133:data<=16'd8957;
      33134:data<=16'd9121;
      33135:data<=16'd8152;
      33136:data<=16'd8466;
      33137:data<=16'd10169;
      33138:data<=16'd10182;
      33139:data<=16'd9576;
      33140:data<=16'd9539;
      33141:data<=16'd8913;
      33142:data<=16'd9227;
      33143:data<=16'd10800;
      33144:data<=16'd10872;
      33145:data<=16'd10241;
      33146:data<=16'd10414;
      33147:data<=16'd9791;
      33148:data<=16'd9505;
      33149:data<=16'd10983;
      33150:data<=16'd11291;
      33151:data<=16'd10445;
      33152:data<=16'd10665;
      33153:data<=16'd9988;
      33154:data<=16'd9248;
      33155:data<=16'd11171;
      33156:data<=16'd10815;
      33157:data<=16'd6061;
      33158:data<=16'd3953;
      33159:data<=16'd4854;
      33160:data<=16'd4108;
      33161:data<=16'd4504;
      33162:data<=16'd6601;
      33163:data<=16'd6438;
      33164:data<=16'd6038;
      33165:data<=16'd6501;
      33166:data<=16'd5749;
      33167:data<=16'd6219;
      33168:data<=16'd7932;
      33169:data<=16'd7850;
      33170:data<=16'd7526;
      33171:data<=16'd7548;
      33172:data<=16'd6713;
      33173:data<=16'd6796;
      33174:data<=16'd8105;
      33175:data<=16'd8816;
      33176:data<=16'd8651;
      33177:data<=16'd8052;
      33178:data<=16'd7318;
      33179:data<=16'd7013;
      33180:data<=16'd7794;
      33181:data<=16'd8724;
      33182:data<=16'd8354;
      33183:data<=16'd7882;
      33184:data<=16'd7746;
      33185:data<=16'd6940;
      33186:data<=16'd7292;
      33187:data<=16'd8751;
      33188:data<=16'd8498;
      33189:data<=16'd7791;
      33190:data<=16'd7774;
      33191:data<=16'd6909;
      33192:data<=16'd6918;
      33193:data<=16'd8410;
      33194:data<=16'd8361;
      33195:data<=16'd7653;
      33196:data<=16'd7715;
      33197:data<=16'd6928;
      33198:data<=16'd6711;
      33199:data<=16'd7888;
      33200:data<=16'd8090;
      33201:data<=16'd7656;
      33202:data<=16'd7197;
      33203:data<=16'd6855;
      33204:data<=16'd7078;
      33205:data<=16'd6091;
      33206:data<=16'd6566;
      33207:data<=16'd10683;
      33208:data<=16'd11900;
      33209:data<=16'd10292;
      33210:data<=16'd10636;
      33211:data<=16'd9357;
      33212:data<=16'd6731;
      33213:data<=16'd6228;
      33214:data<=16'd5565;
      33215:data<=16'd5197;
      33216:data<=16'd5513;
      33217:data<=16'd3883;
      33218:data<=16'd1961;
      33219:data<=16'd1406;
      33220:data<=16'd1202;
      33221:data<=16'd948;
      33222:data<=16'd616;
      33223:data<=16'd241;
      33224:data<=-16'd1042;
      33225:data<=-16'd2464;
      33226:data<=-16'd2549;
      33227:data<=-16'd2963;
      33228:data<=-16'd3169;
      33229:data<=-16'd2461;
      33230:data<=-16'd3645;
      33231:data<=-16'd5385;
      33232:data<=-16'd5521;
      33233:data<=-16'd5632;
      33234:data<=-16'd5456;
      33235:data<=-16'd5018;
      33236:data<=-16'd5940;
      33237:data<=-16'd7494;
      33238:data<=-16'd7934;
      33239:data<=-16'd7413;
      33240:data<=-16'd7344;
      33241:data<=-16'd7382;
      33242:data<=-16'd7577;
      33243:data<=-16'd8921;
      33244:data<=-16'd9356;
      33245:data<=-16'd8950;
      33246:data<=-16'd9335;
      33247:data<=-16'd8728;
      33248:data<=-16'd8537;
      33249:data<=-16'd9976;
      33250:data<=-16'd10477;
      33251:data<=-16'd10710;
      33252:data<=-16'd10684;
      33253:data<=-16'd10006;
      33254:data<=-16'd10181;
      33255:data<=-16'd10392;
      33256:data<=-16'd12797;
      33257:data<=-16'd17344;
      33258:data<=-16'd18227;
      33259:data<=-16'd17112;
      33260:data<=-16'd16936;
      33261:data<=-16'd16572;
      33262:data<=-16'd17306;
      33263:data<=-16'd17341;
      33264:data<=-16'd16255;
      33265:data<=-16'd16421;
      33266:data<=-16'd15402;
      33267:data<=-16'd14610;
      33268:data<=-16'd16042;
      33269:data<=-16'd16099;
      33270:data<=-16'd15452;
      33271:data<=-16'd15006;
      33272:data<=-16'd13820;
      33273:data<=-16'd13843;
      33274:data<=-16'd14578;
      33275:data<=-16'd14897;
      33276:data<=-16'd14571;
      33277:data<=-16'd13247;
      33278:data<=-16'd12704;
      33279:data<=-16'd12446;
      33280:data<=-16'd12328;
      33281:data<=-16'd13418;
      33282:data<=-16'd13120;
      33283:data<=-16'd12258;
      33284:data<=-16'd12149;
      33285:data<=-16'd10851;
      33286:data<=-16'd10945;
      33287:data<=-16'd12196;
      33288:data<=-16'd11681;
      33289:data<=-16'd11630;
      33290:data<=-16'd11333;
      33291:data<=-16'd9741;
      33292:data<=-16'd9638;
      33293:data<=-16'd10545;
      33294:data<=-16'd10872;
      33295:data<=-16'd10266;
      33296:data<=-16'd9454;
      33297:data<=-16'd9144;
      33298:data<=-16'd8299;
      33299:data<=-16'd8636;
      33300:data<=-16'd9752;
      33301:data<=-16'd8683;
      33302:data<=-16'd8237;
      33303:data<=-16'd8120;
      33304:data<=-16'd6570;
      33305:data<=-16'd6790;
      33306:data<=-16'd5271;
      33307:data<=-16'd458;
      33308:data<=16'd1193;
      33309:data<=16'd848;
      33310:data<=16'd1494;
      33311:data<=16'd2197;
      33312:data<=16'd3627;
      33313:data<=16'd4184;
      33314:data<=16'd3779;
      33315:data<=16'd4309;
      33316:data<=16'd4258;
      33317:data<=16'd4349;
      33318:data<=16'd5629;
      33319:data<=16'd6167;
      33320:data<=16'd6179;
      33321:data<=16'd6219;
      33322:data<=16'd5955;
      33323:data<=16'd6038;
      33324:data<=16'd7113;
      33325:data<=16'd8716;
      33326:data<=16'd8866;
      33327:data<=16'd7952;
      33328:data<=16'd7811;
      33329:data<=16'd7683;
      33330:data<=16'd8343;
      33331:data<=16'd9990;
      33332:data<=16'd10110;
      33333:data<=16'd9677;
      33334:data<=16'd9673;
      33335:data<=16'd9250;
      33336:data<=16'd9709;
      33337:data<=16'd10646;
      33338:data<=16'd10828;
      33339:data<=16'd10948;
      33340:data<=16'd10800;
      33341:data<=16'd10317;
      33342:data<=16'd10208;
      33343:data<=16'd10997;
      33344:data<=16'd12029;
      33345:data<=16'd11585;
      33346:data<=16'd11035;
      33347:data<=16'd11126;
      33348:data<=16'd10208;
      33349:data<=16'd10742;
      33350:data<=16'd12424;
      33351:data<=16'd11502;
      33352:data<=16'd10968;
      33353:data<=16'd11420;
      33354:data<=16'd10287;
      33355:data<=16'd11186;
      33356:data<=16'd11976;
      33357:data<=16'd7827;
      33358:data<=16'd4975;
      33359:data<=16'd5727;
      33360:data<=16'd5075;
      33361:data<=16'd4896;
      33362:data<=16'd6701;
      33363:data<=16'd7203;
      33364:data<=16'd6605;
      33365:data<=16'd6319;
      33366:data<=16'd6043;
      33367:data<=16'd6000;
      33368:data<=16'd6796;
      33369:data<=16'd7978;
      33370:data<=16'd7861;
      33371:data<=16'd7178;
      33372:data<=16'd7413;
      33373:data<=16'd6934;
      33374:data<=16'd6721;
      33375:data<=16'd8294;
      33376:data<=16'd8631;
      33377:data<=16'd7999;
      33378:data<=16'd8062;
      33379:data<=16'd7274;
      33380:data<=16'd7350;
      33381:data<=16'd8872;
      33382:data<=16'd8849;
      33383:data<=16'd8352;
      33384:data<=16'd8282;
      33385:data<=16'd7400;
      33386:data<=16'd7262;
      33387:data<=16'd8534;
      33388:data<=16'd9382;
      33389:data<=16'd9004;
      33390:data<=16'd8361;
      33391:data<=16'd8082;
      33392:data<=16'd7386;
      33393:data<=16'd7448;
      33394:data<=16'd8904;
      33395:data<=16'd8969;
      33396:data<=16'd8119;
      33397:data<=16'd8019;
      33398:data<=16'd7389;
      33399:data<=16'd7377;
      33400:data<=16'd8549;
      33401:data<=16'd8683;
      33402:data<=16'd8120;
      33403:data<=16'd7890;
      33404:data<=16'd7553;
      33405:data<=16'd6669;
      33406:data<=16'd6699;
      33407:data<=16'd9881;
      33408:data<=16'd12747;
      33409:data<=16'd12007;
      33410:data<=16'd11276;
      33411:data<=16'd10754;
      33412:data<=16'd8419;
      33413:data<=16'd7151;
      33414:data<=16'd7127;
      33415:data<=16'd6448;
      33416:data<=16'd6184;
      33417:data<=16'd5937;
      33418:data<=16'd4411;
      33419:data<=16'd2663;
      33420:data<=16'd2111;
      33421:data<=16'd2118;
      33422:data<=16'd1659;
      33423:data<=16'd1453;
      33424:data<=16'd670;
      33425:data<=-16'd1251;
      33426:data<=-16'd1701;
      33427:data<=-16'd1448;
      33428:data<=-16'd2040;
      33429:data<=-16'd1685;
      33430:data<=-16'd1988;
      33431:data<=-16'd3868;
      33432:data<=-16'd4482;
      33433:data<=-16'd4517;
      33434:data<=-16'd4734;
      33435:data<=-16'd4106;
      33436:data<=-16'd4225;
      33437:data<=-16'd5727;
      33438:data<=-16'd6975;
      33439:data<=-16'd7065;
      33440:data<=-16'd6684;
      33441:data<=-16'd6692;
      33442:data<=-16'd6531;
      33443:data<=-16'd7065;
      33444:data<=-16'd8604;
      33445:data<=-16'd8719;
      33446:data<=-16'd8363;
      33447:data<=-16'd8583;
      33448:data<=-16'd7874;
      33449:data<=-16'd8276;
      33450:data<=-16'd9790;
      33451:data<=-16'd9747;
      33452:data<=-16'd9633;
      33453:data<=-16'd9694;
      33454:data<=-16'd8951;
      33455:data<=-16'd8919;
      33456:data<=-16'd10386;
      33457:data<=-16'd13782;
      33458:data<=-16'd16980;
      33459:data<=-16'd16944;
      33460:data<=-16'd15887;
      33461:data<=-16'd15590;
      33462:data<=-16'd15743;
      33463:data<=-16'd16550;
      33464:data<=-16'd16296;
      33465:data<=-16'd15599;
      33466:data<=-16'd15608;
      33467:data<=-16'd14492;
      33468:data<=-16'd14051;
      33469:data<=-16'd15135;
      33470:data<=-16'd14915;
      33471:data<=-16'd14455;
      33472:data<=-16'd14207;
      33473:data<=-16'd12977;
      33474:data<=-16'd12768;
      33475:data<=-16'd13717;
      33476:data<=-16'd13916;
      33477:data<=-16'd13273;
      33478:data<=-16'd12401;
      33479:data<=-16'd11849;
      33480:data<=-16'd11765;
      33481:data<=-16'd12440;
      33482:data<=-16'd12971;
      33483:data<=-16'd12061;
      33484:data<=-16'd11626;
      33485:data<=-16'd11659;
      33486:data<=-16'd10552;
      33487:data<=-16'd10836;
      33488:data<=-16'd12002;
      33489:data<=-16'd11314;
      33490:data<=-16'd10865;
      33491:data<=-16'd10760;
      33492:data<=-16'd9532;
      33493:data<=-16'd9497;
      33494:data<=-16'd10713;
      33495:data<=-16'd10602;
      33496:data<=-16'd9765;
      33497:data<=-16'd9603;
      33498:data<=-16'd8903;
      33499:data<=-16'd8128;
      33500:data<=-16'd9336;
      33501:data<=-16'd9859;
      33502:data<=-16'd8533;
      33503:data<=-16'd8573;
      33504:data<=-16'd8155;
      33505:data<=-16'd6949;
      33506:data<=-16'd7577;
      33507:data<=-16'd5292;
      33508:data<=-16'd308;
      33509:data<=16'd738;
      33510:data<=16'd253;
      33511:data<=16'd943;
      33512:data<=16'd1556;
      33513:data<=16'd3089;
      33514:data<=16'd3771;
      33515:data<=16'd3318;
      33516:data<=16'd3836;
      33517:data<=16'd3653;
      33518:data<=16'd3874;
      33519:data<=16'd5506;
      33520:data<=16'd5611;
      33521:data<=16'd5548;
      33522:data<=16'd6152;
      33523:data<=16'd5641;
      33524:data<=16'd5949;
      33525:data<=16'd7078;
      33526:data<=16'd7289;
      33527:data<=16'd7506;
      33528:data<=16'd7344;
      33529:data<=16'd6701;
      33530:data<=16'd7028;
      33531:data<=16'd7950;
      33532:data<=16'd8469;
      33533:data<=16'd8410;
      33534:data<=16'd8445;
      33535:data<=16'd8537;
      33536:data<=16'd7955;
      33537:data<=16'd8273;
      33538:data<=16'd9573;
      33539:data<=16'd9609;
      33540:data<=16'd9489;
      33541:data<=16'd9693;
      33542:data<=16'd8843;
      33543:data<=16'd8987;
      33544:data<=16'd10502;
      33545:data<=16'd10607;
      33546:data<=16'd9958;
      33547:data<=16'd9829;
      33548:data<=16'd9107;
      33549:data<=16'd8777;
      33550:data<=16'd10176;
      33551:data<=16'd10705;
      33552:data<=16'd9576;
      33553:data<=16'd9652;
      33554:data<=16'd9721;
      33555:data<=16'd8903;
      33556:data<=16'd10144;
      33557:data<=16'd9630;
      33558:data<=16'd4819;
      33559:data<=16'd3190;
      33560:data<=16'd4457;
      33561:data<=16'd3195;
      33562:data<=16'd3425;
      33563:data<=16'd5518;
      33564:data<=16'd5203;
      33565:data<=16'd4874;
      33566:data<=16'd4971;
      33567:data<=16'd3961;
      33568:data<=16'd4619;
      33569:data<=16'd6423;
      33570:data<=16'd6578;
      33571:data<=16'd5921;
      33572:data<=16'd5497;
      33573:data<=16'd5131;
      33574:data<=16'd5134;
      33575:data<=16'd6258;
      33576:data<=16'd7350;
      33577:data<=16'd6561;
      33578:data<=16'd5947;
      33579:data<=16'd6326;
      33580:data<=16'd5586;
      33581:data<=16'd5920;
      33582:data<=16'd7711;
      33583:data<=16'd7288;
      33584:data<=16'd6460;
      33585:data<=16'd6751;
      33586:data<=16'd5877;
      33587:data<=16'd5823;
      33588:data<=16'd7486;
      33589:data<=16'd7697;
      33590:data<=16'd7010;
      33591:data<=16'd6684;
      33592:data<=16'd5755;
      33593:data<=16'd5777;
      33594:data<=16'd7409;
      33595:data<=16'd7806;
      33596:data<=16'd6924;
      33597:data<=16'd6654;
      33598:data<=16'd6349;
      33599:data<=16'd6150;
      33600:data<=16'd6907;
      33601:data<=16'd7439;
      33602:data<=16'd7292;
      33603:data<=16'd6754;
      33604:data<=16'd6119;
      33605:data<=16'd5709;
      33606:data<=16'd4789;
      33607:data<=16'd5912;
      33608:data<=16'd10226;
      33609:data<=16'd11204;
      33610:data<=16'd9059;
      33611:data<=16'd9542;
      33612:data<=16'd8954;
      33613:data<=16'd6208;
      33614:data<=16'd5914;
      33615:data<=16'd5632;
      33616:data<=16'd4437;
      33617:data<=16'd4781;
      33618:data<=16'd4058;
      33619:data<=16'd1838;
      33620:data<=16'd1002;
      33621:data<=16'd1086;
      33622:data<=16'd716;
      33623:data<=16'd174;
      33624:data<=-16'd235;
      33625:data<=-16'd1386;
      33626:data<=-16'd2622;
      33627:data<=-16'd2463;
      33628:data<=-16'd2858;
      33629:data<=-16'd3798;
      33630:data<=-16'd3140;
      33631:data<=-16'd3541;
      33632:data<=-16'd5450;
      33633:data<=-16'd5745;
      33634:data<=-16'd5752;
      33635:data<=-16'd6253;
      33636:data<=-16'd5711;
      33637:data<=-16'd5827;
      33638:data<=-16'd7538;
      33639:data<=-16'd8423;
      33640:data<=-16'd7926;
      33641:data<=-16'd7597;
      33642:data<=-16'd7242;
      33643:data<=-16'd7189;
      33644:data<=-16'd8884;
      33645:data<=-16'd10026;
      33646:data<=-16'd9230;
      33647:data<=-16'd9115;
      33648:data<=-16'd9163;
      33649:data<=-16'd8677;
      33650:data<=-16'd9550;
      33651:data<=-16'd10561;
      33652:data<=-16'd10360;
      33653:data<=-16'd10009;
      33654:data<=-16'd9928;
      33655:data<=-16'd9667;
      33656:data<=-16'd9550;
      33657:data<=-16'd12222;
      33658:data<=-16'd16562;
      33659:data<=-16'd17379;
      33660:data<=-16'd16180;
      33661:data<=-16'd16069;
      33662:data<=-16'd16054;
      33663:data<=-16'd16832;
      33664:data<=-16'd17164;
      33665:data<=-16'd15767;
      33666:data<=-16'd15200;
      33667:data<=-16'd14882;
      33668:data<=-16'd14343;
      33669:data<=-16'd15086;
      33670:data<=-16'd15487;
      33671:data<=-16'd15079;
      33672:data<=-16'd14607;
      33673:data<=-16'd13705;
      33674:data<=-16'd13101;
      33675:data<=-16'd13352;
      33676:data<=-16'd14308;
      33677:data<=-16'd14317;
      33678:data<=-16'd12777;
      33679:data<=-16'd12176;
      33680:data<=-16'd11859;
      33681:data<=-16'd11462;
      33682:data<=-16'd12659;
      33683:data<=-16'd12700;
      33684:data<=-16'd11483;
      33685:data<=-16'd11159;
      33686:data<=-16'd10176;
      33687:data<=-16'd10090;
      33688:data<=-16'd11335;
      33689:data<=-16'd11098;
      33690:data<=-16'd10687;
      33691:data<=-16'd10533;
      33692:data<=-16'd9770;
      33693:data<=-16'd9424;
      33694:data<=-16'd9547;
      33695:data<=-16'd10176;
      33696:data<=-16'd10060;
      33697:data<=-16'd9030;
      33698:data<=-16'd8787;
      33699:data<=-16'd7785;
      33700:data<=-16'd7424;
      33701:data<=-16'd9213;
      33702:data<=-16'd9063;
      33703:data<=-16'd8034;
      33704:data<=-16'd7855;
      33705:data<=-16'd6781;
      33706:data<=-16'd6714;
      33707:data<=-16'd5486;
      33708:data<=-16'd1061;
      33709:data<=16'd1419;
      33710:data<=16'd1562;
      33711:data<=16'd1603;
      33712:data<=16'd1804;
      33713:data<=16'd3369;
      33714:data<=16'd4353;
      33715:data<=16'd4020;
      33716:data<=16'd4272;
      33717:data<=16'd4329;
      33718:data<=16'd4514;
      33719:data<=16'd5406;
      33720:data<=16'd6161;
      33721:data<=16'd6793;
      33722:data<=16'd6862;
      33723:data<=16'd6675;
      33724:data<=16'd6529;
      33725:data<=16'd6904;
      33726:data<=16'd8719;
      33727:data<=16'd9219;
      33728:data<=16'd8298;
      33729:data<=16'd8505;
      33730:data<=16'd7924;
      33731:data<=16'd7879;
      33732:data<=16'd9834;
      33733:data<=16'd10137;
      33734:data<=16'd9740;
      33735:data<=16'd9683;
      33736:data<=16'd8760;
      33737:data<=16'd9274;
      33738:data<=16'd10519;
      33739:data<=16'd10763;
      33740:data<=16'd10942;
      33741:data<=16'd10557;
      33742:data<=16'd10110;
      33743:data<=16'd9887;
      33744:data<=16'd10105;
      33745:data<=16'd11571;
      33746:data<=16'd11503;
      33747:data<=16'd10528;
      33748:data<=16'd10883;
      33749:data<=16'd9820;
      33750:data<=16'd9594;
      33751:data<=16'd11803;
      33752:data<=16'd11755;
      33753:data<=16'd11077;
      33754:data<=16'd11233;
      33755:data<=16'd10008;
      33756:data<=16'd10616;
      33757:data<=16'd11715;
      33758:data<=16'd8379;
      33759:data<=16'd4987;
      33760:data<=16'd5066;
      33761:data<=16'd5187;
      33762:data<=16'd4931;
      33763:data<=16'd5952;
      33764:data<=16'd6757;
      33765:data<=16'd6558;
      33766:data<=16'd6549;
      33767:data<=16'd6200;
      33768:data<=16'd5391;
      33769:data<=16'd6114;
      33770:data<=16'd7624;
      33771:data<=16'd7606;
      33772:data<=16'd6948;
      33773:data<=16'd6721;
      33774:data<=16'd6432;
      33775:data<=16'd6901;
      33776:data<=16'd8090;
      33777:data<=16'd8041;
      33778:data<=16'd7391;
      33779:data<=16'd7430;
      33780:data<=16'd7098;
      33781:data<=16'd7307;
      33782:data<=16'd8684;
      33783:data<=16'd8624;
      33784:data<=16'd7796;
      33785:data<=16'd8135;
      33786:data<=16'd7787;
      33787:data<=16'd6796;
      33788:data<=16'd7480;
      33789:data<=16'd8781;
      33790:data<=16'd8624;
      33791:data<=16'd8023;
      33792:data<=16'd7865;
      33793:data<=16'd7074;
      33794:data<=16'd7242;
      33795:data<=16'd9065;
      33796:data<=16'd8989;
      33797:data<=16'd7877;
      33798:data<=16'd7976;
      33799:data<=16'd7398;
      33800:data<=16'd7536;
      33801:data<=16'd8881;
      33802:data<=16'd8508;
      33803:data<=16'd7849;
      33804:data<=16'd7809;
      33805:data<=16'd7274;
      33806:data<=16'd6766;
      33807:data<=16'd6529;
      33808:data<=16'd8804;
      33809:data<=16'd12361;
      33810:data<=16'd11932;
      33811:data<=16'd10305;
      33812:data<=16'd10360;
      33813:data<=16'd8904;
      33814:data<=16'd7224;
      33815:data<=16'd6801;
      33816:data<=16'd5937;
      33817:data<=16'd5598;
      33818:data<=16'd5802;
      33819:data<=16'd4719;
      33820:data<=16'd2840;
      33821:data<=16'd1861;
      33822:data<=16'd1855;
      33823:data<=16'd1880;
      33824:data<=16'd2030;
      33825:data<=16'd1296;
      33826:data<=-16'd707;
      33827:data<=-16'd1407;
      33828:data<=-16'd1281;
      33829:data<=-16'd1647;
      33830:data<=-16'd1392;
      33831:data<=-16'd2056;
      33832:data<=-16'd3762;
      33833:data<=-16'd4278;
      33834:data<=-16'd4361;
      33835:data<=-16'd4416;
      33836:data<=-16'd4215;
      33837:data<=-16'd4164;
      33838:data<=-16'd4523;
      33839:data<=-16'd6087;
      33840:data<=-16'd6945;
      33841:data<=-16'd6329;
      33842:data<=-16'd6334;
      33843:data<=-16'd5824;
      33844:data<=-16'd5993;
      33845:data<=-16'd8294;
      33846:data<=-16'd8775;
      33847:data<=-16'd8006;
      33848:data<=-16'd7808;
      33849:data<=-16'd6969;
      33850:data<=-16'd7744;
      33851:data<=-16'd9282;
      33852:data<=-16'd9242;
      33853:data<=-16'd9347;
      33854:data<=-16'd8966;
      33855:data<=-16'd8633;
      33856:data<=-16'd9156;
      33857:data<=-16'd9182;
      33858:data<=-16'd12026;
      33859:data<=-16'd16410;
      33860:data<=-16'd16662;
      33861:data<=-16'd15471;
      33862:data<=-16'd15094;
      33863:data<=-16'd14985;
      33864:data<=-16'd16177;
      33865:data<=-16'd16048;
      33866:data<=-16'd14604;
      33867:data<=-16'd14404;
      33868:data<=-16'd13869;
      33869:data<=-16'd13899;
      33870:data<=-16'd15098;
      33871:data<=-16'd14595;
      33872:data<=-16'd13626;
      33873:data<=-16'd13637;
      33874:data<=-16'd13126;
      33875:data<=-16'd12845;
      33876:data<=-16'd13673;
      33877:data<=-16'd13825;
      33878:data<=-16'd12671;
      33879:data<=-16'd12187;
      33880:data<=-16'd12041;
      33881:data<=-16'd11024;
      33882:data<=-16'd11476;
      33883:data<=-16'd12481;
      33884:data<=-16'd11324;
      33885:data<=-16'd10757;
      33886:data<=-16'd10771;
      33887:data<=-16'd9574;
      33888:data<=-16'd10105;
      33889:data<=-16'd11203;
      33890:data<=-16'd10201;
      33891:data<=-16'd9705;
      33892:data<=-16'd9753;
      33893:data<=-16'd8834;
      33894:data<=-16'd8772;
      33895:data<=-16'd9674;
      33896:data<=-16'd9564;
      33897:data<=-16'd8710;
      33898:data<=-16'd8323;
      33899:data<=-16'd7589;
      33900:data<=-16'd6951;
      33901:data<=-16'd8276;
      33902:data<=-16'd8986;
      33903:data<=-16'd7638;
      33904:data<=-16'd7248;
      33905:data<=-16'd6842;
      33906:data<=-16'd5940;
      33907:data<=-16'd6297;
      33908:data<=-16'd4058;
      33909:data<=16'd842;
      33910:data<=16'd2681;
      33911:data<=16'd2250;
      33912:data<=16'd2329;
      33913:data<=16'd3033;
      33914:data<=16'd4467;
      33915:data<=16'd4946;
      33916:data<=16'd4683;
      33917:data<=16'd5112;
      33918:data<=16'd4986;
      33919:data<=16'd5489;
      33920:data<=16'd7192;
      33921:data<=16'd7435;
      33922:data<=16'd7213;
      33923:data<=16'd7479;
      33924:data<=16'd7109;
      33925:data<=16'd7550;
      33926:data<=16'd8604;
      33927:data<=16'd8783;
      33928:data<=16'd8807;
      33929:data<=16'd8583;
      33930:data<=16'd8249;
      33931:data<=16'd8392;
      33932:data<=16'd8689;
      33933:data<=16'd9505;
      33934:data<=16'd9961;
      33935:data<=16'd9517;
      33936:data<=16'd9206;
      33937:data<=16'd8599;
      33938:data<=16'd9041;
      33939:data<=16'd10951;
      33940:data<=16'd10856;
      33941:data<=16'd9887;
      33942:data<=16'd10040;
      33943:data<=16'd9386;
      33944:data<=16'd9497;
      33945:data<=16'd10942;
      33946:data<=16'd10809;
      33947:data<=16'd10135;
      33948:data<=16'd10208;
      33949:data<=16'd9875;
      33950:data<=16'd9550;
      33951:data<=16'd10202;
      33952:data<=16'd11032;
      33953:data<=16'd10724;
      33954:data<=16'd10240;
      33955:data<=16'd9721;
      33956:data<=16'd8589;
      33957:data<=16'd9647;
      33958:data<=16'd10073;
      33959:data<=16'd5588;
      33960:data<=16'd3131;
      33961:data<=16'd4250;
      33962:data<=16'd3294;
      33963:data<=16'd3714;
      33964:data<=16'd5786;
      33965:data<=16'd5277;
      33966:data<=16'd5016;
      33967:data<=16'd5222;
      33968:data<=16'd4259;
      33969:data<=16'd4541;
      33970:data<=16'd5777;
      33971:data<=16'd6290;
      33972:data<=16'd5941;
      33973:data<=16'd5407;
      33974:data<=16'd5110;
      33975:data<=16'd4501;
      33976:data<=16'd5406;
      33977:data<=16'd7084;
      33978:data<=16'd6205;
      33979:data<=16'd5615;
      33980:data<=16'd6018;
      33981:data<=16'd4958;
      33982:data<=16'd5603;
      33983:data<=16'd7374;
      33984:data<=16'd6702;
      33985:data<=16'd5949;
      33986:data<=16'd6128;
      33987:data<=16'd5796;
      33988:data<=16'd5758;
      33989:data<=16'd6501;
      33990:data<=16'd6966;
      33991:data<=16'd6575;
      33992:data<=16'd6276;
      33993:data<=16'd5941;
      33994:data<=16'd5541;
      33995:data<=16'd6672;
      33996:data<=16'd7335;
      33997:data<=16'd6267;
      33998:data<=16'd5935;
      33999:data<=16'd5545;
      34000:data<=16'd5028;
      34001:data<=16'd5971;
      34002:data<=16'd6689;
      34003:data<=16'd6388;
      34004:data<=16'd5553;
      34005:data<=16'd5363;
      34006:data<=16'd5758;
      34007:data<=16'd4320;
      34008:data<=16'd5134;
      34009:data<=16'd9665;
      34010:data<=16'd10325;
      34011:data<=16'd8969;
      34012:data<=16'd9758;
      34013:data<=16'd8316;
      34014:data<=16'd6021;
      34015:data<=16'd5568;
      34016:data<=16'd4908;
      34017:data<=16'd4566;
      34018:data<=16'd4273;
      34019:data<=16'd3213;
      34020:data<=16'd1902;
      34021:data<=16'd531;
      34022:data<=16'd522;
      34023:data<=16'd717;
      34024:data<=16'd89;
      34025:data<=16'd305;
      34026:data<=-16'd775;
      34027:data<=-16'd2960;
      34028:data<=-16'd3121;
      34029:data<=-16'd3254;
      34030:data<=-16'd3563;
      34031:data<=-16'd2968;
      34032:data<=-16'd4144;
      34033:data<=-16'd6028;
      34034:data<=-16'd5909;
      34035:data<=-16'd5345;
      34036:data<=-16'd5470;
      34037:data<=-16'd5526;
      34038:data<=-16'd6015;
      34039:data<=-16'd7394;
      34040:data<=-16'd7931;
      34041:data<=-16'd7485;
      34042:data<=-16'd7645;
      34043:data<=-16'd7482;
      34044:data<=-16'd7430;
      34045:data<=-16'd8853;
      34046:data<=-16'd9588;
      34047:data<=-16'd9283;
      34048:data<=-16'd9062;
      34049:data<=-16'd8410;
      34050:data<=-16'd8308;
      34051:data<=-16'd9256;
      34052:data<=-16'd10437;
      34053:data<=-16'd10830;
      34054:data<=-16'd9890;
      34055:data<=-16'd9800;
      34056:data<=-16'd10026;
      34057:data<=-16'd9391;
      34058:data<=-16'd12087;
      34059:data<=-16'd16627;
      34060:data<=-16'd17570;
      34061:data<=-16'd16876;
      34062:data<=-16'd16524;
      34063:data<=-16'd16322;
      34064:data<=-16'd17051;
      34065:data<=-16'd17256;
      34066:data<=-16'd16587;
      34067:data<=-16'd15885;
      34068:data<=-16'd14863;
      34069:data<=-16'd14741;
      34070:data<=-16'd15700;
      34071:data<=-16'd16199;
      34072:data<=-16'd15822;
      34073:data<=-16'd15042;
      34074:data<=-16'd14446;
      34075:data<=-16'd13711;
      34076:data<=-16'd13740;
      34077:data<=-16'd15060;
      34078:data<=-16'd14619;
      34079:data<=-16'd13124;
      34080:data<=-16'd13068;
      34081:data<=-16'd12237;
      34082:data<=-16'd11646;
      34083:data<=-16'd12868;
      34084:data<=-16'd12812;
      34085:data<=-16'd12249;
      34086:data<=-16'd12452;
      34087:data<=-16'd11356;
      34088:data<=-16'd10642;
      34089:data<=-16'd11670;
      34090:data<=-16'd11953;
      34091:data<=-16'd11139;
      34092:data<=-16'd10757;
      34093:data<=-16'd10516;
      34094:data<=-16'd9800;
      34095:data<=-16'd10113;
      34096:data<=-16'd11144;
      34097:data<=-16'd10240;
      34098:data<=-16'd9250;
      34099:data<=-16'd9655;
      34100:data<=-16'd8725;
      34101:data<=-16'd8208;
      34102:data<=-16'd9429;
      34103:data<=-16'd9083;
      34104:data<=-16'd8399;
      34105:data<=-16'd8395;
      34106:data<=-16'd7348;
      34107:data<=-16'd7257;
      34108:data<=-16'd6381;
      34109:data<=-16'd1909;
      34110:data<=16'd989;
      34111:data<=16'd842;
      34112:data<=16'd1289;
      34113:data<=16'd1715;
      34114:data<=16'd2343;
      34115:data<=16'd3647;
      34116:data<=16'd3653;
      34117:data<=16'd3512;
      34118:data<=16'd3714;
      34119:data<=16'd3369;
      34120:data<=16'd4707;
      34121:data<=16'd6727;
      34122:data<=16'd6522;
      34123:data<=16'd6059;
      34124:data<=16'd6184;
      34125:data<=16'd5720;
      34126:data<=16'd6398;
      34127:data<=16'd8097;
      34128:data<=16'd8119;
      34129:data<=16'd7426;
      34130:data<=16'd7661;
      34131:data<=16'd7386;
      34132:data<=16'd7301;
      34133:data<=16'd8739;
      34134:data<=16'd9206;
      34135:data<=16'd8696;
      34136:data<=16'd9056;
      34137:data<=16'd8525;
      34138:data<=16'd7987;
      34139:data<=16'd9505;
      34140:data<=16'd10340;
      34141:data<=16'd9824;
      34142:data<=16'd9715;
      34143:data<=16'd9326;
      34144:data<=16'd8878;
      34145:data<=16'd9527;
      34146:data<=16'd10710;
      34147:data<=16'd10860;
      34148:data<=16'd9891;
      34149:data<=16'd9511;
      34150:data<=16'd9324;
      34151:data<=16'd9289;
      34152:data<=16'd10654;
      34153:data<=16'd10921;
      34154:data<=16'd10085;
      34155:data<=16'd10437;
      34156:data<=16'd9724;
      34157:data<=16'd9500;
      34158:data<=16'd10989;
      34159:data<=16'd8530;
      34160:data<=16'd4432;
      34161:data<=16'd4267;
      34162:data<=16'd4581;
      34163:data<=16'd4214;
      34164:data<=16'd5394;
      34165:data<=16'd6517;
      34166:data<=16'd6361;
      34167:data<=16'd5724;
      34168:data<=16'd5554;
      34169:data<=16'd5668;
      34170:data<=16'd5849;
      34171:data<=16'd6783;
      34172:data<=16'd7010;
      34173:data<=16'd6372;
      34174:data<=16'd6514;
      34175:data<=16'd6106;
      34176:data<=16'd6144;
      34177:data<=16'd7762;
      34178:data<=16'd7720;
      34179:data<=16'd7068;
      34180:data<=16'd7492;
      34181:data<=16'd6681;
      34182:data<=16'd6391;
      34183:data<=16'd7964;
      34184:data<=16'd8595;
      34185:data<=16'd8082;
      34186:data<=16'd7571;
      34187:data<=16'd7172;
      34188:data<=16'd6909;
      34189:data<=16'd7154;
      34190:data<=16'd8111;
      34191:data<=16'd8152;
      34192:data<=16'd7585;
      34193:data<=16'd7818;
      34194:data<=16'd7274;
      34195:data<=16'd7113;
      34196:data<=16'd8528;
      34197:data<=16'd8454;
      34198:data<=16'd7680;
      34199:data<=16'd7702;
      34200:data<=16'd7144;
      34201:data<=16'd7444;
      34202:data<=16'd8454;
      34203:data<=16'd8425;
      34204:data<=16'd8100;
      34205:data<=16'd7370;
      34206:data<=16'd7131;
      34207:data<=16'd7279;
      34208:data<=16'd6055;
      34209:data<=16'd7409;
      34210:data<=16'd11650;
      34211:data<=16'd12205;
      34212:data<=16'd10596;
      34213:data<=16'd10522;
      34214:data<=16'd9268;
      34215:data<=16'd7335;
      34216:data<=16'd7004;
      34217:data<=16'd6661;
      34218:data<=16'd5882;
      34219:data<=16'd5635;
      34220:data<=16'd4927;
      34221:data<=16'd3460;
      34222:data<=16'd2740;
      34223:data<=16'd2551;
      34224:data<=16'd2011;
      34225:data<=16'd1968;
      34226:data<=16'd1645;
      34227:data<=16'd68;
      34228:data<=-16'd840;
      34229:data<=-16'd913;
      34230:data<=-16'd1292;
      34231:data<=-16'd1262;
      34232:data<=-16'd1463;
      34233:data<=-16'd2922;
      34234:data<=-16'd4223;
      34235:data<=-16'd4114;
      34236:data<=-16'd3536;
      34237:data<=-16'd3750;
      34238:data<=-16'd4074;
      34239:data<=-16'd4514;
      34240:data<=-16'd5847;
      34241:data<=-16'd6134;
      34242:data<=-16'd5451;
      34243:data<=-16'd5805;
      34244:data<=-16'd5650;
      34245:data<=-16'd5604;
      34246:data<=-16'd7147;
      34247:data<=-16'd7494;
      34248:data<=-16'd6983;
      34249:data<=-16'd7106;
      34250:data<=-16'd6526;
      34251:data<=-16'd6793;
      34252:data<=-16'd8313;
      34253:data<=-16'd8834;
      34254:data<=-16'd8589;
      34255:data<=-16'd8085;
      34256:data<=-16'd8059;
      34257:data<=-16'd8305;
      34258:data<=-16'd8058;
      34259:data<=-16'd10768;
      34260:data<=-16'd15440;
      34261:data<=-16'd16333;
      34262:data<=-16'd15130;
      34263:data<=-16'd14439;
      34264:data<=-16'd14072;
      34265:data<=-16'd15198;
      34266:data<=-16'd15523;
      34267:data<=-16'd14421;
      34268:data<=-16'd14248;
      34269:data<=-16'd13289;
      34270:data<=-16'd12897;
      34271:data<=-16'd14660;
      34272:data<=-16'd14545;
      34273:data<=-16'd13579;
      34274:data<=-16'd13670;
      34275:data<=-16'd12304;
      34276:data<=-16'd11588;
      34277:data<=-16'd12921;
      34278:data<=-16'd13144;
      34279:data<=-16'd12413;
      34280:data<=-16'd12069;
      34281:data<=-16'd11453;
      34282:data<=-16'd10593;
      34283:data<=-16'd10757;
      34284:data<=-16'd11731;
      34285:data<=-16'd11286;
      34286:data<=-16'd10445;
      34287:data<=-16'd10665;
      34288:data<=-16'd9696;
      34289:data<=-16'd9065;
      34290:data<=-16'd10499;
      34291:data<=-16'd10625;
      34292:data<=-16'd9949;
      34293:data<=-16'd9881;
      34294:data<=-16'd8645;
      34295:data<=-16'd8363;
      34296:data<=-16'd9888;
      34297:data<=-16'd9817;
      34298:data<=-16'd8671;
      34299:data<=-16'd8357;
      34300:data<=-16'd7967;
      34301:data<=-16'd7720;
      34302:data<=-16'd8382;
      34303:data<=-16'd8569;
      34304:data<=-16'd8131;
      34305:data<=-16'd8169;
      34306:data<=-16'd7225;
      34307:data<=-16'd6156;
      34308:data<=-16'd6909;
      34309:data<=-16'd4848;
      34310:data<=16'd337;
      34311:data<=16'd1953;
      34312:data<=16'd1231;
      34313:data<=16'd1704;
      34314:data<=16'd2338;
      34315:data<=16'd3621;
      34316:data<=16'd4478;
      34317:data<=16'd4212;
      34318:data<=16'd4679;
      34319:data<=16'd4525;
      34320:data<=16'd4402;
      34321:data<=16'd6073;
      34322:data<=16'd6745;
      34323:data<=16'd6470;
      34324:data<=16'd6708;
      34325:data<=16'd6223;
      34326:data<=16'd6237;
      34327:data<=16'd7562;
      34328:data<=16'd8231;
      34329:data<=16'd7799;
      34330:data<=16'd7633;
      34331:data<=16'd8053;
      34332:data<=16'd7767;
      34333:data<=16'd7946;
      34334:data<=16'd9489;
      34335:data<=16'd9333;
      34336:data<=16'd8514;
      34337:data<=16'd9085;
      34338:data<=16'd8557;
      34339:data<=16'd8452;
      34340:data<=16'd9876;
      34341:data<=16'd9849;
      34342:data<=16'd9717;
      34343:data<=16'd9906;
      34344:data<=16'd8878;
      34345:data<=16'd9021;
      34346:data<=16'd10395;
      34347:data<=16'd10766;
      34348:data<=16'd10128;
      34349:data<=16'd9270;
      34350:data<=16'd9215;
      34351:data<=16'd9541;
      34352:data<=16'd10016;
      34353:data<=16'd10813;
      34354:data<=16'd10489;
      34355:data<=16'd10123;
      34356:data<=16'd9905;
      34357:data<=16'd8849;
      34358:data<=16'd10049;
      34359:data<=16'd10379;
      34360:data<=16'd5843;
      34361:data<=16'd3548;
      34362:data<=16'd4464;
      34363:data<=16'd3447;
      34364:data<=16'd3657;
      34365:data<=16'd5665;
      34366:data<=16'd5938;
      34367:data<=16'd5288;
      34368:data<=16'd4693;
      34369:data<=16'd4525;
      34370:data<=16'd4952;
      34371:data<=16'd5717;
      34372:data<=16'd6504;
      34373:data<=16'd5873;
      34374:data<=16'd5430;
      34375:data<=16'd5944;
      34376:data<=16'd4911;
      34377:data<=16'd5124;
      34378:data<=16'd7138;
      34379:data<=16'd6764;
      34380:data<=16'd6222;
      34381:data<=16'd6246;
      34382:data<=16'd4965;
      34383:data<=16'd5529;
      34384:data<=16'd7077;
      34385:data<=16'd6916;
      34386:data<=16'd6830;
      34387:data<=16'd6378;
      34388:data<=16'd5398;
      34389:data<=16'd5867;
      34390:data<=16'd7072;
      34391:data<=16'd7319;
      34392:data<=16'd6340;
      34393:data<=16'd5838;
      34394:data<=16'd6246;
      34395:data<=16'd6122;
      34396:data<=16'd6569;
      34397:data<=16'd7162;
      34398:data<=16'd6498;
      34399:data<=16'd6566;
      34400:data<=16'd6451;
      34401:data<=16'd5250;
      34402:data<=16'd5824;
      34403:data<=16'd7089;
      34404:data<=16'd6825;
      34405:data<=16'd6005;
      34406:data<=16'd5662;
      34407:data<=16'd5577;
      34408:data<=16'd4692;
      34409:data<=16'd5603;
      34410:data<=16'd9514;
      34411:data<=16'd10645;
      34412:data<=16'd9191;
      34413:data<=16'd9377;
      34414:data<=16'd8648;
      34415:data<=16'd6684;
      34416:data<=16'd5788;
      34417:data<=16'd5239;
      34418:data<=16'd4987;
      34419:data<=16'd4545;
      34420:data<=16'd3792;
      34421:data<=16'd3021;
      34422:data<=16'd1618;
      34423:data<=16'd1392;
      34424:data<=16'd1503;
      34425:data<=16'd232;
      34426:data<=16'd456;
      34427:data<=16'd297;
      34428:data<=-16'd1967;
      34429:data<=-16'd2167;
      34430:data<=-16'd1851;
      34431:data<=-16'd2717;
      34432:data<=-16'd2309;
      34433:data<=-16'd2749;
      34434:data<=-16'd4473;
      34435:data<=-16'd4992;
      34436:data<=-16'd5178;
      34437:data<=-16'd5124;
      34438:data<=-16'd4567;
      34439:data<=-16'd4907;
      34440:data<=-16'd6237;
      34441:data<=-16'd7159;
      34442:data<=-16'd6667;
      34443:data<=-16'd6343;
      34444:data<=-16'd6960;
      34445:data<=-16'd6995;
      34446:data<=-16'd7555;
      34447:data<=-16'd8631;
      34448:data<=-16'd8246;
      34449:data<=-16'd8088;
      34450:data<=-16'd8466;
      34451:data<=-16'd7914;
      34452:data<=-16'd8399;
      34453:data<=-16'd9946;
      34454:data<=-16'd9994;
      34455:data<=-16'd9307;
      34456:data<=-16'd9357;
      34457:data<=-16'd8939;
      34458:data<=-16'd8555;
      34459:data<=-16'd11373;
      34460:data<=-16'd15756;
      34461:data<=-16'd17020;
      34462:data<=-16'd16119;
      34463:data<=-16'd15714;
      34464:data<=-16'd15700;
      34465:data<=-16'd16225;
      34466:data<=-16'd16662;
      34467:data<=-16'd16073;
      34468:data<=-16'd15409;
      34469:data<=-16'd15017;
      34470:data<=-16'd14551;
      34471:data<=-16'd14845;
      34472:data<=-16'd15850;
      34473:data<=-16'd15720;
      34474:data<=-16'd14606;
      34475:data<=-16'd14099;
      34476:data<=-16'd13368;
      34477:data<=-16'd12988;
      34478:data<=-16'd14245;
      34479:data<=-16'd14202;
      34480:data<=-16'd12856;
      34481:data<=-16'd12722;
      34482:data<=-16'd11952;
      34483:data<=-16'd11474;
      34484:data<=-16'd13030;
      34485:data<=-16'd12877;
      34486:data<=-16'd11323;
      34487:data<=-16'd11441;
      34488:data<=-16'd11380;
      34489:data<=-16'd10689;
      34490:data<=-16'd11185;
      34491:data<=-16'd11759;
      34492:data<=-16'd11294;
      34493:data<=-16'd10851;
      34494:data<=-16'd10399;
      34495:data<=-16'd9279;
      34496:data<=-16'd9353;
      34497:data<=-16'd10678;
      34498:data<=-16'd10235;
      34499:data<=-16'd9148;
      34500:data<=-16'd9238;
      34501:data<=-16'd8730;
      34502:data<=-16'd8517;
      34503:data<=-16'd9488;
      34504:data<=-16'd9351;
      34505:data<=-16'd8595;
      34506:data<=-16'd8279;
      34507:data<=-16'd7676;
      34508:data<=-16'd7624;
      34509:data<=-16'd6740;
      34510:data<=-16'd2560;
      34511:data<=16'd1128;
      34512:data<=16'd1213;
      34513:data<=16'd978;
      34514:data<=16'd1491;
      34515:data<=16'd1929;
      34516:data<=16'd3274;
      34517:data<=16'd3862;
      34518:data<=16'd3530;
      34519:data<=16'd4199;
      34520:data<=16'd3952;
      34521:data<=16'd3896;
      34522:data<=16'd5908;
      34523:data<=16'd6278;
      34524:data<=16'd5832;
      34525:data<=16'd6554;
      34526:data<=16'd5817;
      34527:data<=16'd5796;
      34528:data<=16'd7664;
      34529:data<=16'd7832;
      34530:data<=16'd7327;
      34531:data<=16'd7423;
      34532:data<=16'd7013;
      34533:data<=16'd7272;
      34534:data<=16'd8481;
      34535:data<=16'd8948;
      34536:data<=16'd8225;
      34537:data<=16'd8091;
      34538:data<=16'd8765;
      34539:data<=16'd8208;
      34540:data<=16'd8272;
      34541:data<=16'd9823;
      34542:data<=16'd9652;
      34543:data<=16'd9148;
      34544:data<=16'd9356;
      34545:data<=16'd8314;
      34546:data<=16'd8607;
      34547:data<=16'd10516;
      34548:data<=16'd10458;
      34549:data<=16'd9480;
      34550:data<=16'd9259;
      34551:data<=16'd8963;
      34552:data<=16'd9182;
      34553:data<=16'd10502;
      34554:data<=16'd10991;
      34555:data<=16'd10140;
      34556:data<=16'd10022;
      34557:data<=16'd9765;
      34558:data<=16'd9488;
      34559:data<=16'd11066;
      34560:data<=16'd9488;
      34561:data<=16'd4408;
      34562:data<=16'd3668;
      34563:data<=16'd4705;
      34564:data<=16'd3419;
      34565:data<=16'd4217;
      34566:data<=16'd5930;
      34567:data<=16'd5592;
      34568:data<=16'd5278;
      34569:data<=16'd4901;
      34570:data<=16'd4232;
      34571:data<=16'd4969;
      34572:data<=16'd6496;
      34573:data<=16'd6633;
      34574:data<=16'd5650;
      34575:data<=16'd5510;
      34576:data<=16'd5482;
      34577:data<=16'd5518;
      34578:data<=16'd6956;
      34579:data<=16'd7306;
      34580:data<=16'd6319;
      34581:data<=16'd6370;
      34582:data<=16'd6052;
      34583:data<=16'd5685;
      34584:data<=16'd6746;
      34585:data<=16'd7488;
      34586:data<=16'd7335;
      34587:data<=16'd6836;
      34588:data<=16'd6155;
      34589:data<=16'd5658;
      34590:data<=16'd6043;
      34591:data<=16'd7533;
      34592:data<=16'd7780;
      34593:data<=16'd6883;
      34594:data<=16'd6868;
      34595:data<=16'd6222;
      34596:data<=16'd6358;
      34597:data<=16'd7994;
      34598:data<=16'd7571;
      34599:data<=16'd7209;
      34600:data<=16'd7608;
      34601:data<=16'd6414;
      34602:data<=16'd6758;
      34603:data<=16'd7677;
      34604:data<=16'd7141;
      34605:data<=16'd7494;
      34606:data<=16'd6928;
      34607:data<=16'd6217;
      34608:data<=16'd6660;
      34609:data<=16'd5348;
      34610:data<=16'd6780;
      34611:data<=16'd11482;
      34612:data<=16'd11588;
      34613:data<=16'd9824;
      34614:data<=16'd10334;
      34615:data<=16'd9342;
      34616:data<=16'd7172;
      34617:data<=16'd6382;
      34618:data<=16'd6270;
      34619:data<=16'd6202;
      34620:data<=16'd6216;
      34621:data<=16'd5363;
      34622:data<=16'd3366;
      34623:data<=16'd2596;
      34624:data<=16'd2910;
      34625:data<=16'd2159;
      34626:data<=16'd1898;
      34627:data<=16'd1729;
      34628:data<=16'd67;
      34629:data<=-16'd631;
      34630:data<=-16'd378;
      34631:data<=-16'd735;
      34632:data<=-16'd802;
      34633:data<=-16'd901;
      34634:data<=-16'd1871;
      34635:data<=-16'd3257;
      34636:data<=-16'd3553;
      34637:data<=-16'd2837;
      34638:data<=-16'd2952;
      34639:data<=-16'd2863;
      34640:data<=-16'd3200;
      34641:data<=-16'd5363;
      34642:data<=-16'd5557;
      34643:data<=-16'd4637;
      34644:data<=-16'd5312;
      34645:data<=-16'd4790;
      34646:data<=-16'd5109;
      34647:data<=-16'd7133;
      34648:data<=-16'd6754;
      34649:data<=-16'd6364;
      34650:data<=-16'd6934;
      34651:data<=-16'd6167;
      34652:data<=-16'd6367;
      34653:data<=-16'd7442;
      34654:data<=-16'd7859;
      34655:data<=-16'd7932;
      34656:data<=-16'd7303;
      34657:data<=-16'd7304;
      34658:data<=-16'd7100;
      34659:data<=-16'd6725;
      34660:data<=-16'd10546;
      34661:data<=-16'd14973;
      34662:data<=-16'd14812;
      34663:data<=-16'd13816;
      34664:data<=-16'd13549;
      34665:data<=-16'd13546;
      34666:data<=-16'd14841;
      34667:data<=-16'd14883;
      34668:data<=-16'd13671;
      34669:data<=-16'd13591;
      34670:data<=-16'd13209;
      34671:data<=-16'd12933;
      34672:data<=-16'd13850;
      34673:data<=-16'd13665;
      34674:data<=-16'd12668;
      34675:data<=-16'd12448;
      34676:data<=-16'd11846;
      34677:data<=-16'd11294;
      34678:data<=-16'd12069;
      34679:data<=-16'd12575;
      34680:data<=-16'd11997;
      34681:data<=-16'd11496;
      34682:data<=-16'd10915;
      34683:data<=-16'd10260;
      34684:data<=-16'd10780;
      34685:data<=-16'd11609;
      34686:data<=-16'd11056;
      34687:data<=-16'd10264;
      34688:data<=-16'd10043;
      34689:data<=-16'd9470;
      34690:data<=-16'd9517;
      34691:data<=-16'd10328;
      34692:data<=-16'd9894;
      34693:data<=-16'd9133;
      34694:data<=-16'd8987;
      34695:data<=-16'd8169;
      34696:data<=-16'd7965;
      34697:data<=-16'd9025;
      34698:data<=-16'd9276;
      34699:data<=-16'd8871;
      34700:data<=-16'd8370;
      34701:data<=-16'd7430;
      34702:data<=-16'd7288;
      34703:data<=-16'd8196;
      34704:data<=-16'd8564;
      34705:data<=-16'd8128;
      34706:data<=-16'd7649;
      34707:data<=-16'd6974;
      34708:data<=-16'd6699;
      34709:data<=-16'd7147;
      34710:data<=-16'd4714;
      34711:data<=16'd432;
      34712:data<=16'd2053;
      34713:data<=16'd989;
      34714:data<=16'd1513;
      34715:data<=16'd2419;
      34716:data<=16'd3674;
      34717:data<=16'd4751;
      34718:data<=16'd4070;
      34719:data<=16'd4173;
      34720:data<=16'd4790;
      34721:data<=16'd4686;
      34722:data<=16'd5858;
      34723:data<=16'd6575;
      34724:data<=16'd6049;
      34725:data<=16'd6537;
      34726:data<=16'd6617;
      34727:data<=16'd6044;
      34728:data<=16'd6865;
      34729:data<=16'd8135;
      34730:data<=16'd8220;
      34731:data<=16'd7765;
      34732:data<=16'd7844;
      34733:data<=16'd7577;
      34734:data<=16'd7709;
      34735:data<=16'd9530;
      34736:data<=16'd9817;
      34737:data<=16'd8819;
      34738:data<=16'd9289;
      34739:data<=16'd8801;
      34740:data<=16'd8616;
      34741:data<=16'd10481;
      34742:data<=16'd10592;
      34743:data<=16'd9914;
      34744:data<=16'd10035;
      34745:data<=16'd9298;
      34746:data<=16'd9179;
      34747:data<=16'd9962;
      34748:data<=16'd10746;
      34749:data<=16'd11153;
      34750:data<=16'd10187;
      34751:data<=16'd9474;
      34752:data<=16'd9380;
      34753:data<=16'd9700;
      34754:data<=16'd11271;
      34755:data<=16'd11195;
      34756:data<=16'd10191;
      34757:data<=16'd10404;
      34758:data<=16'd9756;
      34759:data<=16'd10709;
      34760:data<=16'd11638;
      34761:data<=16'd7830;
      34762:data<=16'd5765;
      34763:data<=16'd6940;
      34764:data<=16'd6185;
      34765:data<=16'd6206;
      34766:data<=16'd7215;
      34767:data<=16'd7063;
      34768:data<=16'd7232;
      34769:data<=16'd6898;
      34770:data<=16'd6223;
      34771:data<=16'd6276;
      34772:data<=16'd6942;
      34773:data<=16'd8122;
      34774:data<=16'd7661;
      34775:data<=16'd6745;
      34776:data<=16'd7130;
      34777:data<=16'd6548;
      34778:data<=16'd7065;
      34779:data<=16'd8772;
      34780:data<=16'd7935;
      34781:data<=16'd7368;
      34782:data<=16'd7570;
      34783:data<=16'd6428;
      34784:data<=16'd7031;
      34785:data<=16'd8316;
      34786:data<=16'd7514;
      34787:data<=16'd7069;
      34788:data<=16'd7294;
      34789:data<=16'd6780;
      34790:data<=16'd6686;
      34791:data<=16'd7524;
      34792:data<=16'd7712;
      34793:data<=16'd7060;
      34794:data<=16'd7086;
      34795:data<=16'd6793;
      34796:data<=16'd6120;
      34797:data<=16'd7174;
      34798:data<=16'd7659;
      34799:data<=16'd6563;
      34800:data<=16'd6739;
      34801:data<=16'd6810;
      34802:data<=16'd5874;
      34803:data<=16'd6269;
      34804:data<=16'd7092;
      34805:data<=16'd6677;
      34806:data<=16'd5952;
      34807:data<=16'd6085;
      34808:data<=16'd5985;
      34809:data<=16'd4686;
      34810:data<=16'd5175;
      34811:data<=16'd7971;
      34812:data<=16'd8986;
      34813:data<=16'd8069;
      34814:data<=16'd7424;
      34815:data<=16'd6845;
      34816:data<=16'd5723;
      34817:data<=16'd4153;
      34818:data<=16'd3287;
      34819:data<=16'd3319;
      34820:data<=16'd3172;
      34821:data<=16'd2892;
      34822:data<=16'd1642;
      34823:data<=-16'd379;
      34824:data<=-16'd705;
      34825:data<=-16'd325;
      34826:data<=-16'd741;
      34827:data<=-16'd864;
      34828:data<=-16'd1745;
      34829:data<=-16'd3582;
      34830:data<=-16'd4015;
      34831:data<=-16'd3659;
      34832:data<=-16'd3755;
      34833:data<=-16'd3642;
      34834:data<=-16'd4288;
      34835:data<=-16'd5965;
      34836:data<=-16'd6452;
      34837:data<=-16'd6031;
      34838:data<=-16'd6209;
      34839:data<=-16'd6085;
      34840:data<=-16'd6191;
      34841:data<=-16'd7692;
      34842:data<=-16'd8640;
      34843:data<=-16'd8338;
      34844:data<=-16'd8160;
      34845:data<=-16'd7841;
      34846:data<=-16'd7668;
      34847:data<=-16'd8812;
      34848:data<=-16'd10049;
      34849:data<=-16'd9788;
      34850:data<=-16'd9271;
      34851:data<=-16'd9414;
      34852:data<=-16'd8980;
      34853:data<=-16'd9047;
      34854:data<=-16'd10619;
      34855:data<=-16'd10649;
      34856:data<=-16'd9505;
      34857:data<=-16'd9997;
      34858:data<=-16'd9826;
      34859:data<=-16'd9091;
      34860:data<=-16'd11573;
      34861:data<=-16'd14985;
      34862:data<=-16'd15675;
      34863:data<=-16'd15064;
      34864:data<=-16'd14613;
      34865:data<=-16'd14402;
      34866:data<=-16'd15036;
      34867:data<=-16'd15643;
      34868:data<=-16'd14853;
      34869:data<=-16'd14137;
      34870:data<=-16'd14234;
      34871:data<=-16'd13576;
      34872:data<=-16'd13429;
      34873:data<=-16'd14439;
      34874:data<=-16'd14008;
      34875:data<=-16'd13174;
      34876:data<=-16'd13198;
      34877:data<=-16'd12345;
      34878:data<=-16'd12240;
      34879:data<=-16'd13364;
      34880:data<=-16'd12951;
      34881:data<=-16'd12366;
      34882:data<=-16'd12583;
      34883:data<=-16'd11702;
      34884:data<=-16'd11215;
      34885:data<=-16'd12248;
      34886:data<=-16'd12558;
      34887:data<=-16'd11825;
      34888:data<=-16'd11282;
      34889:data<=-16'd10854;
      34890:data<=-16'd10568;
      34891:data<=-16'd10975;
      34892:data<=-16'd11379;
      34893:data<=-16'd10840;
      34894:data<=-16'd10310;
      34895:data<=-16'd10032;
      34896:data<=-16'd9007;
      34897:data<=-16'd8928;
      34898:data<=-16'd10355;
      34899:data<=-16'd10137;
      34900:data<=-16'd9086;
      34901:data<=-16'd9400;
      34902:data<=-16'd8827;
      34903:data<=-16'd8284;
      34904:data<=-16'd9740;
      34905:data<=-16'd10006;
      34906:data<=-16'd9145;
      34907:data<=-16'd8884;
      34908:data<=-16'd7981;
      34909:data<=-16'd7897;
      34910:data<=-16'd7218;
      34911:data<=-16'd3253;
      34912:data<=-16'd1177;
      34913:data<=-16'd2015;
      34914:data<=-16'd1627;
      34915:data<=-16'd1327;
      34916:data<=-16'd526;
      34917:data<=16'd1459;
      34918:data<=16'd1527;
      34919:data<=16'd1454;
      34920:data<=16'd2126;
      34921:data<=16'd1671;
      34922:data<=16'd2540;
      34923:data<=16'd4196;
      34924:data<=16'd4094;
      34925:data<=16'd4226;
      34926:data<=16'd4666;
      34927:data<=16'd4275;
      34928:data<=16'd4731;
      34929:data<=16'd6075;
      34930:data<=16'd6575;
      34931:data<=16'd6378;
      34932:data<=16'd6467;
      34933:data<=16'd6228;
      34934:data<=16'd5955;
      34935:data<=16'd7253;
      34936:data<=16'd8352;
      34937:data<=16'd7858;
      34938:data<=16'd7808;
      34939:data<=16'd7806;
      34940:data<=16'd7257;
      34941:data<=16'd8052;
      34942:data<=16'd9371;
      34943:data<=16'd9348;
      34944:data<=16'd8951;
      34945:data<=16'd8883;
      34946:data<=16'd8222;
      34947:data<=16'd8135;
      34948:data<=16'd9814;
      34949:data<=16'd10251;
      34950:data<=16'd9250;
      34951:data<=16'd9583;
      34952:data<=16'd9226;
      34953:data<=16'd8580;
      34954:data<=16'd10210;
      34955:data<=16'd10928;
      34956:data<=16'd10248;
      34957:data<=16'd9962;
      34958:data<=16'd9144;
      34959:data<=16'd9404;
      34960:data<=16'd9674;
      34961:data<=16'd7441;
      34962:data<=16'd6034;
      34963:data<=16'd6272;
      34964:data<=16'd6117;
      34965:data<=16'd5900;
      34966:data<=16'd5900;
      34967:data<=16'd6736;
      34968:data<=16'd7288;
      34969:data<=16'd6689;
      34970:data<=16'd6734;
      34971:data<=16'd6435;
      34972:data<=16'd6322;
      34973:data<=16'd7903;
      34974:data<=16'd8035;
      34975:data<=16'd7303;
      34976:data<=16'd7403;
      34977:data<=16'd6482;
      34978:data<=16'd6599;
      34979:data<=16'd8152;
      34980:data<=16'd8199;
      34981:data<=16'd7585;
      34982:data<=16'd7122;
      34983:data<=16'd6892;
      34984:data<=16'd7124;
      34985:data<=16'd7300;
      34986:data<=16'd7865;
      34987:data<=16'd7723;
      34988:data<=16'd7022;
      34989:data<=16'd7250;
      34990:data<=16'd6522;
      34991:data<=16'd6197;
      34992:data<=16'd7689;
      34993:data<=16'd7632;
      34994:data<=16'd7210;
      34995:data<=16'd7356;
      34996:data<=16'd6170;
      34997:data<=16'd6373;
      34998:data<=16'd7802;
      34999:data<=16'd7744;
      35000:data<=16'd7374;
      35001:data<=16'd6717;
      35002:data<=16'd6058;
      35003:data<=16'd6569;
      35004:data<=16'd7204;
      35005:data<=16'd7348;
      35006:data<=16'd6828;
      35007:data<=16'd6569;
      35008:data<=16'd6780;
      35009:data<=16'd5714;
      35010:data<=16'd6006;
      35011:data<=16'd8827;
      35012:data<=16'd9600;
      35013:data<=16'd8522;
      35014:data<=16'd8313;
      35015:data<=16'd8213;
      35016:data<=16'd7250;
      35017:data<=16'd5468;
      35018:data<=16'd4502;
      35019:data<=16'd4262;
      35020:data<=16'd3284;
      35021:data<=16'd3213;
      35022:data<=16'd2984;
      35023:data<=16'd911;
      35024:data<=16'd56;
      35025:data<=16'd15;
      35026:data<=-16'd738;
      35027:data<=-16'd417;
      35028:data<=-16'd573;
      35029:data<=-16'd2343;
      35030:data<=-16'd3237;
      35031:data<=-16'd3028;
      35032:data<=-16'd3146;
      35033:data<=-16'd3612;
      35034:data<=-16'd3771;
      35035:data<=-16'd4416;
      35036:data<=-16'd5636;
      35037:data<=-16'd5448;
      35038:data<=-16'd5151;
      35039:data<=-16'd5783;
      35040:data<=-16'd5177;
      35041:data<=-16'd5441;
      35042:data<=-16'd7316;
      35043:data<=-16'd7483;
      35044:data<=-16'd7520;
      35045:data<=-16'd7985;
      35046:data<=-16'd6954;
      35047:data<=-16'd6927;
      35048:data<=-16'd8276;
      35049:data<=-16'd8734;
      35050:data<=-16'd8640;
      35051:data<=-16'd8340;
      35052:data<=-16'd8150;
      35053:data<=-16'd8293;
      35054:data<=-16'd8795;
      35055:data<=-16'd9603;
      35056:data<=-16'd9247;
      35057:data<=-16'd9056;
      35058:data<=-16'd9715;
      35059:data<=-16'd8560;
      35060:data<=-16'd9345;
      35061:data<=-16'd13759;
      35062:data<=-16'd14956;
      35063:data<=-16'd13955;
      35064:data<=-16'd14539;
      35065:data<=-16'd13829;
      35066:data<=-16'd13273;
      35067:data<=-16'd14380;
      35068:data<=-16'd14161;
      35069:data<=-16'd13644;
      35070:data<=-16'd13511;
      35071:data<=-16'd12416;
      35072:data<=-16'd12198;
      35073:data<=-16'd13107;
      35074:data<=-16'd13185;
      35075:data<=-16'd12569;
      35076:data<=-16'd12132;
      35077:data<=-16'd11835;
      35078:data<=-16'd11300;
      35079:data<=-16'd11251;
      35080:data<=-16'd11964;
      35081:data<=-16'd11928;
      35082:data<=-16'd11386;
      35083:data<=-16'd10974;
      35084:data<=-16'd9897;
      35085:data<=-16'd9667;
      35086:data<=-16'd10969;
      35087:data<=-16'd11257;
      35088:data<=-16'd10493;
      35089:data<=-16'd10035;
      35090:data<=-16'd9309;
      35091:data<=-16'd9085;
      35092:data<=-16'd10170;
      35093:data<=-16'd10451;
      35094:data<=-16'd9555;
      35095:data<=-16'd9183;
      35096:data<=-16'd8549;
      35097:data<=-16'd7987;
      35098:data<=-16'd9162;
      35099:data<=-16'd9706;
      35100:data<=-16'd8819;
      35101:data<=-16'd8742;
      35102:data<=-16'd8184;
      35103:data<=-16'd7075;
      35104:data<=-16'd7538;
      35105:data<=-16'd8320;
      35106:data<=-16'd8436;
      35107:data<=-16'd7744;
      35108:data<=-16'd6593;
      35109:data<=-16'd6643;
      35110:data<=-16'd5353;
      35111:data<=-16'd1844;
      35112:data<=-16'd641;
      35113:data<=-16'd628;
      35114:data<=16'd393;
      35115:data<=16'd279;
      35116:data<=16'd560;
      35117:data<=16'd2106;
      35118:data<=16'd2743;
      35119:data<=16'd3113;
      35120:data<=16'd3338;
      35121:data<=16'd3005;
      35122:data<=16'd3401;
      35123:data<=16'd4551;
      35124:data<=16'd5621;
      35125:data<=16'd5888;
      35126:data<=16'd5762;
      35127:data<=16'd5984;
      35128:data<=16'd5739;
      35129:data<=16'd6081;
      35130:data<=16'd7454;
      35131:data<=16'd7694;
      35132:data<=16'd7780;
      35133:data<=16'd8052;
      35134:data<=16'd7359;
      35135:data<=16'd8075;
      35136:data<=16'd9605;
      35137:data<=16'd9521;
      35138:data<=16'd9468;
      35139:data<=16'd9383;
      35140:data<=16'd8672;
      35141:data<=16'd9186;
      35142:data<=16'd10343;
      35143:data<=16'd10595;
      35144:data<=16'd10269;
      35145:data<=16'd10056;
      35146:data<=16'd9966;
      35147:data<=16'd9828;
      35148:data<=16'd10449;
      35149:data<=16'd11274;
      35150:data<=16'd11048;
      35151:data<=16'd10901;
      35152:data<=16'd10786;
      35153:data<=16'd10196;
      35154:data<=16'd10572;
      35155:data<=16'd11354;
      35156:data<=16'd11438;
      35157:data<=16'd11174;
      35158:data<=16'd10769;
      35159:data<=16'd10610;
      35160:data<=16'd9732;
      35161:data<=16'd8067;
      35162:data<=16'd7671;
      35163:data<=16'd7711;
      35164:data<=16'd7163;
      35165:data<=16'd6946;
      35166:data<=16'd7078;
      35167:data<=16'd8119;
      35168:data<=16'd8898;
      35169:data<=16'd7968;
      35170:data<=16'd7791;
      35171:data<=16'd8093;
      35172:data<=16'd7291;
      35173:data<=16'd7824;
      35174:data<=16'd9147;
      35175:data<=16'd9019;
      35176:data<=16'd8775;
      35177:data<=16'd8570;
      35178:data<=16'd7802;
      35179:data<=16'd8158;
      35180:data<=16'd9756;
      35181:data<=16'd10023;
      35182:data<=16'd8687;
      35183:data<=16'd8035;
      35184:data<=16'd7979;
      35185:data<=16'd8140;
      35186:data<=16'd9385;
      35187:data<=16'd9720;
      35188:data<=16'd8668;
      35189:data<=16'd8454;
      35190:data<=16'd8119;
      35191:data<=16'd7723;
      35192:data<=16'd8763;
      35193:data<=16'd9277;
      35194:data<=16'd8766;
      35195:data<=16'd8680;
      35196:data<=16'd8161;
      35197:data<=16'd7106;
      35198:data<=16'd7417;
      35199:data<=16'd8898;
      35200:data<=16'd8956;
      35201:data<=16'd7991;
      35202:data<=16'd7870;
      35203:data<=16'd7144;
      35204:data<=16'd6942;
      35205:data<=16'd8748;
      35206:data<=16'd8664;
      35207:data<=16'd7420;
      35208:data<=16'd7567;
      35209:data<=16'd6708;
      35210:data<=16'd7342;
      35211:data<=16'd10446;
      35212:data<=16'd10480;
      35213:data<=16'd8983;
      35214:data<=16'd9091;
      35215:data<=16'd8677;
      35216:data<=16'd7720;
      35217:data<=16'd6322;
      35218:data<=16'd4848;
      35219:data<=16'd4764;
      35220:data<=16'd4290;
      35221:data<=16'd3450;
      35222:data<=16'd3557;
      35223:data<=16'd2535;
      35224:data<=16'd878;
      35225:data<=16'd391;
      35226:data<=-16'd123;
      35227:data<=-16'd513;
      35228:data<=-16'd305;
      35229:data<=-16'd1227;
      35230:data<=-16'd2936;
      35231:data<=-16'd3298;
      35232:data<=-16'd3113;
      35233:data<=-16'd3620;
      35234:data<=-16'd3588;
      35235:data<=-16'd3830;
      35236:data<=-16'd5404;
      35237:data<=-16'd5923;
      35238:data<=-16'd5594;
      35239:data<=-16'd6017;
      35240:data<=-16'd5934;
      35241:data<=-16'd5947;
      35242:data<=-16'd6912;
      35243:data<=-16'd7562;
      35244:data<=-16'd7967;
      35245:data<=-16'd8205;
      35246:data<=-16'd7984;
      35247:data<=-16'd7595;
      35248:data<=-16'd7650;
      35249:data<=-16'd9018;
      35250:data<=-16'd9802;
      35251:data<=-16'd8951;
      35252:data<=-16'd8657;
      35253:data<=-16'd8376;
      35254:data<=-16'd8517;
      35255:data<=-16'd10272;
      35256:data<=-16'd10475;
      35257:data<=-16'd9732;
      35258:data<=-16'd9770;
      35259:data<=-16'd8818;
      35260:data<=-16'd10326;
      35261:data<=-16'd14781;
      35262:data<=-16'd16014;
      35263:data<=-16'd15089;
      35264:data<=-16'd15185;
      35265:data<=-16'd14792;
      35266:data<=-16'd14099;
      35267:data<=-16'd14189;
      35268:data<=-16'd14865;
      35269:data<=-16'd15092;
      35270:data<=-16'd14354;
      35271:data<=-16'd13668;
      35272:data<=-16'd12936;
      35273:data<=-16'd12957;
      35274:data<=-16'd14416;
      35275:data<=-16'd14546;
      35276:data<=-16'd13562;
      35277:data<=-16'd13051;
      35278:data<=-16'd12011;
      35279:data<=-16'd12066;
      35280:data<=-16'd13382;
      35281:data<=-16'd13364;
      35282:data<=-16'd12754;
      35283:data<=-16'd12082;
      35284:data<=-16'd11173;
      35285:data<=-16'd11210;
      35286:data<=-16'd11987;
      35287:data<=-16'd12633;
      35288:data<=-16'd12208;
      35289:data<=-16'd11110;
      35290:data<=-16'd10554;
      35291:data<=-16'd9758;
      35292:data<=-16'd10003;
      35293:data<=-16'd11605;
      35294:data<=-16'd11119;
      35295:data<=-16'd9940;
      35296:data<=-16'd9749;
      35297:data<=-16'd8866;
      35298:data<=-16'd9256;
      35299:data<=-16'd10602;
      35300:data<=-16'd10187;
      35301:data<=-16'd9559;
      35302:data<=-16'd9062;
      35303:data<=-16'd8355;
      35304:data<=-16'd8731;
      35305:data<=-16'd9515;
      35306:data<=-16'd9826;
      35307:data<=-16'd9080;
      35308:data<=-16'd8160;
      35309:data<=-16'd8411;
      35310:data<=-16'd6758;
      35311:data<=-16'd3066;
      35312:data<=-16'd1856;
      35313:data<=-16'd2130;
      35314:data<=-16'd1328;
      35315:data<=-16'd875;
      35316:data<=-16'd1233;
      35317:data<=-16'd690;
      35318:data<=16'd923;
      35319:data<=16'd1486;
      35320:data<=16'd1401;
      35321:data<=16'd2033;
      35322:data<=16'd1824;
      35323:data<=16'd2258;
      35324:data<=16'd4397;
      35325:data<=16'd4670;
      35326:data<=16'd4252;
      35327:data<=16'd4884;
      35328:data<=16'd4405;
      35329:data<=16'd4579;
      35330:data<=16'd6058;
      35331:data<=16'd6458;
      35332:data<=16'd6481;
      35333:data<=16'd6373;
      35334:data<=16'd6123;
      35335:data<=16'd6540;
      35336:data<=16'd7063;
      35337:data<=16'd7827;
      35338:data<=16'd8187;
      35339:data<=16'd7699;
      35340:data<=16'd7589;
      35341:data<=16'd7244;
      35342:data<=16'd7592;
      35343:data<=16'd9298;
      35344:data<=16'd9274;
      35345:data<=16'd8352;
      35346:data<=16'd8223;
      35347:data<=16'd7729;
      35348:data<=16'd8449;
      35349:data<=16'd9765;
      35350:data<=16'd9386;
      35351:data<=16'd8960;
      35352:data<=16'd8616;
      35353:data<=16'd8128;
      35354:data<=16'd8856;
      35355:data<=16'd9828;
      35356:data<=16'd10263;
      35357:data<=16'd9950;
      35358:data<=16'd9459;
      35359:data<=16'd9724;
      35360:data<=16'd8043;
      35361:data<=16'd5432;
      35362:data<=16'd6228;
      35363:data<=16'd7316;
      35364:data<=16'd6590;
      35365:data<=16'd6561;
      35366:data<=16'd6285;
      35367:data<=16'd6461;
      35368:data<=16'd8017;
      35369:data<=16'd8055;
      35370:data<=16'd7507;
      35371:data<=16'd7671;
      35372:data<=16'd7030;
      35373:data<=16'd7310;
      35374:data<=16'd8731;
      35375:data<=16'd8774;
      35376:data<=16'd8246;
      35377:data<=16'd8046;
      35378:data<=16'd7523;
      35379:data<=16'd7429;
      35380:data<=16'd8458;
      35381:data<=16'd9471;
      35382:data<=16'd9191;
      35383:data<=16'd8578;
      35384:data<=16'd8261;
      35385:data<=16'd7545;
      35386:data<=16'd8146;
      35387:data<=16'd9894;
      35388:data<=16'd9677;
      35389:data<=16'd8839;
      35390:data<=16'd8713;
      35391:data<=16'd7841;
      35392:data<=16'd7993;
      35393:data<=16'd9368;
      35394:data<=16'd9398;
      35395:data<=16'd9128;
      35396:data<=16'd9153;
      35397:data<=16'd8319;
      35398:data<=16'd8078;
      35399:data<=16'd9062;
      35400:data<=16'd9395;
      35401:data<=16'd8812;
      35402:data<=16'd8381;
      35403:data<=16'd7764;
      35404:data<=16'd7198;
      35405:data<=16'd7905;
      35406:data<=16'd8627;
      35407:data<=16'd8354;
      35408:data<=16'd7827;
      35409:data<=16'd6852;
      35410:data<=16'd7500;
      35411:data<=16'd10272;
      35412:data<=16'd10584;
      35413:data<=16'd9057;
      35414:data<=16'd8760;
      35415:data<=16'd8294;
      35416:data<=16'd7937;
      35417:data<=16'd7045;
      35418:data<=16'd4642;
      35419:data<=16'd4085;
      35420:data<=16'd4364;
      35421:data<=16'd3331;
      35422:data<=16'd3281;
      35423:data<=16'd2623;
      35424:data<=16'd641;
      35425:data<=16'd256;
      35426:data<=16'd144;
      35427:data<=-16'd553;
      35428:data<=-16'd526;
      35429:data<=-16'd826;
      35430:data<=-16'd2076;
      35431:data<=-16'd3469;
      35432:data<=-16'd3982;
      35433:data<=-16'd3824;
      35434:data<=-16'd3983;
      35435:data<=-16'd3874;
      35436:data<=-16'd4441;
      35437:data<=-16'd6203;
      35438:data<=-16'd6614;
      35439:data<=-16'd6272;
      35440:data<=-16'd6285;
      35441:data<=-16'd5741;
      35442:data<=-16'd6526;
      35443:data<=-16'd8358;
      35444:data<=-16'd8449;
      35445:data<=-16'd7971;
      35446:data<=-16'd8031;
      35447:data<=-16'd7823;
      35448:data<=-16'd8026;
      35449:data<=-16'd9169;
      35450:data<=-16'd9979;
      35451:data<=-16'd9659;
      35452:data<=-16'd9552;
      35453:data<=-16'd9664;
      35454:data<=-16'd9028;
      35455:data<=-16'd9524;
      35456:data<=-16'd10992;
      35457:data<=-16'd10988;
      35458:data<=-16'd10216;
      35459:data<=-16'd9579;
      35460:data<=-16'd10369;
      35461:data<=-16'd13758;
      35462:data<=-16'd16031;
      35463:data<=-16'd15424;
      35464:data<=-16'd14847;
      35465:data<=-16'd14580;
      35466:data<=-16'd13932;
      35467:data<=-16'd13940;
      35468:data<=-16'd14751;
      35469:data<=-16'd15059;
      35470:data<=-16'd14216;
      35471:data<=-16'd13743;
      35472:data<=-16'd13735;
      35473:data<=-16'd13076;
      35474:data<=-16'd13514;
      35475:data<=-16'd14744;
      35476:data<=-16'd14108;
      35477:data<=-16'd13038;
      35478:data<=-16'd12797;
      35479:data<=-16'd12196;
      35480:data<=-16'd12346;
      35481:data<=-16'd13565;
      35482:data<=-16'd13361;
      35483:data<=-16'd12141;
      35484:data<=-16'd11887;
      35485:data<=-16'd11492;
      35486:data<=-16'd11209;
      35487:data<=-16'd12346;
      35488:data<=-16'd12299;
      35489:data<=-16'd10991;
      35490:data<=-16'd11047;
      35491:data<=-16'd10648;
      35492:data<=-16'd9919;
      35493:data<=-16'd11050;
      35494:data<=-16'd11502;
      35495:data<=-16'd10455;
      35496:data<=-16'd9756;
      35497:data<=-16'd9144;
      35498:data<=-16'd8968;
      35499:data<=-16'd9597;
      35500:data<=-16'd10147;
      35501:data<=-16'd9787;
      35502:data<=-16'd8765;
      35503:data<=-16'd8519;
      35504:data<=-16'd8211;
      35505:data<=-16'd7820;
      35506:data<=-16'd9125;
      35507:data<=-16'd9125;
      35508:data<=-16'd7683;
      35509:data<=-16'd8167;
      35510:data<=-16'd6487;
      35511:data<=-16'd2161;
      35512:data<=-16'd1099;
      35513:data<=-16'd1632;
      35514:data<=-16'd1039;
      35515:data<=-16'd926;
      35516:data<=-16'd839;
      35517:data<=-16'd50;
      35518:data<=16'd1148;
      35519:data<=16'd2005;
      35520:data<=16'd2109;
      35521:data<=16'd2664;
      35522:data<=16'd2946;
      35523:data<=16'd2569;
      35524:data<=16'd3697;
      35525:data<=16'd5297;
      35526:data<=16'd5474;
      35527:data<=16'd5363;
      35528:data<=16'd5280;
      35529:data<=16'd5022;
      35530:data<=16'd5839;
      35531:data<=16'd7467;
      35532:data<=16'd7817;
      35533:data<=16'd7332;
      35534:data<=16'd7503;
      35535:data<=16'd7451;
      35536:data<=16'd7749;
      35537:data<=16'd8849;
      35538:data<=16'd8690;
      35539:data<=16'd8552;
      35540:data<=16'd9195;
      35541:data<=16'd8470;
      35542:data<=16'd8272;
      35543:data<=16'd9497;
      35544:data<=16'd9958;
      35545:data<=16'd9923;
      35546:data<=16'd9435;
      35547:data<=16'd8912;
      35548:data<=16'd9081;
      35549:data<=16'd9244;
      35550:data<=16'd10416;
      35551:data<=16'd11136;
      35552:data<=16'd9797;
      35553:data<=16'd9717;
      35554:data<=16'd10125;
      35555:data<=16'd9794;
      35556:data<=16'd11039;
      35557:data<=16'd11109;
      35558:data<=16'd10066;
      35559:data<=16'd10821;
      35560:data<=16'd9342;
      35561:data<=16'd6384;
      35562:data<=16'd6887;
      35563:data<=16'd8008;
      35564:data<=16'd7614;
      35565:data<=16'd7388;
      35566:data<=16'd7012;
      35567:data<=16'd6673;
      35568:data<=16'd7389;
      35569:data<=16'd8561;
      35570:data<=16'd8572;
      35571:data<=16'd7743;
      35572:data<=16'd7688;
      35573:data<=16'd7536;
      35574:data<=16'd7551;
      35575:data<=16'd8833;
      35576:data<=16'd8950;
      35577:data<=16'd8294;
      35578:data<=16'd8652;
      35579:data<=16'd7985;
      35580:data<=16'd7743;
      35581:data<=16'd9468;
      35582:data<=16'd9723;
      35583:data<=16'd8903;
      35584:data<=16'd8942;
      35585:data<=16'd8307;
      35586:data<=16'd7997;
      35587:data<=16'd9465;
      35588:data<=16'd10313;
      35589:data<=16'd9166;
      35590:data<=16'd8070;
      35591:data<=16'd8134;
      35592:data<=16'd8173;
      35593:data<=16'd8827;
      35594:data<=16'd10117;
      35595:data<=16'd9407;
      35596:data<=16'd8487;
      35597:data<=16'd9097;
      35598:data<=16'd8392;
      35599:data<=16'd8296;
      35600:data<=16'd9876;
      35601:data<=16'd9175;
      35602:data<=16'd8332;
      35603:data<=16'd8733;
      35604:data<=16'd7539;
      35605:data<=16'd7430;
      35606:data<=16'd8921;
      35607:data<=16'd9018;
      35608:data<=16'd8567;
      35609:data<=16'd7706;
      35610:data<=16'd8020;
      35611:data<=16'd10713;
      35612:data<=16'd11311;
      35613:data<=16'd10066;
      35614:data<=16'd9814;
      35615:data<=16'd8790;
      35616:data<=16'd8096;
      35617:data<=16'd8322;
      35618:data<=16'd6886;
      35619:data<=16'd5068;
      35620:data<=16'd4375;
      35621:data<=16'd4149;
      35622:data<=16'd4199;
      35623:data<=16'd3917;
      35624:data<=16'd2833;
      35625:data<=16'd1290;
      35626:data<=16'd728;
      35627:data<=16'd1137;
      35628:data<=16'd669;
      35629:data<=16'd230;
      35630:data<=-16'd415;
      35631:data<=-16'd2350;
      35632:data<=-16'd2796;
      35633:data<=-16'd2602;
      35634:data<=-16'd3363;
      35635:data<=-16'd2707;
      35636:data<=-16'd2743;
      35637:data<=-16'd4440;
      35638:data<=-16'd4778;
      35639:data<=-16'd4919;
      35640:data<=-16'd5180;
      35641:data<=-16'd4645;
      35642:data<=-16'd4705;
      35643:data<=-16'd5462;
      35644:data<=-16'd6734;
      35645:data<=-16'd7188;
      35646:data<=-16'd6493;
      35647:data<=-16'd6866;
      35648:data<=-16'd6880;
      35649:data<=-16'd6893;
      35650:data<=-16'd8407;
      35651:data<=-16'd8044;
      35652:data<=-16'd7391;
      35653:data<=-16'd8153;
      35654:data<=-16'd7306;
      35655:data<=-16'd7615;
      35656:data<=-16'd9298;
      35657:data<=-16'd9135;
      35658:data<=-16'd9323;
      35659:data<=-16'd9200;
      35660:data<=-16'd9166;
      35661:data<=-16'd12266;
      35662:data<=-16'd14533;
      35663:data<=-16'd14424;
      35664:data<=-16'd14193;
      35665:data<=-16'd13239;
      35666:data<=-16'd12842;
      35667:data<=-16'd12938;
      35668:data<=-16'd12783;
      35669:data<=-16'd13649;
      35670:data<=-16'd13609;
      35671:data<=-16'd12901;
      35672:data<=-16'd13035;
      35673:data<=-16'd12047;
      35674:data<=-16'd11765;
      35675:data<=-16'd13053;
      35676:data<=-16'd12868;
      35677:data<=-16'd12458;
      35678:data<=-16'd12546;
      35679:data<=-16'd11646;
      35680:data<=-16'd11365;
      35681:data<=-16'd12434;
      35682:data<=-16'd13032;
      35683:data<=-16'd12302;
      35684:data<=-16'd11593;
      35685:data<=-16'd11606;
      35686:data<=-16'd11244;
      35687:data<=-16'd11414;
      35688:data<=-16'd12205;
      35689:data<=-16'd11652;
      35690:data<=-16'd11045;
      35691:data<=-16'd10809;
      35692:data<=-16'd9799;
      35693:data<=-16'd9902;
      35694:data<=-16'd10787;
      35695:data<=-16'd10490;
      35696:data<=-16'd9990;
      35697:data<=-16'd9456;
      35698:data<=-16'd8604;
      35699:data<=-16'd8798;
      35700:data<=-16'd9976;
      35701:data<=-16'd10161;
      35702:data<=-16'd9315;
      35703:data<=-16'd8980;
      35704:data<=-16'd8223;
      35705:data<=-16'd7649;
      35706:data<=-16'd9257;
      35707:data<=-16'd9473;
      35708:data<=-16'd7894;
      35709:data<=-16'd8225;
      35710:data<=-16'd6683;
      35711:data<=-16'd2867;
      35712:data<=-16'd2344;
      35713:data<=-16'd2787;
      35714:data<=-16'd1914;
      35715:data<=-16'd1823;
      35716:data<=-16'd1618;
      35717:data<=-16'd1069;
      35718:data<=-16'd224;
      35719:data<=16'd1165;
      35720:data<=16'd1441;
      35721:data<=16'd1621;
      35722:data<=16'd2232;
      35723:data<=16'd1991;
      35724:data<=16'd2673;
      35725:data<=16'd3899;
      35726:data<=16'd4006;
      35727:data<=16'd4619;
      35728:data<=16'd5139;
      35729:data<=16'd4444;
      35730:data<=16'd4587;
      35731:data<=16'd6014;
      35732:data<=16'd7016;
      35733:data<=16'd6854;
      35734:data<=16'd6328;
      35735:data<=16'd6050;
      35736:data<=16'd5984;
      35737:data<=16'd6786;
      35738:data<=16'd7711;
      35739:data<=16'd7511;
      35740:data<=16'd7407;
      35741:data<=16'd7447;
      35742:data<=16'd6943;
      35743:data<=16'd7244;
      35744:data<=16'd7935;
      35745:data<=16'd7850;
      35746:data<=16'd7817;
      35747:data<=16'd7702;
      35748:data<=16'd7121;
      35749:data<=16'd7353;
      35750:data<=16'd8540;
      35751:data<=16'd9085;
      35752:data<=16'd8853;
      35753:data<=16'd8651;
      35754:data<=16'd8002;
      35755:data<=16'd7932;
      35756:data<=16'd9476;
      35757:data<=16'd9767;
      35758:data<=16'd8630;
      35759:data<=16'd8762;
      35760:data<=16'd7574;
      35761:data<=16'd4276;
      35762:data<=16'd3968;
      35763:data<=16'd6068;
      35764:data<=16'd6155;
      35765:data<=16'd5685;
      35766:data<=16'd6222;
      35767:data<=16'd5741;
      35768:data<=16'd5432;
      35769:data<=16'd6874;
      35770:data<=16'd7379;
      35771:data<=16'd6717;
      35772:data<=16'd6567;
      35773:data<=16'd5767;
      35774:data<=16'd5588;
      35775:data<=16'd7304;
      35776:data<=16'd7689;
      35777:data<=16'd6831;
      35778:data<=16'd6980;
      35779:data<=16'd6749;
      35780:data<=16'd6091;
      35781:data<=16'd6470;
      35782:data<=16'd7141;
      35783:data<=16'd7263;
      35784:data<=16'd7219;
      35785:data<=16'd7160;
      35786:data<=16'd6534;
      35787:data<=16'd6516;
      35788:data<=16'd8012;
      35789:data<=16'd8140;
      35790:data<=16'd7086;
      35791:data<=16'd7407;
      35792:data<=16'd6936;
      35793:data<=16'd6328;
      35794:data<=16'd8025;
      35795:data<=16'd8560;
      35796:data<=16'd7482;
      35797:data<=16'd7272;
      35798:data<=16'd6798;
      35799:data<=16'd6716;
      35800:data<=16'd7498;
      35801:data<=16'd7342;
      35802:data<=16'd7086;
      35803:data<=16'd6995;
      35804:data<=16'd6228;
      35805:data<=16'd5799;
      35806:data<=16'd6302;
      35807:data<=16'd7277;
      35808:data<=16'd7250;
      35809:data<=16'd6487;
      35810:data<=16'd7859;
      35811:data<=16'd9873;
      35812:data<=16'd9609;
      35813:data<=16'd8980;
      35814:data<=16'd8892;
      35815:data<=16'd7997;
      35816:data<=16'd6828;
      35817:data<=16'd6443;
      35818:data<=16'd6213;
      35819:data<=16'd4631;
      35820:data<=16'd3037;
      35821:data<=16'd3195;
      35822:data<=16'd2913;
      35823:data<=16'd2120;
      35824:data<=16'd2262;
      35825:data<=16'd983;
      35826:data<=-16'd740;
      35827:data<=-16'd255;
      35828:data<=-16'd399;
      35829:data<=-16'd1507;
      35830:data<=-16'd1052;
      35831:data<=-16'd1290;
      35832:data<=-16'd3281;
      35833:data<=-16'd4135;
      35834:data<=-16'd3876;
      35835:data<=-16'd4014;
      35836:data<=-16'd4162;
      35837:data<=-16'd4819;
      35838:data<=-16'd6229;
      35839:data<=-16'd6673;
      35840:data<=-16'd6573;
      35841:data<=-16'd6990;
      35842:data<=-16'd6495;
      35843:data<=-16'd6214;
      35844:data<=-16'd7935;
      35845:data<=-16'd8846;
      35846:data<=-16'd8072;
      35847:data<=-16'd8172;
      35848:data<=-16'd8704;
      35849:data<=-16'd8602;
      35850:data<=-16'd8916;
      35851:data<=-16'd9494;
      35852:data<=-16'd9312;
      35853:data<=-16'd9122;
      35854:data<=-16'd9482;
      35855:data<=-16'd9323;
      35856:data<=-16'd9468;
      35857:data<=-16'd10642;
      35858:data<=-16'd10405;
      35859:data<=-16'd9903;
      35860:data<=-16'd11844;
      35861:data<=-16'd13470;
      35862:data<=-16'd14098;
      35863:data<=-16'd15540;
      35864:data<=-16'd15869;
      35865:data<=-16'd15092;
      35866:data<=-16'd14474;
      35867:data<=-16'd13392;
      35868:data<=-16'd13321;
      35869:data<=-16'd14155;
      35870:data<=-16'd14214;
      35871:data<=-16'd14537;
      35872:data<=-16'd14769;
      35873:data<=-16'd13996;
      35874:data<=-16'd13294;
      35875:data<=-16'd13221;
      35876:data<=-16'd13897;
      35877:data<=-16'd14125;
      35878:data<=-16'd13389;
      35879:data<=-16'd13074;
      35880:data<=-16'd12452;
      35881:data<=-16'd12146;
      35882:data<=-16'd13267;
      35883:data<=-16'd13168;
      35884:data<=-16'd12490;
      35885:data<=-16'd12596;
      35886:data<=-16'd11506;
      35887:data<=-16'd11232;
      35888:data<=-16'd12349;
      35889:data<=-16'd11879;
      35890:data<=-16'd11374;
      35891:data<=-16'd11233;
      35892:data<=-16'd10069;
      35893:data<=-16'd10002;
      35894:data<=-16'd10769;
      35895:data<=-16'd10540;
      35896:data<=-16'd10170;
      35897:data<=-16'd9909;
      35898:data<=-16'd9194;
      35899:data<=-16'd8496;
      35900:data<=-16'd9028;
      35901:data<=-16'd10144;
      35902:data<=-16'd9823;
      35903:data<=-16'd8956;
      35904:data<=-16'd8167;
      35905:data<=-16'd7128;
      35906:data<=-16'd7805;
      35907:data<=-16'd8936;
      35908:data<=-16'd8282;
      35909:data<=-16'd7382;
      35910:data<=-16'd5362;
      35911:data<=-16'd2381;
      35912:data<=-16'd1859;
      35913:data<=-16'd2302;
      35914:data<=-16'd1579;
      35915:data<=-16'd1283;
      35916:data<=-16'd1407;
      35917:data<=-16'd1086;
      35918:data<=-16'd229;
      35919:data<=16'd1248;
      35920:data<=16'd2531;
      35921:data<=16'd3021;
      35922:data<=16'd3222;
      35923:data<=16'd3278;
      35924:data<=16'd2786;
      35925:data<=16'd3130;
      35926:data<=16'd5156;
      35927:data<=16'd5888;
      35928:data<=16'd5272;
      35929:data<=16'd5692;
      35930:data<=16'd5153;
      35931:data<=16'd4643;
      35932:data<=16'd6849;
      35933:data<=16'd8170;
      35934:data<=16'd7896;
      35935:data<=16'd8228;
      35936:data<=16'd7821;
      35937:data<=16'd7652;
      35938:data<=16'd8657;
      35939:data<=16'd9263;
      35940:data<=16'd9632;
      35941:data<=16'd9118;
      35942:data<=16'd8150;
      35943:data<=16'd8698;
      35944:data<=16'd9555;
      35945:data<=16'd9903;
      35946:data<=16'd10129;
      35947:data<=16'd10245;
      35948:data<=16'd10408;
      35949:data<=16'd9529;
      35950:data<=16'd9239;
      35951:data<=16'd10784;
      35952:data<=16'd10677;
      35953:data<=16'd9937;
      35954:data<=16'd10373;
      35955:data<=16'd9746;
      35956:data<=16'd10107;
      35957:data<=16'd11538;
      35958:data<=16'd11042;
      35959:data<=16'd10329;
      35960:data<=16'd8492;
      35961:data<=16'd5385;
      35962:data<=16'd5797;
      35963:data<=16'd7858;
      35964:data<=16'd7918;
      35965:data<=16'd7674;
      35966:data<=16'd7526;
      35967:data<=16'd7006;
      35968:data<=16'd6692;
      35969:data<=16'd7225;
      35970:data<=16'd8384;
      35971:data<=16'd8507;
      35972:data<=16'd8279;
      35973:data<=16'd8291;
      35974:data<=16'd7450;
      35975:data<=16'd7928;
      35976:data<=16'd9615;
      35977:data<=16'd9424;
      35978:data<=16'd8713;
      35979:data<=16'd8469;
      35980:data<=16'd7944;
      35981:data<=16'd8627;
      35982:data<=16'd10182;
      35983:data<=16'd10625;
      35984:data<=16'd9826;
      35985:data<=16'd8746;
      35986:data<=16'd8357;
      35987:data<=16'd8751;
      35988:data<=16'd9392;
      35989:data<=16'd9671;
      35990:data<=16'd9647;
      35991:data<=16'd9561;
      35992:data<=16'd8520;
      35993:data<=16'd7952;
      35994:data<=16'd9553;
      35995:data<=16'd10320;
      35996:data<=16'd9509;
      35997:data<=16'd9347;
      35998:data<=16'd8536;
      35999:data<=16'd7421;
      36000:data<=16'd8614;
      36001:data<=16'd10258;
      36002:data<=16'd9811;
      36003:data<=16'd8877;
      36004:data<=16'd8816;
      36005:data<=16'd8355;
      36006:data<=16'd8282;
      36007:data<=16'd9814;
      36008:data<=16'd10298;
      36009:data<=16'd9846;
      36010:data<=16'd10998;
      36011:data<=16'd11850;
      36012:data<=16'd11468;
      36013:data<=16'd11212;
      36014:data<=16'd10845;
      36015:data<=16'd10569;
      36016:data<=16'd9985;
      36017:data<=16'd9445;
      36018:data<=16'd9876;
      36019:data<=16'd8812;
      36020:data<=16'd6625;
      36021:data<=16'd5912;
      36022:data<=16'd4949;
      36023:data<=16'd3794;
      36024:data<=16'd3892;
      36025:data<=16'd3354;
      36026:data<=16'd1757;
      36027:data<=16'd607;
      36028:data<=16'd356;
      36029:data<=16'd246;
      36030:data<=-16'd323;
      36031:data<=-16'd614;
      36032:data<=-16'd1128;
      36033:data<=-16'd2106;
      36034:data<=-16'd2290;
      36035:data<=-16'd2464;
      36036:data<=-16'd2563;
      36037:data<=-16'd2077;
      36038:data<=-16'd2928;
      36039:data<=-16'd4090;
      36040:data<=-16'd4176;
      36041:data<=-16'd5049;
      36042:data<=-16'd5805;
      36043:data<=-16'd5125;
      36044:data<=-16'd5377;
      36045:data<=-16'd6963;
      36046:data<=-16'd7373;
      36047:data<=-16'd6860;
      36048:data<=-16'd7054;
      36049:data<=-16'd6837;
      36050:data<=-16'd6865;
      36051:data<=-16'd8577;
      36052:data<=-16'd8997;
      36053:data<=-16'd8119;
      36054:data<=-16'd8185;
      36055:data<=-16'd7541;
      36056:data<=-16'd7617;
      36057:data<=-16'd9277;
      36058:data<=-16'd9141;
      36059:data<=-16'd9133;
      36060:data<=-16'd11194;
      36061:data<=-16'd12554;
      36062:data<=-16'd12938;
      36063:data<=-16'd13397;
      36064:data<=-16'd14038;
      36065:data<=-16'd14070;
      36066:data<=-16'd13239;
      36067:data<=-16'd12969;
      36068:data<=-16'd12519;
      36069:data<=-16'd12552;
      36070:data<=-16'd14149;
      36071:data<=-16'd13982;
      36072:data<=-16'd13365;
      36073:data<=-16'd13902;
      36074:data<=-16'd12445;
      36075:data<=-16'd12204;
      36076:data<=-16'd13808;
      36077:data<=-16'd12678;
      36078:data<=-16'd11872;
      36079:data<=-16'd12249;
      36080:data<=-16'd11320;
      36081:data<=-16'd11435;
      36082:data<=-16'd12011;
      36083:data<=-16'd11785;
      36084:data<=-16'd11665;
      36085:data<=-16'd10749;
      36086:data<=-16'd9970;
      36087:data<=-16'd10085;
      36088:data<=-16'd10658;
      36089:data<=-16'd11637;
      36090:data<=-16'd11433;
      36091:data<=-16'd10924;
      36092:data<=-16'd10422;
      36093:data<=-16'd8784;
      36094:data<=-16'd9553;
      36095:data<=-16'd11630;
      36096:data<=-16'd10748;
      36097:data<=-16'd9996;
      36098:data<=-16'd9856;
      36099:data<=-16'd8463;
      36100:data<=-16'd8689;
      36101:data<=-16'd9917;
      36102:data<=-16'd9837;
      36103:data<=-16'd9614;
      36104:data<=-16'd9292;
      36105:data<=-16'd8284;
      36106:data<=-16'd7524;
      36107:data<=-16'd8223;
      36108:data<=-16'd9532;
      36109:data<=-16'd8475;
      36110:data<=-16'd5168;
      36111:data<=-16'd2869;
      36112:data<=-16'd2270;
      36113:data<=-16'd1776;
      36114:data<=-16'd1360;
      36115:data<=-16'd1447;
      36116:data<=-16'd1152;
      36117:data<=-16'd873;
      36118:data<=-16'd717;
      36119:data<=16'd911;
      36120:data<=16'd2455;
      36121:data<=16'd2594;
      36122:data<=16'd3021;
      36123:data<=16'd2877;
      36124:data<=16'd2290;
      36125:data<=16'd3416;
      36126:data<=16'd4616;
      36127:data<=16'd4464;
      36128:data<=16'd4291;
      36129:data<=16'd4811;
      36130:data<=16'd5262;
      36131:data<=16'd5039;
      36132:data<=16'd5780;
      36133:data<=16'd7068;
      36134:data<=16'd6731;
      36135:data<=16'd6640;
      36136:data<=16'd7028;
      36137:data<=16'd6607;
      36138:data<=16'd7582;
      36139:data<=16'd8789;
      36140:data<=16'd8244;
      36141:data<=16'd8229;
      36142:data<=16'd8326;
      36143:data<=16'd7551;
      36144:data<=16'd8143;
      36145:data<=16'd9647;
      36146:data<=16'd9511;
      36147:data<=16'd8692;
      36148:data<=16'd9166;
      36149:data<=16'd9188;
      36150:data<=16'd8158;
      36151:data<=16'd8649;
      36152:data<=16'd9617;
      36153:data<=16'd9172;
      36154:data<=16'd8862;
      36155:data<=16'd9022;
      36156:data<=16'd8783;
      36157:data<=16'd8963;
      36158:data<=16'd10568;
      36159:data<=16'd10948;
      36160:data<=16'd7598;
      36161:data<=16'd4711;
      36162:data<=16'd4557;
      36163:data<=16'd5265;
      36164:data<=16'd7485;
      36165:data<=16'd8267;
      36166:data<=16'd6557;
      36167:data<=16'd6626;
      36168:data<=16'd6441;
      36169:data<=16'd6216;
      36170:data<=16'd8182;
      36171:data<=16'd7735;
      36172:data<=16'd6669;
      36173:data<=16'd7318;
      36174:data<=16'd6112;
      36175:data<=16'd6081;
      36176:data<=16'd7852;
      36177:data<=16'd8225;
      36178:data<=16'd8413;
      36179:data<=16'd7388;
      36180:data<=16'd6002;
      36181:data<=16'd6487;
      36182:data<=16'd7300;
      36183:data<=16'd8425;
      36184:data<=16'd8170;
      36185:data<=16'd6871;
      36186:data<=16'd7385;
      36187:data<=16'd6862;
      36188:data<=16'd6755;
      36189:data<=16'd8796;
      36190:data<=16'd8232;
      36191:data<=16'd7206;
      36192:data<=16'd7718;
      36193:data<=16'd7292;
      36194:data<=16'd7256;
      36195:data<=16'd7292;
      36196:data<=16'd7383;
      36197:data<=16'd7474;
      36198:data<=16'd5874;
      36199:data<=16'd5721;
      36200:data<=16'd6846;
      36201:data<=16'd7368;
      36202:data<=16'd8711;
      36203:data<=16'd7887;
      36204:data<=16'd6018;
      36205:data<=16'd6114;
      36206:data<=16'd5298;
      36207:data<=16'd5288;
      36208:data<=16'd6373;
      36209:data<=16'd6511;
      36210:data<=16'd8282;
      36211:data<=16'd9712;
      36212:data<=16'd9435;
      36213:data<=16'd8745;
      36214:data<=16'd6755;
      36215:data<=16'd6488;
      36216:data<=16'd6943;
      36217:data<=16'd5800;
      36218:data<=16'd6225;
      36219:data<=16'd4963;
      36220:data<=16'd1923;
      36221:data<=16'd2469;
      36222:data<=16'd2945;
      36223:data<=16'd1234;
      36224:data<=16'd341;
      36225:data<=16'd741;
      36226:data<=16'd573;
      36227:data<=-16'd2023;
      36228:data<=-16'd3187;
      36229:data<=-16'd2400;
      36230:data<=-16'd3203;
      36231:data<=-16'd2731;
      36232:data<=-16'd3134;
      36233:data<=-16'd5764;
      36234:data<=-16'd5479;
      36235:data<=-16'd5241;
      36236:data<=-16'd4896;
      36237:data<=-16'd3416;
      36238:data<=-16'd5959;
      36239:data<=-16'd7494;
      36240:data<=-16'd6431;
      36241:data<=-16'd7144;
      36242:data<=-16'd6413;
      36243:data<=-16'd6525;
      36244:data<=-16'd7877;
      36245:data<=-16'd7823;
      36246:data<=-16'd10110;
      36247:data<=-16'd10671;
      36248:data<=-16'd8987;
      36249:data<=-16'd9506;
      36250:data<=-16'd8348;
      36251:data<=-16'd9360;
      36252:data<=-16'd12425;
      36253:data<=-16'd8793;
      36254:data<=-16'd2065;
      36255:data<=16'd2663;
      36256:data<=-16'd252;
      36257:data<=-16'd9774;
      36258:data<=-16'd11342;
      36259:data<=-16'd8943;
      36260:data<=-16'd10707;
      36261:data<=-16'd10454;
      36262:data<=-16'd10204;
      36263:data<=-16'd9938;
      36264:data<=-16'd9280;
      36265:data<=-16'd10473;
      36266:data<=-16'd9130;
      36267:data<=-16'd14856;
      36268:data<=-16'd23340;
      36269:data<=-16'd16263;
      36270:data<=-16'd15659;
      36271:data<=-16'd29645;
      36272:data<=-16'd31216;
      36273:data<=-16'd26368;
      36274:data<=-16'd26491;
      36275:data<=-16'd24996;
      36276:data<=-16'd24714;
      36277:data<=-16'd23971;
      36278:data<=-16'd21946;
      36279:data<=-16'd22316;
      36280:data<=-16'd20971;
      36281:data<=-16'd20519;
      36282:data<=-16'd21961;
      36283:data<=-16'd20600;
      36284:data<=-16'd19381;
      36285:data<=-16'd18586;
      36286:data<=-16'd17917;
      36287:data<=-16'd18315;
      36288:data<=-16'd16666;
      36289:data<=-16'd15368;
      36290:data<=-16'd15600;
      36291:data<=-16'd14898;
      36292:data<=-16'd13999;
      36293:data<=-16'd12460;
      36294:data<=-16'd12975;
      36295:data<=-16'd14753;
      36296:data<=-16'd12546;
      36297:data<=-16'd11324;
      36298:data<=-16'd11975;
      36299:data<=-16'd10066;
      36300:data<=-16'd9450;
      36301:data<=-16'd9398;
      36302:data<=-16'd7858;
      36303:data<=-16'd7295;
      36304:data<=-16'd6473;
      36305:data<=-16'd6428;
      36306:data<=-16'd7442;
      36307:data<=-16'd7286;
      36308:data<=-16'd7212;
      36309:data<=-16'd6473;
      36310:data<=-16'd6119;
      36311:data<=-16'd6642;
      36312:data<=-16'd4760;
      36313:data<=-16'd4158;
      36314:data<=-16'd4875;
      36315:data<=-16'd3501;
      36316:data<=-16'd3659;
      36317:data<=-16'd2235;
      36318:data<=-16'd829;
      36319:data<=-16'd5383;
      36320:data<=-16'd1383;
      36321:data<=16'd12571;
      36322:data<=16'd16184;
      36323:data<=16'd13159;
      36324:data<=16'd13882;
      36325:data<=16'd12872;
      36326:data<=16'd12061;
      36327:data<=16'd13773;
      36328:data<=16'd12599;
      36329:data<=16'd11103;
      36330:data<=16'd12311;
      36331:data<=16'd12085;
      36332:data<=16'd10207;
      36333:data<=16'd9864;
      36334:data<=16'd10392;
      36335:data<=16'd9887;
      36336:data<=16'd8827;
      36337:data<=16'd8445;
      36338:data<=16'd8646;
      36339:data<=16'd8202;
      36340:data<=16'd7412;
      36341:data<=16'd8003;
      36342:data<=16'd8939;
      36343:data<=16'd8358;
      36344:data<=16'd7172;
      36345:data<=16'd6055;
      36346:data<=16'd5441;
      36347:data<=16'd5817;
      36348:data<=16'd5758;
      36349:data<=16'd5388;
      36350:data<=16'd5600;
      36351:data<=16'd5356;
      36352:data<=16'd4990;
      36353:data<=16'd4813;
      36354:data<=16'd4760;
      36355:data<=16'd5429;
      36356:data<=16'd4481;
      36357:data<=16'd2362;
      36358:data<=16'd2252;
      36359:data<=16'd1803;
      36360:data<=16'd1245;
      36361:data<=16'd2469;
      36362:data<=16'd1783;
      36363:data<=16'd702;
      36364:data<=16'd1563;
      36365:data<=16'd1950;
      36366:data<=16'd3253;
      36367:data<=16'd2930;
      36368:data<=16'd789;
      36369:data<=16'd2532;
      36370:data<=-16'd1985;
      36371:data<=-16'd15073;
      36372:data<=-16'd18295;
      36373:data<=-16'd14665;
      36374:data<=-16'd15429;
      36375:data<=-16'd14515;
      36376:data<=-16'd12951;
      36377:data<=-16'd13438;
      36378:data<=-16'd12007;
      36379:data<=-16'd11543;
      36380:data<=-16'd11835;
      36381:data<=-16'd10830;
      36382:data<=-16'd11294;
      36383:data<=-16'd11503;
      36384:data<=-16'd10813;
      36385:data<=-16'd10434;
      36386:data<=-16'd9229;
      36387:data<=-16'd8957;
      36388:data<=-16'd8774;
      36389:data<=-16'd6790;
      36390:data<=-16'd5764;
      36391:data<=-16'd6021;
      36392:data<=-16'd6159;
      36393:data<=-16'd5695;
      36394:data<=-16'd5206;
      36395:data<=-16'd6044;
      36396:data<=-16'd5985;
      36397:data<=-16'd5236;
      36398:data<=-16'd5786;
      36399:data<=-16'd4566;
      36400:data<=-16'd2801;
      36401:data<=-16'd3230;
      36402:data<=-16'd3263;
      36403:data<=-16'd2957;
      36404:data<=-16'd2590;
      36405:data<=-16'd1964;
      36406:data<=-16'd3010;
      36407:data<=-16'd4027;
      36408:data<=-16'd3692;
      36409:data<=-16'd3048;
      36410:data<=-16'd2237;
      36411:data<=-16'd1888;
      36412:data<=-16'd1445;
      36413:data<=-16'd1130;
      36414:data<=-16'd688;
      36415:data<=16'd447;
      36416:data<=-16'd694;
      36417:data<=-16'd252;
      36418:data<=16'd2478;
      36419:data<=-16'd657;
      36420:data<=16'd1492;
      36421:data<=16'd15092;
      36422:data<=16'd19688;
      36423:data<=16'd15791;
      36424:data<=16'd16995;
      36425:data<=16'd17191;
      36426:data<=16'd15744;
      36427:data<=16'd16433;
      36428:data<=16'd15500;
      36429:data<=16'd15249;
      36430:data<=16'd16049;
      36431:data<=16'd14709;
      36432:data<=16'd13362;
      36433:data<=16'd12775;
      36434:data<=16'd12478;
      36435:data<=16'd12134;
      36436:data<=16'd11482;
      36437:data<=16'd11734;
      36438:data<=16'd11079;
      36439:data<=16'd9943;
      36440:data<=16'd11039;
      36441:data<=16'd11236;
      36442:data<=16'd9994;
      36443:data<=16'd10067;
      36444:data<=16'd9276;
      36445:data<=16'd7069;
      36446:data<=16'd6492;
      36447:data<=16'd7514;
      36448:data<=16'd7439;
      36449:data<=16'd6294;
      36450:data<=16'd6514;
      36451:data<=16'd7133;
      36452:data<=16'd6865;
      36453:data<=16'd6987;
      36454:data<=16'd6989;
      36455:data<=16'd6672;
      36456:data<=16'd6422;
      36457:data<=16'd6041;
      36458:data<=16'd6478;
      36459:data<=16'd6470;
      36460:data<=16'd5882;
      36461:data<=16'd6443;
      36462:data<=16'd6206;
      36463:data<=16'd5592;
      36464:data<=16'd5483;
      36465:data<=16'd4915;
      36466:data<=16'd6476;
      36467:data<=16'd6711;
      36468:data<=16'd4150;
      36469:data<=16'd6305;
      36470:data<=16'd5259;
      36471:data<=-16'd5624;
      36472:data<=-16'd11291;
      36473:data<=-16'd9436;
      36474:data<=-16'd9518;
      36475:data<=-16'd9153;
      36476:data<=-16'd8034;
      36477:data<=-16'd8140;
      36478:data<=-16'd7344;
      36479:data<=-16'd7210;
      36480:data<=-16'd7617;
      36481:data<=-16'd6432;
      36482:data<=-16'd4831;
      36483:data<=-16'd3588;
      36484:data<=-16'd2998;
      36485:data<=-16'd2689;
      36486:data<=-16'd2507;
      36487:data<=-16'd2849;
      36488:data<=-16'd1603;
      36489:data<=-16'd14;
      36490:data<=-16'd685;
      36491:data<=-16'd696;
      36492:data<=-16'd21;
      36493:data<=-16'd375;
      36494:data<=16'd1034;
      36495:data<=16'd3582;
      36496:data<=16'd3996;
      36497:data<=16'd3193;
      36498:data<=16'd3362;
      36499:data<=16'd3971;
      36500:data<=16'd3533;
      36501:data<=16'd3433;
      36502:data<=16'd4077;
      36503:data<=16'd3497;
      36504:data<=16'd3177;
      36505:data<=16'd3586;
      36506:data<=16'd3566;
      36507:data<=16'd4928;
      36508:data<=16'd6003;
      36509:data<=16'd5369;
      36510:data<=16'd5932;
      36511:data<=16'd6279;
      36512:data<=16'd5457;
      36513:data<=16'd5752;
      36514:data<=16'd6146;
      36515:data<=16'd5764;
      36516:data<=16'd5109;
      36517:data<=16'd5491;
      36518:data<=16'd6375;
      36519:data<=16'd4972;
      36520:data<=16'd8536;
      36521:data<=16'd20381;
      36522:data<=16'd25857;
      36523:data<=16'd23052;
      36524:data<=16'd22838;
      36525:data<=16'd23008;
      36526:data<=16'd21789;
      36527:data<=16'd21547;
      36528:data<=16'd19943;
      36529:data<=16'd18782;
      36530:data<=16'd18956;
      36531:data<=16'd18574;
      36532:data<=16'd19382;
      36533:data<=16'd19590;
      36534:data<=16'd18158;
      36535:data<=16'd17678;
      36536:data<=16'd16283;
      36537:data<=16'd14465;
      36538:data<=16'd14842;
      36539:data<=16'd14842;
      36540:data<=16'd13718;
      36541:data<=16'd13065;
      36542:data<=16'd12501;
      36543:data<=16'd12151;
      36544:data<=16'd12408;
      36545:data<=16'd13018;
      36546:data<=16'd12862;
      36547:data<=16'd11621;
      36548:data<=16'd11242;
      36549:data<=16'd11527;
      36550:data<=16'd10804;
      36551:data<=16'd9859;
      36552:data<=16'd9570;
      36553:data<=16'd9541;
      36554:data<=16'd8819;
      36555:data<=16'd7485;
      36556:data<=16'd7250;
      36557:data<=16'd8217;
      36558:data<=16'd9362;
      36559:data<=16'd9828;
      36560:data<=16'd8831;
      36561:data<=16'd7782;
      36562:data<=16'd7524;
      36563:data<=16'd7118;
      36564:data<=16'd6540;
      36565:data<=16'd5715;
      36566:data<=16'd5900;
      36567:data<=16'd6605;
      36568:data<=16'd4772;
      36569:data<=16'd4071;
      36570:data<=16'd4364;
      36571:data<=-16'd3019;
      36572:data<=-16'd12029;
      36573:data<=-16'd12546;
      36574:data<=-16'd11594;
      36575:data<=-16'd12804;
      36576:data<=-16'd11855;
      36577:data<=-16'd11088;
      36578:data<=-16'd11304;
      36579:data<=-16'd10739;
      36580:data<=-16'd11148;
      36581:data<=-16'd11679;
      36582:data<=-16'd10416;
      36583:data<=-16'd8701;
      36584:data<=-16'd7797;
      36585:data<=-16'd7439;
      36586:data<=-16'd6969;
      36587:data<=-16'd6798;
      36588:data<=-16'd7094;
      36589:data<=-16'd7107;
      36590:data<=-16'd7145;
      36591:data<=-16'd7000;
      36592:data<=-16'd6622;
      36593:data<=-16'd6771;
      36594:data<=-16'd6020;
      36595:data<=-16'd4141;
      36596:data<=-16'd3156;
      36597:data<=-16'd3283;
      36598:data<=-16'd3891;
      36599:data<=-16'd4012;
      36600:data<=-16'd3621;
      36601:data<=-16'd3668;
      36602:data<=-16'd3339;
      36603:data<=-16'd3216;
      36604:data<=-16'd3724;
      36605:data<=-16'd3415;
      36606:data<=-16'd3682;
      36607:data<=-16'd3756;
      36608:data<=-16'd2182;
      36609:data<=-16'd2302;
      36610:data<=-16'd3159;
      36611:data<=-16'd2608;
      36612:data<=-16'd2428;
      36613:data<=-16'd1665;
      36614:data<=-16'd1196;
      36615:data<=-16'd2044;
      36616:data<=-16'd2246;
      36617:data<=-16'd2887;
      36618:data<=-16'd2223;
      36619:data<=-16'd746;
      36620:data<=-16'd1409;
      36621:data<=16'd4951;
      36622:data<=16'd16613;
      36623:data<=16'd17970;
      36624:data<=16'd14559;
      36625:data<=16'd15288;
      36626:data<=16'd14458;
      36627:data<=16'd13047;
      36628:data<=16'd13142;
      36629:data<=16'd12098;
      36630:data<=16'd11350;
      36631:data<=16'd11312;
      36632:data<=16'd11823;
      36633:data<=16'd12637;
      36634:data<=16'd12069;
      36635:data<=16'd11288;
      36636:data<=16'd10064;
      36637:data<=16'd8627;
      36638:data<=16'd9342;
      36639:data<=16'd9386;
      36640:data<=16'd7802;
      36641:data<=16'd7514;
      36642:data<=16'd7309;
      36643:data<=16'd6549;
      36644:data<=16'd6551;
      36645:data<=16'd7110;
      36646:data<=16'd7248;
      36647:data<=16'd6184;
      36648:data<=16'd5627;
      36649:data<=16'd5929;
      36650:data<=16'd5225;
      36651:data<=16'd4625;
      36652:data<=16'd4355;
      36653:data<=16'd3662;
      36654:data<=16'd3166;
      36655:data<=16'd2115;
      36656:data<=16'd1444;
      36657:data<=16'd1988;
      36658:data<=16'd2281;
      36659:data<=16'd2138;
      36660:data<=16'd813;
      36661:data<=-16'd419;
      36662:data<=-16'd203;
      36663:data<=-16'd1174;
      36664:data<=-16'd1550;
      36665:data<=-16'd883;
      36666:data<=-16'd1791;
      36667:data<=-16'd1098;
      36668:data<=-16'd1683;
      36669:data<=-16'd4388;
      36670:data<=-16'd2500;
      36671:data<=-16'd6690;
      36672:data<=-16'd20269;
      36673:data<=-16'd24090;
      36674:data<=-16'd20397;
      36675:data<=-16'd21120;
      36676:data<=-16'd21126;
      36677:data<=-16'd20196;
      36678:data<=-16'd20359;
      36679:data<=-16'd19155;
      36680:data<=-16'd18794;
      36681:data<=-16'd18462;
      36682:data<=-16'd17885;
      36683:data<=-16'd19293;
      36684:data<=-16'd19400;
      36685:data<=-16'd18299;
      36686:data<=-16'd17937;
      36687:data<=-16'd16753;
      36688:data<=-16'd16298;
      36689:data<=-16'd16454;
      36690:data<=-16'd15697;
      36691:data<=-16'd15913;
      36692:data<=-16'd16057;
      36693:data<=-16'd14863;
      36694:data<=-16'd14468;
      36695:data<=-16'd15136;
      36696:data<=-16'd15377;
      36697:data<=-16'd14894;
      36698:data<=-16'd14795;
      36699:data<=-16'd14833;
      36700:data<=-16'd14128;
      36701:data<=-16'd13787;
      36702:data<=-16'd13386;
      36703:data<=-16'd12693;
      36704:data<=-16'd12853;
      36705:data<=-16'd12173;
      36706:data<=-16'd11160;
      36707:data<=-16'd11670;
      36708:data<=-16'd12019;
      36709:data<=-16'd12003;
      36710:data<=-16'd11770;
      36711:data<=-16'd11232;
      36712:data<=-16'd11265;
      36713:data<=-16'd10592;
      36714:data<=-16'd10191;
      36715:data<=-16'd10267;
      36716:data<=-16'd9192;
      36717:data<=-16'd9840;
      36718:data<=-16'd9502;
      36719:data<=-16'd7482;
      36720:data<=-16'd10187;
      36721:data<=-16'd7042;
      36722:data<=16'd6158;
      36723:data<=16'd10196;
      36724:data<=16'd6452;
      36725:data<=16'd7645;
      36726:data<=16'd8217;
      36727:data<=16'd7063;
      36728:data<=16'd7286;
      36729:data<=16'd6560;
      36730:data<=16'd6789;
      36731:data<=16'd7247;
      36732:data<=16'd5965;
      36733:data<=16'd4960;
      36734:data<=16'd3858;
      36735:data<=16'd3529;
      36736:data<=16'd4053;
      36737:data<=16'd3318;
      36738:data<=16'd3118;
      36739:data<=16'd3200;
      36740:data<=16'd2719;
      36741:data<=16'd3460;
      36742:data<=16'd3466;
      36743:data<=16'd2660;
      36744:data<=16'd3066;
      36745:data<=16'd2337;
      36746:data<=16'd516;
      36747:data<=16'd24;
      36748:data<=16'd112;
      36749:data<=16'd36;
      36750:data<=16'd317;
      36751:data<=16'd560;
      36752:data<=16'd50;
      36753:data<=16'd17;
      36754:data<=16'd858;
      36755:data<=16'd743;
      36756:data<=16'd450;
      36757:data<=16'd89;
      36758:data<=-16'd1732;
      36759:data<=-16'd2660;
      36760:data<=-16'd2526;
      36761:data<=-16'd2845;
      36762:data<=-16'd2657;
      36763:data<=-16'd2972;
      36764:data<=-16'd3119;
      36765:data<=-16'd2620;
      36766:data<=-16'd3259;
      36767:data<=-16'd2610;
      36768:data<=-16'd2366;
      36769:data<=-16'd3739;
      36770:data<=-16'd2544;
      36771:data<=-16'd7621;
      36772:data<=-16'd20604;
      36773:data<=-16'd24146;
      36774:data<=-16'd20654;
      36775:data<=-16'd21199;
      36776:data<=-16'd20782;
      36777:data<=-16'd19544;
      36778:data<=-16'd19420;
      36779:data<=-16'd17538;
      36780:data<=-16'd17014;
      36781:data<=-16'd16953;
      36782:data<=-16'd15541;
      36783:data<=-16'd16422;
      36784:data<=-16'd17206;
      36785:data<=-16'd15887;
      36786:data<=-16'd14962;
      36787:data<=-16'd14166;
      36788:data<=-16'd13693;
      36789:data<=-16'd13435;
      36790:data<=-16'd12763;
      36791:data<=-16'd12483;
      36792:data<=-16'd11693;
      36793:data<=-16'd10530;
      36794:data<=-16'd9899;
      36795:data<=-16'd9720;
      36796:data<=-16'd10496;
      36797:data<=-16'd10366;
      36798:data<=-16'd9235;
      36799:data<=-16'd9377;
      36800:data<=-16'd8984;
      36801:data<=-16'd7912;
      36802:data<=-16'd7518;
      36803:data<=-16'd6795;
      36804:data<=-16'd6664;
      36805:data<=-16'd6361;
      36806:data<=-16'd5204;
      36807:data<=-16'd5758;
      36808:data<=-16'd6701;
      36809:data<=-16'd6658;
      36810:data<=-16'd6423;
      36811:data<=-16'd5442;
      36812:data<=-16'd4899;
      36813:data<=-16'd4570;
      36814:data<=-16'd3750;
      36815:data<=-16'd3410;
      36816:data<=-16'd2658;
      36817:data<=-16'd2781;
      36818:data<=-16'd2329;
      36819:data<=16'd64;
      36820:data<=-16'd1762;
      36821:data<=-16'd308;
      36822:data<=16'd11734;
      36823:data<=16'd17468;
      36824:data<=16'd14389;
      36825:data<=16'd15245;
      36826:data<=16'd15662;
      36827:data<=16'd14401;
      36828:data<=16'd14941;
      36829:data<=16'd13068;
      36830:data<=16'd12187;
      36831:data<=16'd13970;
      36832:data<=16'd12957;
      36833:data<=16'd10839;
      36834:data<=16'd10120;
      36835:data<=16'd10125;
      36836:data<=16'd9809;
      36837:data<=16'd8721;
      36838:data<=16'd9122;
      36839:data<=16'd9621;
      36840:data<=16'd8802;
      36841:data<=16'd8989;
      36842:data<=16'd8578;
      36843:data<=16'd7874;
      36844:data<=16'd8651;
      36845:data<=16'd8120;
      36846:data<=16'd7004;
      36847:data<=16'd6849;
      36848:data<=16'd6505;
      36849:data<=16'd6549;
      36850:data<=16'd6445;
      36851:data<=16'd6379;
      36852:data<=16'd6890;
      36853:data<=16'd6487;
      36854:data<=16'd6326;
      36855:data<=16'd6607;
      36856:data<=16'd6144;
      36857:data<=16'd6264;
      36858:data<=16'd6634;
      36859:data<=16'd6614;
      36860:data<=16'd6297;
      36861:data<=16'd5985;
      36862:data<=16'd7175;
      36863:data<=16'd7962;
      36864:data<=16'd7526;
      36865:data<=16'd7627;
      36866:data<=16'd6763;
      36867:data<=16'd6122;
      36868:data<=16'd6041;
      36869:data<=16'd5081;
      36870:data<=16'd7007;
      36871:data<=16'd6078;
      36872:data<=-16'd3977;
      36873:data<=-16'd10431;
      36874:data<=-16'd8674;
      36875:data<=-16'd8153;
      36876:data<=-16'd8254;
      36877:data<=-16'd6818;
      36878:data<=-16'd6617;
      36879:data<=-16'd6569;
      36880:data<=-16'd5990;
      36881:data<=-16'd6103;
      36882:data<=-16'd5940;
      36883:data<=-16'd4244;
      36884:data<=-16'd2543;
      36885:data<=-16'd2278;
      36886:data<=-16'd1600;
      36887:data<=-16'd466;
      36888:data<=-16'd625;
      36889:data<=-16'd775;
      36890:data<=-16'd349;
      36891:data<=-16'd165;
      36892:data<=16'd209;
      36893:data<=16'd456;
      36894:data<=16'd143;
      36895:data<=16'd255;
      36896:data<=16'd1583;
      36897:data<=16'd2526;
      36898:data<=16'd2064;
      36899:data<=16'd2590;
      36900:data<=16'd3501;
      36901:data<=16'd2961;
      36902:data<=16'd3165;
      36903:data<=16'd3215;
      36904:data<=16'd2164;
      36905:data<=16'd2641;
      36906:data<=16'd2826;
      36907:data<=16'd2100;
      36908:data<=16'd3230;
      36909:data<=16'd4319;
      36910:data<=16'd4464;
      36911:data<=16'd5027;
      36912:data<=16'd4992;
      36913:data<=16'd4479;
      36914:data<=16'd4049;
      36915:data<=16'd3918;
      36916:data<=16'd4490;
      36917:data<=16'd4510;
      36918:data<=16'd4666;
      36919:data<=16'd5371;
      36920:data<=16'd4404;
      36921:data<=16'd6466;
      36922:data<=16'd16319;
      36923:data<=16'd24567;
      36924:data<=16'd24110;
      36925:data<=16'd22294;
      36926:data<=16'd22359;
      36927:data<=16'd20830;
      36928:data<=16'd19488;
      36929:data<=16'd19052;
      36930:data<=16'd18063;
      36931:data<=16'd17781;
      36932:data<=16'd17196;
      36933:data<=16'd16481;
      36934:data<=16'd17302;
      36935:data<=16'd17173;
      36936:data<=16'd16172;
      36937:data<=16'd15679;
      36938:data<=16'd14457;
      36939:data<=16'd13849;
      36940:data<=16'd13611;
      36941:data<=16'd12449;
      36942:data<=16'd12038;
      36943:data<=16'd11524;
      36944:data<=16'd10662;
      36945:data<=16'd10937;
      36946:data<=16'd11420;
      36947:data<=16'd12005;
      36948:data<=16'd11755;
      36949:data<=16'd10378;
      36950:data<=16'd10238;
      36951:data<=16'd10120;
      36952:data<=16'd9368;
      36953:data<=16'd9138;
      36954:data<=16'd8381;
      36955:data<=16'd8457;
      36956:data<=16'd8849;
      36957:data<=16'd7407;
      36958:data<=16'd7460;
      36959:data<=16'd9218;
      36960:data<=16'd9427;
      36961:data<=16'd8787;
      36962:data<=16'd8044;
      36963:data<=16'd7548;
      36964:data<=16'd7515;
      36965:data<=16'd6939;
      36966:data<=16'd6108;
      36967:data<=16'd5785;
      36968:data<=16'd5620;
      36969:data<=16'd4296;
      36970:data<=16'd3961;
      36971:data<=16'd5389;
      36972:data<=-16'd509;
      36973:data<=-16'd11586;
      36974:data<=-16'd13323;
      36975:data<=-16'd10563;
      36976:data<=-16'd12073;
      36977:data<=-16'd12002;
      36978:data<=-16'd10743;
      36979:data<=-16'd10748;
      36980:data<=-16'd9764;
      36981:data<=-16'd10122;
      36982:data<=-16'd10784;
      36983:data<=-16'd9207;
      36984:data<=-16'd7602;
      36985:data<=-16'd6388;
      36986:data<=-16'd6009;
      36987:data<=-16'd6332;
      36988:data<=-16'd5796;
      36989:data<=-16'd5680;
      36990:data<=-16'd5956;
      36991:data<=-16'd5912;
      36992:data<=-16'd6178;
      36993:data<=-16'd5984;
      36994:data<=-16'd5524;
      36995:data<=-16'd4958;
      36996:data<=-16'd4184;
      36997:data<=-16'd4067;
      36998:data<=-16'd3654;
      36999:data<=-16'd3265;
      37000:data<=-16'd3648;
      37001:data<=-16'd3298;
      37002:data<=-16'd2795;
      37003:data<=-16'd2889;
      37004:data<=-16'd3385;
      37005:data<=-16'd3970;
      37006:data<=-16'd3595;
      37007:data<=-16'd3821;
      37008:data<=-16'd3773;
      37009:data<=-16'd1566;
      37010:data<=-16'd1130;
      37011:data<=-16'd1812;
      37012:data<=-16'd1315;
      37013:data<=-16'd2074;
      37014:data<=-16'd2033;
      37015:data<=-16'd1336;
      37016:data<=-16'd1945;
      37017:data<=-16'd1383;
      37018:data<=-16'd1691;
      37019:data<=-16'd1794;
      37020:data<=-16'd335;
      37021:data<=-16'd1556;
      37022:data<=16'd3559;
      37023:data<=16'd16155;
      37024:data<=16'd18891;
      37025:data<=16'd15485;
      37026:data<=16'd16264;
      37027:data<=16'd15385;
      37028:data<=16'd13493;
      37029:data<=16'd12992;
      37030:data<=16'd12166;
      37031:data<=16'd12601;
      37032:data<=16'd11969;
      37033:data<=16'd11044;
      37034:data<=16'd12270;
      37035:data<=16'd11402;
      37036:data<=16'd9852;
      37037:data<=16'd9887;
      37038:data<=16'd8960;
      37039:data<=16'd8642;
      37040:data<=16'd8341;
      37041:data<=16'd6749;
      37042:data<=16'd6470;
      37043:data<=16'd6308;
      37044:data<=16'd5415;
      37045:data<=16'd5500;
      37046:data<=16'd6291;
      37047:data<=16'd7327;
      37048:data<=16'd7119;
      37049:data<=16'd5544;
      37050:data<=16'd4939;
      37051:data<=16'd4969;
      37052:data<=16'd4199;
      37053:data<=16'd2742;
      37054:data<=16'd2453;
      37055:data<=16'd3755;
      37056:data<=16'd3676;
      37057:data<=16'd2784;
      37058:data<=16'd2666;
      37059:data<=16'd1791;
      37060:data<=16'd1257;
      37061:data<=16'd1339;
      37062:data<=16'd1011;
      37063:data<=16'd858;
      37064:data<=-16'd223;
      37065:data<=-16'd792;
      37066:data<=-16'd522;
      37067:data<=-16'd1662;
      37068:data<=-16'd1230;
      37069:data<=-16'd1213;
      37070:data<=-16'd2989;
      37071:data<=-16'd1556;
      37072:data<=-16'd6526;
      37073:data<=-16'd19957;
      37074:data<=-16'd23519;
      37075:data<=-16'd19975;
      37076:data<=-16'd20700;
      37077:data<=-16'd20172;
      37078:data<=-16'd18826;
      37079:data<=-16'd19132;
      37080:data<=-16'd18124;
      37081:data<=-16'd18052;
      37082:data<=-16'd18117;
      37083:data<=-16'd17365;
      37084:data<=-16'd18221;
      37085:data<=-16'd17978;
      37086:data<=-16'd16691;
      37087:data<=-16'd16651;
      37088:data<=-16'd16175;
      37089:data<=-16'd15637;
      37090:data<=-16'd15317;
      37091:data<=-16'd14486;
      37092:data<=-16'd13866;
      37093:data<=-16'd13308;
      37094:data<=-16'd13038;
      37095:data<=-16'd12801;
      37096:data<=-16'd13303;
      37097:data<=-16'd15438;
      37098:data<=-16'd15361;
      37099:data<=-16'd13327;
      37100:data<=-16'd13338;
      37101:data<=-16'd13456;
      37102:data<=-16'd12713;
      37103:data<=-16'd11935;
      37104:data<=-16'd10939;
      37105:data<=-16'd11301;
      37106:data<=-16'd11327;
      37107:data<=-16'd10248;
      37108:data<=-16'd10939;
      37109:data<=-16'd11831;
      37110:data<=-16'd11570;
      37111:data<=-16'd11283;
      37112:data<=-16'd11006;
      37113:data<=-16'd10874;
      37114:data<=-16'd10038;
      37115:data<=-16'd9600;
      37116:data<=-16'd9699;
      37117:data<=-16'd8516;
      37118:data<=-16'd8848;
      37119:data<=-16'd8213;
      37120:data<=-16'd5862;
      37121:data<=-16'd8984;
      37122:data<=-16'd6796;
      37123:data<=16'd6537;
      37124:data<=16'd11282;
      37125:data<=16'd7756;
      37126:data<=16'd8484;
      37127:data<=16'd7993;
      37128:data<=16'd6849;
      37129:data<=16'd7958;
      37130:data<=16'd6843;
      37131:data<=16'd6470;
      37132:data<=16'd7319;
      37133:data<=16'd6006;
      37134:data<=16'd4123;
      37135:data<=16'd2716;
      37136:data<=16'd2990;
      37137:data<=16'd3544;
      37138:data<=16'd2466;
      37139:data<=16'd2487;
      37140:data<=16'd2406;
      37141:data<=16'd1762;
      37142:data<=16'd2497;
      37143:data<=16'd1867;
      37144:data<=16'd1309;
      37145:data<=16'd2202;
      37146:data<=16'd1306;
      37147:data<=16'd581;
      37148:data<=16'd684;
      37149:data<=16'd143;
      37150:data<=16'd344;
      37151:data<=16'd235;
      37152:data<=16'd18;
      37153:data<=16'd140;
      37154:data<=-16'd585;
      37155:data<=-16'd318;
      37156:data<=-16'd5;
      37157:data<=-16'd544;
      37158:data<=-16'd378;
      37159:data<=-16'd1547;
      37160:data<=-16'd2761;
      37161:data<=-16'd2291;
      37162:data<=-16'd2508;
      37163:data<=-16'd2244;
      37164:data<=-16'd1689;
      37165:data<=-16'd1932;
      37166:data<=-16'd1835;
      37167:data<=-16'd2373;
      37168:data<=-16'd2291;
      37169:data<=-16'd2211;
      37170:data<=-16'd2626;
      37171:data<=-16'd711;
      37172:data<=-16'd5483;
      37173:data<=-16'd18443;
      37174:data<=-16'd22973;
      37175:data<=-16'd20139;
      37176:data<=-16'd19626;
      37177:data<=-16'd18719;
      37178:data<=-16'd17895;
      37179:data<=-16'd17602;
      37180:data<=-16'd16293;
      37181:data<=-16'd16057;
      37182:data<=-16'd15670;
      37183:data<=-16'd15258;
      37184:data<=-16'd15368;
      37185:data<=-16'd14381;
      37186:data<=-16'd14143;
      37187:data<=-16'd13499;
      37188:data<=-16'd11970;
      37189:data<=-16'd12351;
      37190:data<=-16'd11961;
      37191:data<=-16'd10530;
      37192:data<=-16'd9946;
      37193:data<=-16'd9050;
      37194:data<=-16'd8754;
      37195:data<=-16'd8093;
      37196:data<=-16'd7899;
      37197:data<=-16'd10281;
      37198:data<=-16'd10643;
      37199:data<=-16'd9241;
      37200:data<=-16'd8818;
      37201:data<=-16'd7456;
      37202:data<=-16'd7147;
      37203:data<=-16'd7119;
      37204:data<=-16'd5586;
      37205:data<=-16'd5796;
      37206:data<=-16'd5946;
      37207:data<=-16'd5148;
      37208:data<=-16'd5510;
      37209:data<=-16'd5900;
      37210:data<=-16'd7015;
      37211:data<=-16'd7013;
      37212:data<=-16'd5157;
      37213:data<=-16'd5244;
      37214:data<=-16'd4852;
      37215:data<=-16'd3630;
      37216:data<=-16'd3571;
      37217:data<=-16'd2475;
      37218:data<=-16'd2858;
      37219:data<=-16'd2889;
      37220:data<=-16'd717;
      37221:data<=-16'd3193;
      37222:data<=-16'd2259;
      37223:data<=16'd9148;
      37224:data<=16'd16037;
      37225:data<=16'd14442;
      37226:data<=16'd13476;
      37227:data<=16'd13540;
      37228:data<=16'd13496;
      37229:data<=16'd13288;
      37230:data<=16'd12569;
      37231:data<=16'd12219;
      37232:data<=16'd11913;
      37233:data<=16'd11549;
      37234:data<=16'd10151;
      37235:data<=16'd8379;
      37236:data<=16'd8724;
      37237:data<=16'd8819;
      37238:data<=16'd7973;
      37239:data<=16'd8428;
      37240:data<=16'd8355;
      37241:data<=16'd7574;
      37242:data<=16'd7370;
      37243:data<=16'd6905;
      37244:data<=16'd6743;
      37245:data<=16'd6943;
      37246:data<=16'd6540;
      37247:data<=16'd5404;
      37248:data<=16'd4734;
      37249:data<=16'd5815;
      37250:data<=16'd5887;
      37251:data<=16'd4384;
      37252:data<=16'd4854;
      37253:data<=16'd5459;
      37254:data<=16'd4730;
      37255:data<=16'd4948;
      37256:data<=16'd5221;
      37257:data<=16'd5335;
      37258:data<=16'd5368;
      37259:data<=16'd4537;
      37260:data<=16'd4990;
      37261:data<=16'd5867;
      37262:data<=16'd5197;
      37263:data<=16'd4866;
      37264:data<=16'd4786;
      37265:data<=16'd4654;
      37266:data<=16'd4781;
      37267:data<=16'd4469;
      37268:data<=16'd5122;
      37269:data<=16'd4927;
      37270:data<=16'd3165;
      37271:data<=16'd5010;
      37272:data<=16'd5103;
      37273:data<=-16'd3883;
      37274:data<=-16'd11728;
      37275:data<=-16'd11330;
      37276:data<=-16'd9659;
      37277:data<=-16'd9547;
      37278:data<=-16'd9051;
      37279:data<=-16'd8302;
      37280:data<=-16'd7442;
      37281:data<=-16'd7118;
      37282:data<=-16'd7333;
      37283:data<=-16'd6713;
      37284:data<=-16'd5422;
      37285:data<=-16'd4270;
      37286:data<=-16'd3369;
      37287:data<=-16'd2887;
      37288:data<=-16'd2654;
      37289:data<=-16'd2403;
      37290:data<=-16'd2141;
      37291:data<=-16'd1710;
      37292:data<=-16'd1148;
      37293:data<=-16'd810;
      37294:data<=-16'd751;
      37295:data<=-16'd522;
      37296:data<=16'd311;
      37297:data<=16'd1392;
      37298:data<=16'd1785;
      37299:data<=16'd1647;
      37300:data<=16'd2064;
      37301:data<=16'd2645;
      37302:data<=16'd2564;
      37303:data<=16'd2573;
      37304:data<=16'd2869;
      37305:data<=16'd2878;
      37306:data<=16'd2811;
      37307:data<=16'd2453;
      37308:data<=16'd2285;
      37309:data<=16'd3551;
      37310:data<=16'd4837;
      37311:data<=16'd4792;
      37312:data<=16'd4607;
      37313:data<=16'd4592;
      37314:data<=16'd4720;
      37315:data<=16'd5213;
      37316:data<=16'd5122;
      37317:data<=16'd4745;
      37318:data<=16'd4598;
      37319:data<=16'd4595;
      37320:data<=16'd5471;
      37321:data<=16'd5165;
      37322:data<=16'd5177;
      37323:data<=16'd13291;
      37324:data<=16'd23958;
      37325:data<=16'd24959;
      37326:data<=16'd21992;
      37327:data<=16'd22315;
      37328:data<=16'd21699;
      37329:data<=16'd20377;
      37330:data<=16'd20007;
      37331:data<=16'd18816;
      37332:data<=16'd18073;
      37333:data<=16'd17573;
      37334:data<=16'd17174;
      37335:data<=16'd18325;
      37336:data<=16'd18181;
      37337:data<=16'd16610;
      37338:data<=16'd16512;
      37339:data<=16'd16416;
      37340:data<=16'd15816;
      37341:data<=16'd15267;
      37342:data<=16'd14078;
      37343:data<=16'd13467;
      37344:data<=16'd13085;
      37345:data<=16'd11881;
      37346:data<=16'd11549;
      37347:data<=16'd12555;
      37348:data<=16'd13535;
      37349:data<=16'd13315;
      37350:data<=16'd12125;
      37351:data<=16'd11361;
      37352:data<=16'd10988;
      37353:data<=16'd10672;
      37354:data<=16'd10129;
      37355:data<=16'd8992;
      37356:data<=16'd8698;
      37357:data<=16'd8839;
      37358:data<=16'd7858;
      37359:data<=16'd7770;
      37360:data<=16'd9357;
      37361:data<=16'd9884;
      37362:data<=16'd8915;
      37363:data<=16'd8807;
      37364:data<=16'd8975;
      37365:data<=16'd7696;
      37366:data<=16'd7257;
      37367:data<=16'd7383;
      37368:data<=16'd6390;
      37369:data<=16'd6643;
      37370:data<=16'd5808;
      37371:data<=16'd4940;
      37372:data<=16'd8322;
      37373:data<=16'd3838;
      37374:data<=-16'd9480;
      37375:data<=-16'd12558;
      37376:data<=-16'd9450;
      37377:data<=-16'd10924;
      37378:data<=-16'd10381;
      37379:data<=-16'd9436;
      37380:data<=-16'd10701;
      37381:data<=-16'd9492;
      37382:data<=-16'd8821;
      37383:data<=-16'd9411;
      37384:data<=-16'd8243;
      37385:data<=-16'd6858;
      37386:data<=-16'd6099;
      37387:data<=-16'd6352;
      37388:data<=-16'd6636;
      37389:data<=-16'd6082;
      37390:data<=-16'd6134;
      37391:data<=-16'd5606;
      37392:data<=-16'd5256;
      37393:data<=-16'd5894;
      37394:data<=-16'd4946;
      37395:data<=-16'd4464;
      37396:data<=-16'd4670;
      37397:data<=-16'd3107;
      37398:data<=-16'd2658;
      37399:data<=-16'd3298;
      37400:data<=-16'd3046;
      37401:data<=-16'd2792;
      37402:data<=-16'd2347;
      37403:data<=-16'd2602;
      37404:data<=-16'd3015;
      37405:data<=-16'd2362;
      37406:data<=-16'd2375;
      37407:data<=-16'd2623;
      37408:data<=-16'd2751;
      37409:data<=-16'd2285;
      37410:data<=-16'd259;
      37411:data<=16'd21;
      37412:data<=-16'd757;
      37413:data<=-16'd311;
      37414:data<=-16'd801;
      37415:data<=-16'd852;
      37416:data<=-16'd914;
      37417:data<=-16'd2065;
      37418:data<=-16'd1621;
      37419:data<=-16'd1536;
      37420:data<=-16'd822;
      37421:data<=16'd164;
      37422:data<=-16'd2194;
      37423:data<=16'd3313;
      37424:data<=16'd16349;
      37425:data<=16'd19011;
      37426:data<=16'd16193;
      37427:data<=16'd16910;
      37428:data<=16'd15635;
      37429:data<=16'd14334;
      37430:data<=16'd14392;
      37431:data<=16'd13493;
      37432:data<=16'd13311;
      37433:data<=16'd12342;
      37434:data<=16'd11561;
      37435:data<=16'd12466;
      37436:data<=16'd12091;
      37437:data<=16'd11374;
      37438:data<=16'd10995;
      37439:data<=16'd10322;
      37440:data<=16'd10147;
      37441:data<=16'd9085;
      37442:data<=16'd7988;
      37443:data<=16'd7718;
      37444:data<=16'd7141;
      37445:data<=16'd7019;
      37446:data<=16'd6363;
      37447:data<=16'd6094;
      37448:data<=16'd7567;
      37449:data<=16'd7392;
      37450:data<=16'd6543;
      37451:data<=16'd6305;
      37452:data<=16'd4978;
      37453:data<=16'd4921;
      37454:data<=16'd5039;
      37455:data<=16'd3597;
      37456:data<=16'd3457;
      37457:data<=16'd3416;
      37458:data<=16'd2907;
      37459:data<=16'd2942;
      37460:data<=16'd1989;
      37461:data<=16'd1343;
      37462:data<=16'd1234;
      37463:data<=16'd796;
      37464:data<=16'd867;
      37465:data<=16'd281;
      37466:data<=-16'd2;
      37467:data<=16'd105;
      37468:data<=-16'd672;
      37469:data<=-16'd94;
      37470:data<=-16'd802;
      37471:data<=-16'd1906;
      37472:data<=16'd428;
      37473:data<=-16'd5060;
      37474:data<=-16'd18310;
      37475:data<=-16'd22383;
      37476:data<=-16'd20579;
      37477:data<=-16'd21185;
      37478:data<=-16'd19849;
      37479:data<=-16'd18541;
      37480:data<=-16'd19243;
      37481:data<=-16'd18662;
      37482:data<=-16'd17587;
      37483:data<=-16'd16812;
      37484:data<=-16'd16976;
      37485:data<=-16'd18110;
      37486:data<=-16'd17699;
      37487:data<=-16'd16768;
      37488:data<=-16'd16936;
      37489:data<=-16'd16769;
      37490:data<=-16'd16039;
      37491:data<=-16'd15579;
      37492:data<=-16'd15276;
      37493:data<=-16'd14390;
      37494:data<=-16'd13705;
      37495:data<=-16'd13664;
      37496:data<=-16'd12665;
      37497:data<=-16'd12448;
      37498:data<=-16'd13885;
      37499:data<=-16'd13723;
      37500:data<=-16'd13171;
      37501:data<=-16'd13386;
      37502:data<=-16'd12402;
      37503:data<=-16'd11897;
      37504:data<=-16'd12107;
      37505:data<=-16'd11815;
      37506:data<=-16'd11878;
      37507:data<=-16'd11025;
      37508:data<=-16'd9809;
      37509:data<=-16'd9920;
      37510:data<=-16'd10123;
      37511:data<=-16'd10525;
      37512:data<=-16'd10655;
      37513:data<=-16'd10152;
      37514:data<=-16'd10176;
      37515:data<=-16'd9495;
      37516:data<=-16'd9179;
      37517:data<=-16'd9768;
      37518:data<=-16'd9222;
      37519:data<=-16'd9326;
      37520:data<=-16'd7890;
      37521:data<=-16'd5479;
      37522:data<=-16'd8652;
      37523:data<=-16'd6869;
      37524:data<=16'd5785;
      37525:data<=16'd11532;
      37526:data<=16'd8505;
      37527:data<=16'd8246;
      37528:data<=16'd8202;
      37529:data<=16'd7189;
      37530:data<=16'd7547;
      37531:data<=16'd7154;
      37532:data<=16'd6727;
      37533:data<=16'd6687;
      37534:data<=16'd6062;
      37535:data<=16'd4849;
      37536:data<=16'd2930;
      37537:data<=16'd2300;
      37538:data<=16'd2934;
      37539:data<=16'd3081;
      37540:data<=16'd3366;
      37541:data<=16'd3060;
      37542:data<=16'd2446;
      37543:data<=16'd2475;
      37544:data<=16'd1697;
      37545:data<=16'd1571;
      37546:data<=16'd2525;
      37547:data<=16'd1477;
      37548:data<=-16'd572;
      37549:data<=-16'd1055;
      37550:data<=-16'd411;
      37551:data<=-16'd332;
      37552:data<=-16'd1213;
      37553:data<=-16'd1606;
      37554:data<=-16'd1283;
      37555:data<=-16'd651;
      37556:data<=-16'd328;
      37557:data<=-16'd860;
      37558:data<=-16'd461;
      37559:data<=-16'd637;
      37560:data<=-16'd3090;
      37561:data<=-16'd3983;
      37562:data<=-16'd3527;
      37563:data<=-16'd3365;
      37564:data<=-16'd2643;
      37565:data<=-16'd3196;
      37566:data<=-16'd2974;
      37567:data<=-16'd1492;
      37568:data<=-16'd2364;
      37569:data<=-16'd2315;
      37570:data<=-16'd2429;
      37571:data<=-16'd4027;
      37572:data<=-16'd1751;
      37573:data<=-16'd5016;
      37574:data<=-16'd17685;
      37575:data<=-16'd22944;
      37576:data<=-16'd20644;
      37577:data<=-16'd20538;
      37578:data<=-16'd19790;
      37579:data<=-16'd18128;
      37580:data<=-16'd17288;
      37581:data<=-16'd16684;
      37582:data<=-16'd16601;
      37583:data<=-16'd15203;
      37584:data<=-16'd14236;
      37585:data<=-16'd15027;
      37586:data<=-16'd14471;
      37587:data<=-16'd13688;
      37588:data<=-16'd13399;
      37589:data<=-16'd12859;
      37590:data<=-16'd13189;
      37591:data<=-16'd12519;
      37592:data<=-16'd10977;
      37593:data<=-16'd10243;
      37594:data<=-16'd9135;
      37595:data<=-16'd8581;
      37596:data<=-16'd8467;
      37597:data<=-16'd8099;
      37598:data<=-16'd8877;
      37599:data<=-16'd8893;
      37600:data<=-16'd7809;
      37601:data<=-16'd7658;
      37602:data<=-16'd7432;
      37603:data<=-16'd7022;
      37604:data<=-16'd6410;
      37605:data<=-16'd5553;
      37606:data<=-16'd5689;
      37607:data<=-16'd5515;
      37608:data<=-16'd4834;
      37609:data<=-16'd4519;
      37610:data<=-16'd4309;
      37611:data<=-16'd5206;
      37612:data<=-16'd5468;
      37613:data<=-16'd4508;
      37614:data<=-16'd4690;
      37615:data<=-16'd4335;
      37616:data<=-16'd3842;
      37617:data<=-16'd3776;
      37618:data<=-16'd2126;
      37619:data<=-16'd2443;
      37620:data<=-16'd2993;
      37621:data<=-16'd605;
      37622:data<=-16'd2032;
      37623:data<=-16'd1885;
      37624:data<=16'd8191;
      37625:data<=16'd16032;
      37626:data<=16'd15534;
      37627:data<=16'd14692;
      37628:data<=16'd14601;
      37629:data<=16'd13808;
      37630:data<=16'd13371;
      37631:data<=16'd13135;
      37632:data<=16'd13000;
      37633:data<=16'd12850;
      37634:data<=16'd12631;
      37635:data<=16'd11382;
      37636:data<=16'd9104;
      37637:data<=16'd8301;
      37638:data<=16'd8522;
      37639:data<=16'd8489;
      37640:data<=16'd9006;
      37641:data<=16'd8994;
      37642:data<=16'd8075;
      37643:data<=16'd7324;
      37644:data<=16'd6699;
      37645:data<=16'd6793;
      37646:data<=16'd7124;
      37647:data<=16'd6370;
      37648:data<=16'd5280;
      37649:data<=16'd4555;
      37650:data<=16'd4167;
      37651:data<=16'd4050;
      37652:data<=16'd4043;
      37653:data<=16'd4323;
      37654:data<=16'd4423;
      37655:data<=16'd4178;
      37656:data<=16'd4055;
      37657:data<=16'd3877;
      37658:data<=16'd3961;
      37659:data<=16'd4052;
      37660:data<=16'd3691;
      37661:data<=16'd4061;
      37662:data<=16'd4402;
      37663:data<=16'd3632;
      37664:data<=16'd3580;
      37665:data<=16'd4176;
      37666:data<=16'd4366;
      37667:data<=16'd4352;
      37668:data<=16'd3474;
      37669:data<=16'd3425;
      37670:data<=16'd4317;
      37671:data<=16'd2960;
      37672:data<=16'd3451;
      37673:data<=16'd5453;
      37674:data<=-16'd2077;
      37675:data<=-16'd13200;
      37676:data<=-16'd14207;
      37677:data<=-16'd11906;
      37678:data<=-16'd12248;
      37679:data<=-16'd10675;
      37680:data<=-16'd9656;
      37681:data<=-16'd10270;
      37682:data<=-16'd9699;
      37683:data<=-16'd9359;
      37684:data<=-16'd8510;
      37685:data<=-16'd6702;
      37686:data<=-16'd5664;
      37687:data<=-16'd4537;
      37688:data<=-16'd3917;
      37689:data<=-16'd4056;
      37690:data<=-16'd3850;
      37691:data<=-16'd4005;
      37692:data<=-16'd3544;
      37693:data<=-16'd2419;
      37694:data<=-16'd1895;
      37695:data<=-16'd1401;
      37696:data<=-16'd1926;
      37697:data<=-16'd2018;
      37698:data<=16'd452;
      37699:data<=16'd1842;
      37700:data<=16'd1395;
      37701:data<=16'd1400;
      37702:data<=16'd1600;
      37703:data<=16'd2346;
      37704:data<=16'd2543;
      37705:data<=16'd1648;
      37706:data<=16'd1783;
      37707:data<=16'd2279;
      37708:data<=16'd2055;
      37709:data<=16'd1835;
      37710:data<=16'd2535;
      37711:data<=16'd3947;
      37712:data<=16'd4052;
      37713:data<=16'd4073;
      37714:data<=16'd4890;
      37715:data<=16'd4337;
      37716:data<=16'd3985;
      37717:data<=16'd3886;
      37718:data<=16'd3532;
      37719:data<=16'd4642;
      37720:data<=16'd4168;
      37721:data<=16'd3818;
      37722:data<=16'd5239;
      37723:data<=16'd4256;
      37724:data<=16'd10208;
      37725:data<=16'd23417;
      37726:data<=16'd25872;
      37727:data<=16'd22512;
      37728:data<=16'd23531;
      37729:data<=16'd21872;
      37730:data<=16'd19845;
      37731:data<=16'd20703;
      37732:data<=16'd20331;
      37733:data<=16'd19666;
      37734:data<=16'd18164;
      37735:data<=16'd17321;
      37736:data<=16'd18838;
      37737:data<=16'd18207;
      37738:data<=16'd16845;
      37739:data<=16'd16463;
      37740:data<=16'd15315;
      37741:data<=16'd15440;
      37742:data<=16'd14886;
      37743:data<=16'd13001;
      37744:data<=16'd12880;
      37745:data<=16'd12372;
      37746:data<=16'd11956;
      37747:data<=16'd12731;
      37748:data<=16'd12333;
      37749:data<=16'd12301;
      37750:data<=16'd12486;
      37751:data<=16'd11764;
      37752:data<=16'd11602;
      37753:data<=16'd10821;
      37754:data<=16'd9953;
      37755:data<=16'd9914;
      37756:data<=16'd9494;
      37757:data<=16'd9758;
      37758:data<=16'd9589;
      37759:data<=16'd8464;
      37760:data<=16'd9148;
      37761:data<=16'd10536;
      37762:data<=16'd10740;
      37763:data<=16'd9914;
      37764:data<=16'd9189;
      37765:data<=16'd9332;
      37766:data<=16'd8473;
      37767:data<=16'd7652;
      37768:data<=16'd7548;
      37769:data<=16'd6711;
      37770:data<=16'd7324;
      37771:data<=16'd6370;
      37772:data<=16'd4508;
      37773:data<=16'd8014;
      37774:data<=16'd4532;
      37775:data<=-16'd9163;
      37776:data<=-16'd13170;
      37777:data<=-16'd10345;
      37778:data<=-16'd12137;
      37779:data<=-16'd11673;
      37780:data<=-16'd9703;
      37781:data<=-16'd10169;
      37782:data<=-16'd9682;
      37783:data<=-16'd9417;
      37784:data<=-16'd9169;
      37785:data<=-16'd7758;
      37786:data<=-16'd6802;
      37787:data<=-16'd5818;
      37788:data<=-16'd5500;
      37789:data<=-16'd5518;
      37790:data<=-16'd4757;
      37791:data<=-16'd4842;
      37792:data<=-16'd4632;
      37793:data<=-16'd3660;
      37794:data<=-16'd3557;
      37795:data<=-16'd3533;
      37796:data<=-16'd3824;
      37797:data<=-16'd3798;
      37798:data<=-16'd2470;
      37799:data<=-16'd1791;
      37800:data<=-16'd1838;
      37801:data<=-16'd2046;
      37802:data<=-16'd2127;
      37803:data<=-16'd1433;
      37804:data<=-16'd1371;
      37805:data<=-16'd1453;
      37806:data<=-16'd1560;
      37807:data<=-16'd2637;
      37808:data<=-16'd2223;
      37809:data<=-16'd1654;
      37810:data<=-16'd2262;
      37811:data<=-16'd1025;
      37812:data<=-16'd208;
      37813:data<=-16'd801;
      37814:data<=-16'd503;
      37815:data<=-16'd723;
      37816:data<=-16'd834;
      37817:data<=-16'd869;
      37818:data<=-16'd1190;
      37819:data<=-16'd284;
      37820:data<=-16'd825;
      37821:data<=-16'd805;
      37822:data<=16'd503;
      37823:data<=-16'd1366;
      37824:data<=16'd3844;
      37825:data<=16'd17086;
      37826:data<=16'd20521;
      37827:data<=16'd17846;
      37828:data<=16'd18503;
      37829:data<=16'd17020;
      37830:data<=16'd15209;
      37831:data<=16'd15001;
      37832:data<=16'd14151;
      37833:data<=16'd14049;
      37834:data<=16'd12518;
      37835:data<=16'd11423;
      37836:data<=16'd13109;
      37837:data<=16'd12659;
      37838:data<=16'd11517;
      37839:data<=16'd11524;
      37840:data<=16'd10254;
      37841:data<=16'd9512;
      37842:data<=16'd8871;
      37843:data<=16'd7774;
      37844:data<=16'd7717;
      37845:data<=16'd7128;
      37846:data<=16'd6572;
      37847:data<=16'd6296;
      37848:data<=16'd6059;
      37849:data<=16'd7632;
      37850:data<=16'd7997;
      37851:data<=16'd6526;
      37852:data<=16'd6387;
      37853:data<=16'd5868;
      37854:data<=16'd5042;
      37855:data<=16'd4880;
      37856:data<=16'd4335;
      37857:data<=16'd4258;
      37858:data<=16'd3685;
      37859:data<=16'd3130;
      37860:data<=16'd3933;
      37861:data<=16'd3601;
      37862:data<=16'd2764;
      37863:data<=16'd2159;
      37864:data<=16'd1278;
      37865:data<=16'd1656;
      37866:data<=16'd1292;
      37867:data<=16'd610;
      37868:data<=16'd1036;
      37869:data<=16'd6;
      37870:data<=16'd138;
      37871:data<=16'd285;
      37872:data<=-16'd1801;
      37873:data<=-16'd902;
      37874:data<=-16'd5248;
      37875:data<=-16'd18625;
      37876:data<=-16'd23673;
      37877:data<=-16'd20648;
      37878:data<=-16'd20735;
      37879:data<=-16'd20551;
      37880:data<=-16'd19472;
      37881:data<=-16'd18895;
      37882:data<=-16'd17819;
      37883:data<=-16'd17964;
      37884:data<=-16'd17150;
      37885:data<=-16'd16383;
      37886:data<=-16'd18114;
      37887:data<=-16'd18143;
      37888:data<=-16'd17205;
      37889:data<=-16'd17074;
      37890:data<=-16'd15913;
      37891:data<=-16'd15600;
      37892:data<=-16'd15400;
      37893:data<=-16'd14114;
      37894:data<=-16'd13828;
      37895:data<=-16'd13438;
      37896:data<=-16'd12724;
      37897:data<=-16'd12239;
      37898:data<=-16'd11913;
      37899:data<=-16'd13455;
      37900:data<=-16'd14349;
      37901:data<=-16'd13127;
      37902:data<=-16'd12975;
      37903:data<=-16'd12897;
      37904:data<=-16'd12163;
      37905:data<=-16'd11940;
      37906:data<=-16'd11256;
      37907:data<=-16'd10927;
      37908:data<=-16'd10742;
      37909:data<=-16'd9940;
      37910:data<=-16'd10505;
      37911:data<=-16'd11812;
      37912:data<=-16'd12041;
      37913:data<=-16'd11212;
      37914:data<=-16'd10248;
      37915:data<=-16'd10143;
      37916:data<=-16'd9850;
      37917:data<=-16'd9688;
      37918:data<=-16'd9723;
      37919:data<=-16'd8432;
      37920:data<=-16'd8578;
      37921:data<=-16'd8737;
      37922:data<=-16'd6783;
      37923:data<=-16'd8305;
      37924:data<=-16'd6681;
      37925:data<=16'd4672;
      37926:data<=16'd11156;
      37927:data<=16'd9206;
      37928:data<=16'd9110;
      37929:data<=16'd9141;
      37930:data<=16'd7893;
      37931:data<=16'd7609;
      37932:data<=16'd6667;
      37933:data<=16'd6357;
      37934:data<=16'd6511;
      37935:data<=16'd5676;
      37936:data<=16'd5101;
      37937:data<=16'd4059;
      37938:data<=16'd3389;
      37939:data<=16'd3742;
      37940:data<=16'd2886;
      37941:data<=16'd2340;
      37942:data<=16'd2801;
      37943:data<=16'd2449;
      37944:data<=16'd2134;
      37945:data<=16'd1741;
      37946:data<=16'd1343;
      37947:data<=16'd1701;
      37948:data<=16'd772;
      37949:data<=-16'd980;
      37950:data<=-16'd1096;
      37951:data<=-16'd641;
      37952:data<=-16'd663;
      37953:data<=-16'd591;
      37954:data<=-16'd643;
      37955:data<=-16'd813;
      37956:data<=-16'd669;
      37957:data<=-16'd987;
      37958:data<=-16'd1648;
      37959:data<=-16'd1039;
      37960:data<=-16'd467;
      37961:data<=-16'd1554;
      37962:data<=-16'd2570;
      37963:data<=-16'd3106;
      37964:data<=-16'd3544;
      37965:data<=-16'd3538;
      37966:data<=-16'd3533;
      37967:data<=-16'd2544;
      37968:data<=-16'd1638;
      37969:data<=-16'd2516;
      37970:data<=-16'd2314;
      37971:data<=-16'd2003;
      37972:data<=-16'd3010;
      37973:data<=-16'd2302;
      37974:data<=-16'd5826;
      37975:data<=-16'd17014;
      37976:data<=-16'd23755;
      37977:data<=-16'd22384;
      37978:data<=-16'd21252;
      37979:data<=-16'd21093;
      37980:data<=-16'd19465;
      37981:data<=-16'd18073;
      37982:data<=-16'd17719;
      37983:data<=-16'd17447;
      37984:data<=-16'd16556;
      37985:data<=-16'd15564;
      37986:data<=-16'd15600;
      37987:data<=-16'd16178;
      37988:data<=-16'd15929;
      37989:data<=-16'd15012;
      37990:data<=-16'd14081;
      37991:data<=-16'd12948;
      37992:data<=-16'd12357;
      37993:data<=-16'd12496;
      37994:data<=-16'd11712;
      37995:data<=-16'd10734;
      37996:data<=-16'd10666;
      37997:data<=-16'd9862;
      37998:data<=-16'd9048;
      37999:data<=-16'd9694;
      38000:data<=-16'd9988;
      38001:data<=-16'd9468;
      38002:data<=-16'd9175;
      38003:data<=-16'd8715;
      38004:data<=-16'd8140;
      38005:data<=-16'd7770;
      38006:data<=-16'd7269;
      38007:data<=-16'd6645;
      38008:data<=-16'd6175;
      38009:data<=-16'd5955;
      38010:data<=-16'd5683;
      38011:data<=-16'd5792;
      38012:data<=-16'd6916;
      38013:data<=-16'd7092;
      38014:data<=-16'd5398;
      38015:data<=-16'd4561;
      38016:data<=-16'd4934;
      38017:data<=-16'd5042;
      38018:data<=-16'd4949;
      38019:data<=-16'd4067;
      38020:data<=-16'd3570;
      38021:data<=-16'd3829;
      38022:data<=-16'd2279;
      38023:data<=-16'd2350;
      38024:data<=-16'd3177;
      38025:data<=16'd5012;
      38026:data<=16'd15339;
      38027:data<=16'd15760;
      38028:data<=16'd14088;
      38029:data<=16'd15083;
      38030:data<=16'd14019;
      38031:data<=16'd13192;
      38032:data<=16'd13347;
      38033:data<=16'd12698;
      38034:data<=16'd12367;
      38035:data<=16'd11662;
      38036:data<=16'd10812;
      38037:data<=16'd9694;
      38038:data<=16'd8106;
      38039:data<=16'd8499;
      38040:data<=16'd8686;
      38041:data<=16'd7368;
      38042:data<=16'd7592;
      38043:data<=16'd7689;
      38044:data<=16'd7172;
      38045:data<=16'd7498;
      38046:data<=16'd7007;
      38047:data<=16'd6689;
      38048:data<=16'd6422;
      38049:data<=16'd4561;
      38050:data<=16'd3494;
      38051:data<=16'd3717;
      38052:data<=16'd4084;
      38053:data<=16'd4256;
      38054:data<=16'd3594;
      38055:data<=16'd3579;
      38056:data<=16'd3905;
      38057:data<=16'd3416;
      38058:data<=16'd3792;
      38059:data<=16'd4376;
      38060:data<=16'd4140;
      38061:data<=16'd3670;
      38062:data<=16'd3207;
      38063:data<=16'd3589;
      38064:data<=16'd3471;
      38065:data<=16'd2696;
      38066:data<=16'd3269;
      38067:data<=16'd3850;
      38068:data<=16'd4246;
      38069:data<=16'd4225;
      38070:data<=16'd3447;
      38071:data<=16'd4297;
      38072:data<=16'd3515;
      38073:data<=16'd2405;
      38074:data<=16'd5256;
      38075:data<=16'd171;
      38076:data<=-16'd12260;
      38077:data<=-16'd14413;
      38078:data<=-16'd11470;
      38079:data<=-16'd12461;
      38080:data<=-16'd11518;
      38081:data<=-16'd10053;
      38082:data<=-16'd10017;
      38083:data<=-16'd9007;
      38084:data<=-16'd8651;
      38085:data<=-16'd7967;
      38086:data<=-16'd6398;
      38087:data<=-16'd5400;
      38088:data<=-16'd4426;
      38089:data<=-16'd4173;
      38090:data<=-16'd3823;
      38091:data<=-16'd2966;
      38092:data<=-16'd3128;
      38093:data<=-16'd2878;
      38094:data<=-16'd2475;
      38095:data<=-16'd2425;
      38096:data<=-16'd1447;
      38097:data<=-16'd1263;
      38098:data<=-16'd1037;
      38099:data<=16'd792;
      38100:data<=16'd1700;
      38101:data<=16'd1683;
      38102:data<=16'd1595;
      38103:data<=16'd1606;
      38104:data<=16'd2208;
      38105:data<=16'd2003;
      38106:data<=16'd2053;
      38107:data<=16'd2942;
      38108:data<=16'd2637;
      38109:data<=16'd2409;
      38110:data<=16'd2473;
      38111:data<=16'd2732;
      38112:data<=16'd4317;
      38113:data<=16'd4667;
      38114:data<=16'd4320;
      38115:data<=16'd4890;
      38116:data<=16'd4616;
      38117:data<=16'd4733;
      38118:data<=16'd4516;
      38119:data<=16'd3861;
      38120:data<=16'd4875;
      38121:data<=16'd3971;
      38122:data<=16'd3592;
      38123:data<=16'd5368;
      38124:data<=16'd4009;
      38125:data<=16'd9773;
      38126:data<=16'd23572;
      38127:data<=16'd26260;
      38128:data<=16'd22632;
      38129:data<=16'd23526;
      38130:data<=16'd22151;
      38131:data<=16'd20533;
      38132:data<=16'd20900;
      38133:data<=16'd19397;
      38134:data<=16'd18844;
      38135:data<=16'd18174;
      38136:data<=16'd17159;
      38137:data<=16'd18487;
      38138:data<=16'd18045;
      38139:data<=16'd16644;
      38140:data<=16'd16766;
      38141:data<=16'd15591;
      38142:data<=16'd14836;
      38143:data<=16'd15039;
      38144:data<=16'd14340;
      38145:data<=16'd13899;
      38146:data<=16'd13060;
      38147:data<=16'd12258;
      38148:data<=16'd12525;
      38149:data<=16'd12589;
      38150:data<=16'd12777;
      38151:data<=16'd12478;
      38152:data<=16'd11594;
      38153:data<=16'd11558;
      38154:data<=16'd11217;
      38155:data<=16'd10689;
      38156:data<=16'd10264;
      38157:data<=16'd9189;
      38158:data<=16'd8984;
      38159:data<=16'd9138;
      38160:data<=16'd8819;
      38161:data<=16'd9195;
      38162:data<=16'd9846;
      38163:data<=16'd10332;
      38164:data<=16'd9856;
      38165:data<=16'd8969;
      38166:data<=16'd8960;
      38167:data<=16'd8237;
      38168:data<=16'd8220;
      38169:data<=16'd8575;
      38170:data<=16'd6969;
      38171:data<=16'd7517;
      38172:data<=16'd7501;
      38173:data<=16'd5497;
      38174:data<=16'd8510;
      38175:data<=16'd5313;
      38176:data<=-16'd8533;
      38177:data<=-16'd13106;
      38178:data<=-16'd10151;
      38179:data<=-16'd11326;
      38180:data<=-16'd10871;
      38181:data<=-16'd9718;
      38182:data<=-16'd10172;
      38183:data<=-16'd8640;
      38184:data<=-16'd8273;
      38185:data<=-16'd8760;
      38186:data<=-16'd7630;
      38187:data<=-16'd6581;
      38188:data<=-16'd5419;
      38189:data<=-16'd5233;
      38190:data<=-16'd5501;
      38191:data<=-16'd4473;
      38192:data<=-16'd4385;
      38193:data<=-16'd4475;
      38194:data<=-16'd4085;
      38195:data<=-16'd4584;
      38196:data<=-16'd4068;
      38197:data<=-16'd3510;
      38198:data<=-16'd3946;
      38199:data<=-16'd3045;
      38200:data<=-16'd1833;
      38201:data<=-16'd1377;
      38202:data<=-16'd1139;
      38203:data<=-16'd1310;
      38204:data<=-16'd1381;
      38205:data<=-16'd1395;
      38206:data<=-16'd977;
      38207:data<=-16'd466;
      38208:data<=-16'd933;
      38209:data<=-16'd1154;
      38210:data<=-16'd1510;
      38211:data<=-16'd1600;
      38212:data<=16'd162;
      38213:data<=16'd787;
      38214:data<=16'd199;
      38215:data<=16'd523;
      38216:data<=16'd516;
      38217:data<=16'd685;
      38218:data<=16'd108;
      38219:data<=-16'd983;
      38220:data<=-16'd284;
      38221:data<=-16'd893;
      38222:data<=-16'd1151;
      38223:data<=-16'd8;
      38224:data<=-16'd1409;
      38225:data<=16'd4382;
      38226:data<=16'd17576;
      38227:data<=16'd20886;
      38228:data<=16'd18255;
      38229:data<=16'd18748;
      38230:data<=16'd17484;
      38231:data<=16'd16644;
      38232:data<=16'd16612;
      38233:data<=16'd14524;
      38234:data<=16'd14292;
      38235:data<=16'd14041;
      38236:data<=16'd12913;
      38237:data<=16'd13958;
      38238:data<=16'd13668;
      38239:data<=16'd12431;
      38240:data<=16'd12434;
      38241:data<=16'd11147;
      38242:data<=16'd9919;
      38243:data<=16'd9694;
      38244:data<=16'd9139;
      38245:data<=16'd8715;
      38246:data<=16'd7868;
      38247:data<=16'd7112;
      38248:data<=16'd6913;
      38249:data<=16'd6831;
      38250:data<=16'd7647;
      38251:data<=16'd7679;
      38252:data<=16'd6441;
      38253:data<=16'd5926;
      38254:data<=16'd5582;
      38255:data<=16'd5486;
      38256:data<=16'd5242;
      38257:data<=16'd4002;
      38258:data<=16'd3651;
      38259:data<=16'd3515;
      38260:data<=16'd2786;
      38261:data<=16'd2975;
      38262:data<=16'd3080;
      38263:data<=16'd2746;
      38264:data<=16'd2355;
      38265:data<=16'd1562;
      38266:data<=16'd1177;
      38267:data<=16'd896;
      38268:data<=16'd1061;
      38269:data<=16'd1254;
      38270:data<=16'd397;
      38271:data<=16'd822;
      38272:data<=16'd425;
      38273:data<=-16'd1359;
      38274:data<=-16'd182;
      38275:data<=-16'd4576;
      38276:data<=-16'd17159;
      38277:data<=-16'd22553;
      38278:data<=-16'd20836;
      38279:data<=-16'd20999;
      38280:data<=-16'd20434;
      38281:data<=-16'd19503;
      38282:data<=-16'd19464;
      38283:data<=-16'd18374;
      38284:data<=-16'd18010;
      38285:data<=-16'd17609;
      38286:data<=-16'd16691;
      38287:data<=-16'd17437;
      38288:data<=-16'd17785;
      38289:data<=-16'd16892;
      38290:data<=-16'd16607;
      38291:data<=-16'd16463;
      38292:data<=-16'd15593;
      38293:data<=-16'd14390;
      38294:data<=-16'd14175;
      38295:data<=-16'd14454;
      38296:data<=-16'd13805;
      38297:data<=-16'd13180;
      38298:data<=-16'd12809;
      38299:data<=-16'd12877;
      38300:data<=-16'd13684;
      38301:data<=-16'd13282;
      38302:data<=-16'd12345;
      38303:data<=-16'd12252;
      38304:data<=-16'd12016;
      38305:data<=-16'd12044;
      38306:data<=-16'd11714;
      38307:data<=-16'd10701;
      38308:data<=-16'd10540;
      38309:data<=-16'd10266;
      38310:data<=-16'd9862;
      38311:data<=-16'd10040;
      38312:data<=-16'd10261;
      38313:data<=-16'd11286;
      38314:data<=-16'd11297;
      38315:data<=-16'd9914;
      38316:data<=-16'd10100;
      38317:data<=-16'd10011;
      38318:data<=-16'd9215;
      38319:data<=-16'd9248;
      38320:data<=-16'd8601;
      38321:data<=-16'd9013;
      38322:data<=-16'd8939;
      38323:data<=-16'd6760;
      38324:data<=-16'd8273;
      38325:data<=-16'd6886;
      38326:data<=16'd4208;
      38327:data<=16'd10928;
      38328:data<=16'd9271;
      38329:data<=16'd9359;
      38330:data<=16'd9817;
      38331:data<=16'd8695;
      38332:data<=16'd8617;
      38333:data<=16'd8109;
      38334:data<=16'd7550;
      38335:data<=16'd7457;
      38336:data<=16'd6393;
      38337:data<=16'd5300;
      38338:data<=16'd4522;
      38339:data<=16'd3842;
      38340:data<=16'd3736;
      38341:data<=16'd3680;
      38342:data<=16'd3472;
      38343:data<=16'd3134;
      38344:data<=16'd3051;
      38345:data<=16'd3453;
      38346:data<=16'd3203;
      38347:data<=16'd2719;
      38348:data<=16'd2608;
      38349:data<=16'd1795;
      38350:data<=16'd664;
      38351:data<=-16'd130;
      38352:data<=-16'd534;
      38353:data<=-16'd361;
      38354:data<=-16'd334;
      38355:data<=-16'd343;
      38356:data<=-16'd335;
      38357:data<=-16'd926;
      38358:data<=-16'd1178;
      38359:data<=-16'd1077;
      38360:data<=-16'd993;
      38361:data<=-16'd845;
      38362:data<=-16'd1994;
      38363:data<=-16'd3074;
      38364:data<=-16'd2596;
      38365:data<=-16'd2698;
      38366:data<=-16'd2858;
      38367:data<=-16'd2493;
      38368:data<=-16'd2852;
      38369:data<=-16'd2594;
      38370:data<=-16'd1979;
      38371:data<=-16'd1686;
      38372:data<=-16'd1460;
      38373:data<=-16'd2449;
      38374:data<=-16'd2396;
      38375:data<=-16'd4149;
      38376:data<=-16'd14143;
      38377:data<=-16'd22692;
      38378:data<=-16'd22011;
      38379:data<=-16'd20859;
      38380:data<=-16'd20797;
      38381:data<=-16'd18900;
      38382:data<=-16'd18407;
      38383:data<=-16'd18034;
      38384:data<=-16'd16900;
      38385:data<=-16'd16446;
      38386:data<=-16'd15001;
      38387:data<=-16'd14768;
      38388:data<=-16'd16257;
      38389:data<=-16'd15355;
      38390:data<=-16'd14102;
      38391:data<=-16'd14275;
      38392:data<=-16'd13200;
      38393:data<=-16'd11935;
      38394:data<=-16'd11756;
      38395:data<=-16'd11671;
      38396:data<=-16'd11621;
      38397:data<=-16'd10795;
      38398:data<=-16'd9367;
      38399:data<=-16'd9412;
      38400:data<=-16'd10470;
      38401:data<=-16'd10354;
      38402:data<=-16'd9206;
      38403:data<=-16'd8587;
      38404:data<=-16'd8398;
      38405:data<=-16'd7858;
      38406:data<=-16'd7479;
      38407:data<=-16'd7210;
      38408:data<=-16'd6390;
      38409:data<=-16'd5827;
      38410:data<=-16'd5782;
      38411:data<=-16'd5063;
      38412:data<=-16'd4584;
      38413:data<=-16'd5849;
      38414:data<=-16'd6658;
      38415:data<=-16'd5870;
      38416:data<=-16'd5777;
      38417:data<=-16'd5406;
      38418:data<=-16'd4024;
      38419:data<=-16'd4410;
      38420:data<=-16'd4861;
      38421:data<=-16'd4238;
      38422:data<=-16'd4573;
      38423:data<=-16'd3260;
      38424:data<=-16'd2742;
      38425:data<=-16'd5006;
      38426:data<=16'd1371;
      38427:data<=16'd13541;
      38428:data<=16'd15429;
      38429:data<=16'd12833;
      38430:data<=16'd14342;
      38431:data<=16'd13914;
      38432:data<=16'd12601;
      38433:data<=16'd13248;
      38434:data<=16'd12684;
      38435:data<=16'd11790;
      38436:data<=16'd11163;
      38437:data<=16'd10053;
      38438:data<=16'd9171;
      38439:data<=16'd8090;
      38440:data<=16'd7877;
      38441:data<=16'd8388;
      38442:data<=16'd7741;
      38443:data<=16'd6990;
      38444:data<=16'd6792;
      38445:data<=16'd7321;
      38446:data<=16'd8003;
      38447:data<=16'd7021;
      38448:data<=16'd6514;
      38449:data<=16'd6734;
      38450:data<=16'd4969;
      38451:data<=16'd3739;
      38452:data<=16'd4202;
      38453:data<=16'd4170;
      38454:data<=16'd4027;
      38455:data<=16'd3926;
      38456:data<=16'd3964;
      38457:data<=16'd4138;
      38458:data<=16'd3518;
      38459:data<=16'd3192;
      38460:data<=16'd3683;
      38461:data<=16'd4158;
      38462:data<=16'd4150;
      38463:data<=16'd3582;
      38464:data<=16'd3607;
      38465:data<=16'd3758;
      38466:data<=16'd3489;
      38467:data<=16'd3626;
      38468:data<=16'd3330;
      38469:data<=16'd3761;
      38470:data<=16'd4582;
      38471:data<=16'd3900;
      38472:data<=16'd4499;
      38473:data<=16'd4087;
      38474:data<=16'd2930;
      38475:data<=16'd6470;
      38476:data<=16'd2641;
      38477:data<=-16'd11163;
      38478:data<=-16'd14777;
      38479:data<=-16'd10978;
      38480:data<=-16'd11866;
      38481:data<=-16'd11483;
      38482:data<=-16'd10317;
      38483:data<=-16'd10869;
      38484:data<=-16'd9690;
      38485:data<=-16'd9151;
      38486:data<=-16'd8475;
      38487:data<=-16'd6296;
      38488:data<=-16'd5623;
      38489:data<=-16'd4952;
      38490:data<=-16'd4020;
      38491:data<=-16'd3996;
      38492:data<=-16'd3375;
      38493:data<=-16'd2775;
      38494:data<=-16'd2473;
      38495:data<=-16'd2411;
      38496:data<=-16'd2635;
      38497:data<=-16'd1827;
      38498:data<=-16'd1407;
      38499:data<=-16'd1375;
      38500:data<=16'd196;
      38501:data<=16'd1283;
      38502:data<=16'd1133;
      38503:data<=16'd1260;
      38504:data<=16'd1691;
      38505:data<=16'd2017;
      38506:data<=16'd1704;
      38507:data<=16'd1371;
      38508:data<=16'd1598;
      38509:data<=16'd2079;
      38510:data<=16'd2408;
      38511:data<=16'd1650;
      38512:data<=16'd1779;
      38513:data<=16'd3430;
      38514:data<=16'd3601;
      38515:data<=16'd3582;
      38516:data<=16'd3906;
      38517:data<=16'd3874;
      38518:data<=16'd4968;
      38519:data<=16'd4005;
      38520:data<=16'd2623;
      38521:data<=16'd4247;
      38522:data<=16'd3542;
      38523:data<=16'd3448;
      38524:data<=16'd5083;
      38525:data<=16'd2933;
      38526:data<=16'd8643;
      38527:data<=16'd22016;
      38528:data<=16'd24783;
      38529:data<=16'd22336;
      38530:data<=16'd22838;
      38531:data<=16'd21215;
      38532:data<=16'd20503;
      38533:data<=16'd20610;
      38534:data<=16'd19240;
      38535:data<=16'd19024;
      38536:data<=16'd17358;
      38537:data<=16'd16208;
      38538:data<=16'd17989;
      38539:data<=16'd17379;
      38540:data<=16'd16019;
      38541:data<=16'd16151;
      38542:data<=16'd15227;
      38543:data<=16'd14512;
      38544:data<=16'd13932;
      38545:data<=16'd13286;
      38546:data<=16'd13183;
      38547:data<=16'd12035;
      38548:data<=16'd11414;
      38549:data<=16'd11518;
      38550:data<=16'd11024;
      38551:data<=16'd11752;
      38552:data<=16'd12070;
      38553:data<=16'd11129;
      38554:data<=16'd11027;
      38555:data<=16'd10352;
      38556:data<=16'd9673;
      38557:data<=16'd10072;
      38558:data<=16'd9411;
      38559:data<=16'd8384;
      38560:data<=16'd8194;
      38561:data<=16'd8194;
      38562:data<=16'd8334;
      38563:data<=16'd8918;
      38564:data<=16'd9561;
      38565:data<=16'd8851;
      38566:data<=16'd8258;
      38567:data<=16'd8486;
      38568:data<=16'd6992;
      38569:data<=16'd6607;
      38570:data<=16'd7521;
      38571:data<=16'd6253;
      38572:data<=16'd6479;
      38573:data<=16'd6067;
      38574:data<=16'd3767;
      38575:data<=16'd6358;
      38576:data<=16'd3841;
      38577:data<=-16'd8473;
      38578:data<=-16'd13238;
      38579:data<=-16'd11013;
      38580:data<=-16'd11617;
      38581:data<=-16'd11435;
      38582:data<=-16'd11200;
      38583:data<=-16'd11373;
      38584:data<=-16'd9897;
      38585:data<=-16'd10031;
      38586:data<=-16'd9935;
      38587:data<=-16'd8432;
      38588:data<=-16'd7671;
      38589:data<=-16'd5982;
      38590:data<=-16'd5233;
      38591:data<=-16'd5791;
      38592:data<=-16'd5145;
      38593:data<=-16'd5576;
      38594:data<=-16'd5814;
      38595:data<=-16'd4648;
      38596:data<=-16'd4945;
      38597:data<=-16'd4846;
      38598:data<=-16'd4287;
      38599:data<=-16'd4825;
      38600:data<=-16'd3826;
      38601:data<=-16'd2185;
      38602:data<=-16'd1718;
      38603:data<=-16'd1486;
      38604:data<=-16'd1812;
      38605:data<=-16'd2138;
      38606:data<=-16'd2146;
      38607:data<=-16'd2322;
      38608:data<=-16'd1855;
      38609:data<=-16'd1466;
      38610:data<=-16'd2156;
      38611:data<=-16'd2834;
      38612:data<=-16'd2334;
      38613:data<=-16'd1204;
      38614:data<=-16'd704;
      38615:data<=-16'd505;
      38616:data<=-16'd526;
      38617:data<=-16'd476;
      38618:data<=16'd355;
      38619:data<=16'd73;
      38620:data<=-16'd350;
      38621:data<=16'd24;
      38622:data<=-16'd1585;
      38623:data<=-16'd1313;
      38624:data<=16'd412;
      38625:data<=-16'd1431;
      38626:data<=16'd3706;
      38627:data<=16'd16424;
      38628:data<=16'd20236;
      38629:data<=16'd18301;
      38630:data<=16'd18760;
      38631:data<=16'd17552;
      38632:data<=16'd16615;
      38633:data<=16'd16433;
      38634:data<=16'd14454;
      38635:data<=16'd13759;
      38636:data<=16'd13130;
      38637:data<=16'd11997;
      38638:data<=16'd12936;
      38639:data<=16'd12972;
      38640:data<=16'd11618;
      38641:data<=16'd11260;
      38642:data<=16'd10910;
      38643:data<=16'd10172;
      38644:data<=16'd9300;
      38645:data<=16'd8690;
      38646:data<=16'd8313;
      38647:data<=16'd7354;
      38648:data<=16'd6978;
      38649:data<=16'd7012;
      38650:data<=16'd6734;
      38651:data<=16'd7312;
      38652:data<=16'd7568;
      38653:data<=16'd7010;
      38654:data<=16'd6570;
      38655:data<=16'd5541;
      38656:data<=16'd5086;
      38657:data<=16'd5407;
      38658:data<=16'd4770;
      38659:data<=16'd3999;
      38660:data<=16'd3773;
      38661:data<=16'd4052;
      38662:data<=16'd4281;
      38663:data<=16'd3450;
      38664:data<=16'd2951;
      38665:data<=16'd2817;
      38666:data<=16'd2311;
      38667:data<=16'd2332;
      38668:data<=16'd1707;
      38669:data<=16'd931;
      38670:data<=16'd996;
      38671:data<=16'd500;
      38672:data<=16'd537;
      38673:data<=-16'd197;
      38674:data<=-16'd1712;
      38675:data<=-16'd490;
      38676:data<=-16'd4411;
      38677:data<=-16'd16133;
      38678:data<=-16'd21828;
      38679:data<=-16'd20765;
      38680:data<=-16'd20906;
      38681:data<=-16'd20395;
      38682:data<=-16'd19516;
      38683:data<=-16'd19411;
      38684:data<=-16'd18380;
      38685:data<=-16'd17778;
      38686:data<=-16'd16932;
      38687:data<=-16'd15787;
      38688:data<=-16'd16606;
      38689:data<=-16'd17105;
      38690:data<=-16'd15979;
      38691:data<=-16'd15434;
      38692:data<=-16'd15479;
      38693:data<=-16'd14859;
      38694:data<=-16'd13841;
      38695:data<=-16'd13729;
      38696:data<=-16'd13797;
      38697:data<=-16'd12994;
      38698:data<=-16'd12552;
      38699:data<=-16'd12192;
      38700:data<=-16'd11906;
      38701:data<=-16'd12751;
      38702:data<=-16'd12897;
      38703:data<=-16'd12251;
      38704:data<=-16'd12237;
      38705:data<=-16'd11734;
      38706:data<=-16'd11068;
      38707:data<=-16'd11062;
      38708:data<=-16'd10828;
      38709:data<=-16'd10170;
      38710:data<=-16'd9794;
      38711:data<=-16'd10207;
      38712:data<=-16'd10201;
      38713:data<=-16'd10073;
      38714:data<=-16'd11195;
      38715:data<=-16'd10795;
      38716:data<=-16'd9552;
      38717:data<=-16'd10493;
      38718:data<=-16'd10245;
      38719:data<=-16'd8922;
      38720:data<=-16'd8722;
      38721:data<=-16'd7692;
      38722:data<=-16'd8041;
      38723:data<=-16'd8552;
      38724:data<=-16'd6422;
      38725:data<=-16'd7623;
      38726:data<=-16'd7655;
      38727:data<=16'd2035;
      38728:data<=16'd10401;
      38729:data<=16'd10154;
      38730:data<=16'd9263;
      38731:data<=16'd9691;
      38732:data<=16'd9266;
      38733:data<=16'd9025;
      38734:data<=16'd8643;
      38735:data<=16'd7623;
      38736:data<=16'd6545;
      38737:data<=16'd6070;
      38738:data<=16'd5844;
      38739:data<=16'd4652;
      38740:data<=16'd3462;
      38741:data<=16'd3221;
      38742:data<=16'd2783;
      38743:data<=16'd2203;
      38744:data<=16'd2182;
      38745:data<=16'd2519;
      38746:data<=16'd2690;
      38747:data<=16'd2061;
      38748:data<=16'd1538;
      38749:data<=16'd1873;
      38750:data<=16'd1522;
      38751:data<=16'd337;
      38752:data<=-16'd353;
      38753:data<=-16'd773;
      38754:data<=-16'd1266;
      38755:data<=-16'd1571;
      38756:data<=-16'd1350;
      38757:data<=-16'd604;
      38758:data<=-16'd464;
      38759:data<=-16'd930;
      38760:data<=-16'd773;
      38761:data<=-16'd221;
      38762:data<=16'd38;
      38763:data<=-16'd607;
      38764:data<=-16'd1977;
      38765:data<=-16'd2525;
      38766:data<=-16'd2447;
      38767:data<=-16'd2514;
      38768:data<=-16'd2276;
      38769:data<=-16'd2137;
      38770:data<=-16'd2202;
      38771:data<=-16'd2453;
      38772:data<=-16'd2534;
      38773:data<=-16'd1709;
      38774:data<=-16'd2026;
      38775:data<=-16'd2626;
      38776:data<=-16'd2937;
      38777:data<=-16'd10325;
      38778:data<=-16'd21076;
      38779:data<=-16'd22723;
      38780:data<=-16'd20272;
      38781:data<=-16'd20741;
      38782:data<=-16'd19848;
      38783:data<=-16'd18331;
      38784:data<=-16'd18026;
      38785:data<=-16'd17062;
      38786:data<=-16'd15948;
      38787:data<=-16'd14666;
      38788:data<=-16'd14231;
      38789:data<=-16'd15164;
      38790:data<=-16'd14801;
      38791:data<=-16'd13784;
      38792:data<=-16'd13123;
      38793:data<=-16'd11932;
      38794:data<=-16'd11198;
      38795:data<=-16'd10781;
      38796:data<=-16'd10392;
      38797:data<=-16'd10111;
      38798:data<=-16'd8934;
      38799:data<=-16'd8238;
      38800:data<=-16'd8804;
      38801:data<=-16'd9368;
      38802:data<=-16'd9741;
      38803:data<=-16'd9359;
      38804:data<=-16'd8507;
      38805:data<=-16'd7711;
      38806:data<=-16'd6666;
      38807:data<=-16'd6566;
      38808:data<=-16'd6680;
      38809:data<=-16'd5797;
      38810:data<=-16'd5332;
      38811:data<=-16'd4908;
      38812:data<=-16'd4410;
      38813:data<=-16'd5171;
      38814:data<=-16'd6422;
      38815:data<=-16'd6707;
      38816:data<=-16'd5697;
      38817:data<=-16'd5172;
      38818:data<=-16'd5206;
      38819:data<=-16'd4273;
      38820:data<=-16'd4443;
      38821:data<=-16'd4153;
      38822:data<=-16'd2209;
      38823:data<=-16'd2963;
      38824:data<=-16'd2312;
      38825:data<=-16'd619;
      38826:data<=-16'd4291;
      38827:data<=-16'd461;
      38828:data<=16'd12901;
      38829:data<=16'd16319;
      38830:data<=16'd13621;
      38831:data<=16'd15224;
      38832:data<=16'd14681;
      38833:data<=16'd13335;
      38834:data<=16'd14061;
      38835:data<=16'd13227;
      38836:data<=16'd12634;
      38837:data<=16'd12493;
      38838:data<=16'd10977;
      38839:data<=16'd9259;
      38840:data<=16'd8173;
      38841:data<=16'd8493;
      38842:data<=16'd8586;
      38843:data<=16'd7608;
      38844:data<=16'd7429;
      38845:data<=16'd6993;
      38846:data<=16'd6857;
      38847:data<=16'd7589;
      38848:data<=16'd6815;
      38849:data<=16'd6610;
      38850:data<=16'd7168;
      38851:data<=16'd5623;
      38852:data<=16'd4494;
      38853:data<=16'd4570;
      38854:data<=16'd4276;
      38855:data<=16'd4364;
      38856:data<=16'd4115;
      38857:data<=16'd3680;
      38858:data<=16'd4079;
      38859:data<=16'd4458;
      38860:data<=16'd4432;
      38861:data<=16'd4012;
      38862:data<=16'd4090;
      38863:data<=16'd4801;
      38864:data<=16'd4969;
      38865:data<=16'd4957;
      38866:data<=16'd4247;
      38867:data<=16'd3594;
      38868:data<=16'd4178;
      38869:data<=16'd3638;
      38870:data<=16'd3342;
      38871:data<=16'd3930;
      38872:data<=16'd3204;
      38873:data<=16'd4018;
      38874:data<=16'd3711;
      38875:data<=16'd2132;
      38876:data<=16'd5927;
      38877:data<=16'd3192;
      38878:data<=-16'd9969;
      38879:data<=-16'd13714;
      38880:data<=-16'd10731;
      38881:data<=-16'd12460;
      38882:data<=-16'd11764;
      38883:data<=-16'd9743;
      38884:data<=-16'd10154;
      38885:data<=-16'd9197;
      38886:data<=-16'd8860;
      38887:data<=-16'd8672;
      38888:data<=-16'd6664;
      38889:data<=-16'd5133;
      38890:data<=-16'd4020;
      38891:data<=-16'd3782;
      38892:data<=-16'd3469;
      38893:data<=-16'd2309;
      38894:data<=-16'd2846;
      38895:data<=-16'd2108;
      38896:data<=16'd390;
      38897:data<=16'd406;
      38898:data<=16'd496;
      38899:data<=16'd1139;
      38900:data<=16'd628;
      38901:data<=16'd1750;
      38902:data<=16'd3263;
      38903:data<=16'd3357;
      38904:data<=16'd3395;
      38905:data<=16'd3018;
      38906:data<=16'd2860;
      38907:data<=16'd3265;
      38908:data<=16'd3043;
      38909:data<=16'd2751;
      38910:data<=16'd3122;
      38911:data<=16'd3416;
      38912:data<=16'd2669;
      38913:data<=16'd2663;
      38914:data<=16'd4244;
      38915:data<=16'd4570;
      38916:data<=16'd4590;
      38917:data<=16'd5172;
      38918:data<=16'd4508;
      38919:data<=16'd4699;
      38920:data<=16'd5248;
      38921:data<=16'd4901;
      38922:data<=16'd5118;
      38923:data<=16'd4027;
      38924:data<=16'd4191;
      38925:data<=16'd5580;
      38926:data<=16'd3629;
      38927:data<=16'd8247;
      38928:data<=16'd19722;
      38929:data<=16'd21969;
      38930:data<=16'd19637;
      38931:data<=16'd20862;
      38932:data<=16'd19910;
      38933:data<=16'd18424;
      38934:data<=16'd17914;
      38935:data<=16'd16665;
      38936:data<=16'd16782;
      38937:data<=16'd16257;
      38938:data<=16'd15402;
      38939:data<=16'd15907;
      38940:data<=16'd15121;
      38941:data<=16'd14616;
      38942:data<=16'd14516;
      38943:data<=16'd13112;
      38944:data<=16'd13030;
      38945:data<=16'd13036;
      38946:data<=16'd11934;
      38947:data<=16'd11479;
      38948:data<=16'd10560;
      38949:data<=16'd10049;
      38950:data<=16'd10454;
      38951:data<=16'd10314;
      38952:data<=16'd10745;
      38953:data<=16'd10824;
      38954:data<=16'd10117;
      38955:data<=16'd10336;
      38956:data<=16'd9964;
      38957:data<=16'd9004;
      38958:data<=16'd8886;
      38959:data<=16'd8526;
      38960:data<=16'd7661;
      38961:data<=16'd6783;
      38962:data<=16'd6614;
      38963:data<=16'd7356;
      38964:data<=16'd8028;
      38965:data<=16'd8404;
      38966:data<=16'd7788;
      38967:data<=16'd7101;
      38968:data<=16'd7511;
      38969:data<=16'd6754;
      38970:data<=16'd5780;
      38971:data<=16'd5567;
      38972:data<=16'd4402;
      38973:data<=16'd4717;
      38974:data<=16'd4640;
      38975:data<=16'd2695;
      38976:data<=16'd4576;
      38977:data<=16'd3189;
      38978:data<=-16'd6930;
      38979:data<=-16'd11752;
      38980:data<=-16'd9586;
      38981:data<=-16'd10181;
      38982:data<=-16'd10669;
      38983:data<=-16'd9580;
      38984:data<=-16'd9674;
      38985:data<=-16'd9138;
      38986:data<=-16'd8664;
      38987:data<=-16'd9063;
      38988:data<=-16'd8323;
      38989:data<=-16'd6496;
      38990:data<=-16'd5160;
      38991:data<=-16'd5130;
      38992:data<=-16'd4908;
      38993:data<=-16'd4267;
      38994:data<=-16'd4878;
      38995:data<=-16'd5074;
      38996:data<=-16'd4658;
      38997:data<=-16'd5098;
      38998:data<=-16'd4470;
      38999:data<=-16'd3991;
      39000:data<=-16'd5180;
      39001:data<=-16'd4535;
      39002:data<=-16'd2381;
      39003:data<=-16'd1635;
      39004:data<=-16'd1568;
      39005:data<=-16'd1574;
      39006:data<=-16'd2047;
      39007:data<=-16'd2579;
      39008:data<=-16'd2716;
      39009:data<=-16'd2808;
      39010:data<=-16'd2966;
      39011:data<=-16'd2657;
      39012:data<=-16'd2887;
      39013:data<=-16'd3277;
      39014:data<=-16'd1865;
      39015:data<=-16'd652;
      39016:data<=-16'd757;
      39017:data<=-16'd626;
      39018:data<=-16'd940;
      39019:data<=-16'd1143;
      39020:data<=-16'd672;
      39021:data<=-16'd597;
      39022:data<=-16'd438;
      39023:data<=-16'd817;
      39024:data<=-16'd889;
      39025:data<=-16'd224;
      39026:data<=-16'd1154;
      39027:data<=16'd2645;
      39028:data<=16'd13006;
      39029:data<=16'd17132;
      39030:data<=16'd14965;
      39031:data<=16'd15039;
      39032:data<=16'd14509;
      39033:data<=16'd13148;
      39034:data<=16'd13065;
      39035:data<=16'd11846;
      39036:data<=16'd11133;
      39037:data<=16'd11095;
      39038:data<=16'd10084;
      39039:data<=16'd10314;
      39040:data<=16'd10936;
      39041:data<=16'd10443;
      39042:data<=16'd9814;
      39043:data<=16'd8775;
      39044:data<=16'd8199;
      39045:data<=16'd8251;
      39046:data<=16'd7782;
      39047:data<=16'd7474;
      39048:data<=16'd6951;
      39049:data<=16'd6043;
      39050:data<=16'd5850;
      39051:data<=16'd6260;
      39052:data<=16'd7116;
      39053:data<=16'd7224;
      39054:data<=16'd6269;
      39055:data<=16'd5993;
      39056:data<=16'd5476;
      39057:data<=16'd4772;
      39058:data<=16'd5473;
      39059:data<=16'd5435;
      39060:data<=16'd4226;
      39061:data<=16'd3808;
      39062:data<=16'd3736;
      39063:data<=16'd3657;
      39064:data<=16'd3319;
      39065:data<=16'd2625;
      39066:data<=16'd2452;
      39067:data<=16'd2394;
      39068:data<=16'd2094;
      39069:data<=16'd1492;
      39070:data<=16'd664;
      39071:data<=16'd509;
      39072:data<=16'd176;
      39073:data<=-16'd426;
      39074:data<=-16'd381;
      39075:data<=-16'd440;
      39076:data<=-16'd111;
      39077:data<=-16'd2755;
      39078:data<=-16'd11759;
      39079:data<=-16'd18316;
      39080:data<=-16'd17676;
      39081:data<=-16'd16792;
      39082:data<=-16'd16656;
      39083:data<=-16'd15752;
      39084:data<=-16'd15443;
      39085:data<=-16'd14434;
      39086:data<=-16'd13576;
      39087:data<=-16'd13718;
      39088:data<=-16'd13397;
      39089:data<=-16'd13863;
      39090:data<=-16'd14559;
      39091:data<=-16'd13940;
      39092:data<=-16'd13383;
      39093:data<=-16'd12925;
      39094:data<=-16'd12413;
      39095:data<=-16'd12087;
      39096:data<=-16'd11511;
      39097:data<=-16'd11435;
      39098:data<=-16'd11398;
      39099:data<=-16'd10724;
      39100:data<=-16'd10249;
      39101:data<=-16'd10405;
      39102:data<=-16'd11626;
      39103:data<=-16'd12155;
      39104:data<=-16'd10850;
      39105:data<=-16'd10487;
      39106:data<=-16'd10684;
      39107:data<=-16'd10026;
      39108:data<=-16'd9902;
      39109:data<=-16'd9582;
      39110:data<=-16'd9221;
      39111:data<=-16'd9435;
      39112:data<=-16'd8593;
      39113:data<=-16'd8062;
      39114:data<=-16'd9145;
      39115:data<=-16'd10120;
      39116:data<=-16'd9900;
      39117:data<=-16'd8613;
      39118:data<=-16'd7987;
      39119:data<=-16'd7850;
      39120:data<=-16'd7037;
      39121:data<=-16'd7069;
      39122:data<=-16'd6572;
      39123:data<=-16'd5369;
      39124:data<=-16'd5864;
      39125:data<=-16'd5485;
      39126:data<=-16'd6024;
      39127:data<=-16'd8028;
      39128:data<=-16'd1817;
      39129:data<=16'd8146;
      39130:data<=16'd9289;
      39131:data<=16'd7297;
      39132:data<=16'd8047;
      39133:data<=16'd7406;
      39134:data<=16'd6150;
      39135:data<=16'd6217;
      39136:data<=16'd5927;
      39137:data<=16'd5406;
      39138:data<=16'd5838;
      39139:data<=16'd5633;
      39140:data<=16'd3260;
      39141:data<=16'd2117;
      39142:data<=16'd3407;
      39143:data<=16'd3287;
      39144:data<=16'd2416;
      39145:data<=16'd2578;
      39146:data<=16'd2461;
      39147:data<=16'd2473;
      39148:data<=16'd2049;
      39149:data<=16'd1221;
      39150:data<=16'd1994;
      39151:data<=16'd2115;
      39152:data<=16'd394;
      39153:data<=-16'd481;
      39154:data<=-16'd473;
      39155:data<=-16'd344;
      39156:data<=-16'd277;
      39157:data<=-16'd561;
      39158:data<=-16'd508;
      39159:data<=-16'd458;
      39160:data<=-16'd388;
      39161:data<=-16'd118;
      39162:data<=-16'd646;
      39163:data<=-16'd904;
      39164:data<=-16'd1096;
      39165:data<=-16'd2605;
      39166:data<=-16'd3283;
      39167:data<=-16'd3112;
      39168:data<=-16'd3579;
      39169:data<=-16'd3509;
      39170:data<=-16'd3254;
      39171:data<=-16'd3087;
      39172:data<=-16'd2957;
      39173:data<=-16'd3237;
      39174:data<=-16'd2554;
      39175:data<=-16'd2861;
      39176:data<=-16'd3738;
      39177:data<=-16'd2422;
      39178:data<=-16'd7354;
      39179:data<=-16'd18274;
      39180:data<=-16'd20410;
      39181:data<=-16'd17223;
      39182:data<=-16'd17835;
      39183:data<=-16'd17042;
      39184:data<=-16'd15144;
      39185:data<=-16'd14806;
      39186:data<=-16'd13490;
      39187:data<=-16'd13160;
      39188:data<=-16'd13712;
      39189:data<=-16'd13259;
      39190:data<=-16'd13347;
      39191:data<=-16'd13200;
      39192:data<=-16'd12768;
      39193:data<=-16'd12392;
      39194:data<=-16'd10894;
      39195:data<=-16'd10076;
      39196:data<=-16'd10050;
      39197:data<=-16'd9497;
      39198:data<=-16'd9125;
      39199:data<=-16'd8252;
      39200:data<=-16'd7682;
      39201:data<=-16'd8384;
      39202:data<=-16'd8654;
      39203:data<=-16'd8487;
      39204:data<=-16'd8096;
      39205:data<=-16'd7685;
      39206:data<=-16'd7623;
      39207:data<=-16'd6837;
      39208:data<=-16'd6460;
      39209:data<=-16'd6375;
      39210:data<=-16'd5157;
      39211:data<=-16'd4918;
      39212:data<=-16'd4795;
      39213:data<=-16'd3571;
      39214:data<=-16'd4050;
      39215:data<=-16'd5268;
      39216:data<=-16'd5134;
      39217:data<=-16'd4402;
      39218:data<=-16'd4074;
      39219:data<=-16'd4246;
      39220:data<=-16'd3348;
      39221:data<=-16'd2555;
      39222:data<=-16'd2525;
      39223:data<=-16'd1377;
      39224:data<=-16'd1448;
      39225:data<=-16'd1340;
      39226:data<=-16'd619;
      39227:data<=-16'd3853;
      39228:data<=-16'd820;
      39229:data<=16'd11198;
      39230:data<=16'd14281;
      39231:data<=16'd11013;
      39232:data<=16'd12411;
      39233:data<=16'd12369;
      39234:data<=16'd11220;
      39235:data<=16'd11579;
      39236:data<=16'd10198;
      39237:data<=16'd10055;
      39238:data<=16'd11098;
      39239:data<=16'd10141;
      39240:data<=16'd8492;
      39241:data<=16'd7401;
      39242:data<=16'd7764;
      39243:data<=16'd7485;
      39244:data<=16'd5736;
      39245:data<=16'd5997;
      39246:data<=16'd6619;
      39247:data<=16'd6448;
      39248:data<=16'd6946;
      39249:data<=16'd5994;
      39250:data<=16'd5274;
      39251:data<=16'd6150;
      39252:data<=16'd5380;
      39253:data<=16'd4027;
      39254:data<=16'd3685;
      39255:data<=16'd3650;
      39256:data<=16'd3897;
      39257:data<=16'd3844;
      39258:data<=16'd3980;
      39259:data<=16'd4100;
      39260:data<=16'd3623;
      39261:data<=16'd3586;
      39262:data<=16'd3301;
      39263:data<=16'd3043;
      39264:data<=16'd3410;
      39265:data<=16'd3165;
      39266:data<=16'd3254;
      39267:data<=16'd3224;
      39268:data<=16'd2513;
      39269:data<=16'd2819;
      39270:data<=16'd2786;
      39271:data<=16'd2664;
      39272:data<=16'd2924;
      39273:data<=16'd1988;
      39274:data<=16'd2379;
      39275:data<=16'd2481;
      39276:data<=16'd1635;
      39277:data<=16'd4589;
      39278:data<=16'd2475;
      39279:data<=-16'd8117;
      39280:data<=-16'd11828;
      39281:data<=-16'd9165;
      39282:data<=-16'd9514;
      39283:data<=-16'd9307;
      39284:data<=-16'd8352;
      39285:data<=-16'd8496;
      39286:data<=-16'd7430;
      39287:data<=-16'd6858;
      39288:data<=-16'd7248;
      39289:data<=-16'd6417;
      39290:data<=-16'd4381;
      39291:data<=-16'd2767;
      39292:data<=-16'd3207;
      39293:data<=-16'd3366;
      39294:data<=-16'd1865;
      39295:data<=-16'd1533;
      39296:data<=-16'd1745;
      39297:data<=-16'd1712;
      39298:data<=-16'd2396;
      39299:data<=-16'd1783;
      39300:data<=-16'd690;
      39301:data<=-16'd1239;
      39302:data<=-16'd802;
      39303:data<=16'd1121;
      39304:data<=16'd1780;
      39305:data<=16'd1569;
      39306:data<=16'd1903;
      39307:data<=16'd1877;
      39308:data<=16'd1480;
      39309:data<=16'd1868;
      39310:data<=16'd2006;
      39311:data<=16'd1820;
      39312:data<=16'd2487;
      39313:data<=16'd2594;
      39314:data<=16'd2745;
      39315:data<=16'd4264;
      39316:data<=16'd4746;
      39317:data<=16'd4446;
      39318:data<=16'd4714;
      39319:data<=16'd4564;
      39320:data<=16'd4713;
      39321:data<=16'd4840;
      39322:data<=16'd4696;
      39323:data<=16'd4981;
      39324:data<=16'd4234;
      39325:data<=16'd4570;
      39326:data<=16'd5491;
      39327:data<=16'd3489;
      39328:data<=16'd7404;
      39329:data<=16'd18645;
      39330:data<=16'd22166;
      39331:data<=16'd19130;
      39332:data<=16'd19165;
      39333:data<=16'd19011;
      39334:data<=16'd17805;
      39335:data<=16'd17434;
      39336:data<=16'd16289;
      39337:data<=16'd15793;
      39338:data<=16'd15831;
      39339:data<=16'd15394;
      39340:data<=16'd15599;
      39341:data<=16'd15339;
      39342:data<=16'd14945;
      39343:data<=16'd14891;
      39344:data<=16'd13544;
      39345:data<=16'd12574;
      39346:data<=16'd12605;
      39347:data<=16'd12046;
      39348:data<=16'd11747;
      39349:data<=16'd11444;
      39350:data<=16'd10698;
      39351:data<=16'd10499;
      39352:data<=16'd10546;
      39353:data<=16'd11012;
      39354:data<=16'd11314;
      39355:data<=16'd10311;
      39356:data<=16'd9664;
      39357:data<=16'd9815;
      39358:data<=16'd9415;
      39359:data<=16'd8734;
      39360:data<=16'd7993;
      39361:data<=16'd7213;
      39362:data<=16'd6742;
      39363:data<=16'd6328;
      39364:data<=16'd6176;
      39365:data<=16'd6987;
      39366:data<=16'd8088;
      39367:data<=16'd7808;
      39368:data<=16'd6863;
      39369:data<=16'd6570;
      39370:data<=16'd5902;
      39371:data<=16'd5536;
      39372:data<=16'd5580;
      39373:data<=16'd4261;
      39374:data<=16'd3756;
      39375:data<=16'd3709;
      39376:data<=16'd2760;
      39377:data<=16'd4608;
      39378:data<=16'd3412;
      39379:data<=-16'd5862;
      39380:data<=-16'd11142;
      39381:data<=-16'd9774;
      39382:data<=-16'd10260;
      39383:data<=-16'd10451;
      39384:data<=-16'd9456;
      39385:data<=-16'd9919;
      39386:data<=-16'd9351;
      39387:data<=-16'd8628;
      39388:data<=-16'd9004;
      39389:data<=-16'd8445;
      39390:data<=-16'd7130;
      39391:data<=-16'd5844;
      39392:data<=-16'd5547;
      39393:data<=-16'd5727;
      39394:data<=-16'd5121;
      39395:data<=-16'd5357;
      39396:data<=-16'd5638;
      39397:data<=-16'd5256;
      39398:data<=-16'd6050;
      39399:data<=-16'd5883;
      39400:data<=-16'd4968;
      39401:data<=-16'd5670;
      39402:data<=-16'd5151;
      39403:data<=-16'd3573;
      39404:data<=-16'd3265;
      39405:data<=-16'd2913;
      39406:data<=-16'd2837;
      39407:data<=-16'd3322;
      39408:data<=-16'd3275;
      39409:data<=-16'd3145;
      39410:data<=-16'd3030;
      39411:data<=-16'd2951;
      39412:data<=-16'd2993;
      39413:data<=-16'd3101;
      39414:data<=-16'd3060;
      39415:data<=-16'd1814;
      39416:data<=-16'd638;
      39417:data<=-16'd661;
      39418:data<=-16'd553;
      39419:data<=-16'd638;
      39420:data<=-16'd479;
      39421:data<=16'd103;
      39422:data<=-16'd537;
      39423:data<=-16'd873;
      39424:data<=-16'd549;
      39425:data<=-16'd599;
      39426:data<=-16'd520;
      39427:data<=-16'd1343;
      39428:data<=16'd1468;
      39429:data<=16'd10520;
      39430:data<=16'd15606;
      39431:data<=16'd14393;
      39432:data<=16'd13867;
      39433:data<=16'd13389;
      39434:data<=16'd12586;
      39435:data<=16'd12469;
      39436:data<=16'd11262;
      39437:data<=16'd10533;
      39438:data<=16'd10683;
      39439:data<=16'd10096;
      39440:data<=16'd9917;
      39441:data<=16'd10454;
      39442:data<=16'd10675;
      39443:data<=16'd9815;
      39444:data<=16'd8583;
      39445:data<=16'd8411;
      39446:data<=16'd8147;
      39447:data<=16'd7568;
      39448:data<=16'd7518;
      39449:data<=16'd7009;
      39450:data<=16'd6410;
      39451:data<=16'd6009;
      39452:data<=16'd5865;
      39453:data<=16'd6840;
      39454:data<=16'd7198;
      39455:data<=16'd6508;
      39456:data<=16'd6172;
      39457:data<=16'd5557;
      39458:data<=16'd5172;
      39459:data<=16'd4940;
      39460:data<=16'd3977;
      39461:data<=16'd3682;
      39462:data<=16'd3727;
      39463:data<=16'd3307;
      39464:data<=16'd2795;
      39465:data<=16'd1844;
      39466:data<=16'd1597;
      39467:data<=16'd1742;
      39468:data<=16'd999;
      39469:data<=16'd822;
      39470:data<=16'd520;
      39471:data<=-16'd284;
      39472:data<=16'd96;
      39473:data<=-16'd67;
      39474:data<=-16'd842;
      39475:data<=-16'd608;
      39476:data<=-16'd726;
      39477:data<=-16'd779;
      39478:data<=-16'd2469;
      39479:data<=-16'd9881;
      39480:data<=-16'd17578;
      39481:data<=-16'd18577;
      39482:data<=-16'd16857;
      39483:data<=-16'd16780;
      39484:data<=-16'd16503;
      39485:data<=-16'd15605;
      39486:data<=-16'd15133;
      39487:data<=-16'd14721;
      39488:data<=-16'd14587;
      39489:data<=-16'd14499;
      39490:data<=-16'd14401;
      39491:data<=-16'd15221;
      39492:data<=-16'd15274;
      39493:data<=-16'd14023;
      39494:data<=-16'd14001;
      39495:data<=-16'd14237;
      39496:data<=-16'd13430;
      39497:data<=-16'd13132;
      39498:data<=-16'd12854;
      39499:data<=-16'd12084;
      39500:data<=-16'd11690;
      39501:data<=-16'd11485;
      39502:data<=-16'd11870;
      39503:data<=-16'd12969;
      39504:data<=-16'd13256;
      39505:data<=-16'd12273;
      39506:data<=-16'd11321;
      39507:data<=-16'd11063;
      39508:data<=-16'd10822;
      39509:data<=-16'd10492;
      39510:data<=-16'd10016;
      39511:data<=-16'd9048;
      39512:data<=-16'd8713;
      39513:data<=-16'd8859;
      39514:data<=-16'd8281;
      39515:data<=-16'd8361;
      39516:data<=-16'd9329;
      39517:data<=-16'd9182;
      39518:data<=-16'd8238;
      39519:data<=-16'd8022;
      39520:data<=-16'd7940;
      39521:data<=-16'd7239;
      39522:data<=-16'd7204;
      39523:data<=-16'd7206;
      39524:data<=-16'd6255;
      39525:data<=-16'd6469;
      39526:data<=-16'd6358;
      39527:data<=-16'd6156;
      39528:data<=-16'd8625;
      39529:data<=-16'd4511;
      39530:data<=16'd6839;
      39531:data<=16'd9324;
      39532:data<=16'd6053;
      39533:data<=16'd7359;
      39534:data<=16'd7269;
      39535:data<=16'd5959;
      39536:data<=16'd6860;
      39537:data<=16'd6346;
      39538:data<=16'd6106;
      39539:data<=16'd6633;
      39540:data<=16'd5403;
      39541:data<=16'd4217;
      39542:data<=16'd3471;
      39543:data<=16'd3207;
      39544:data<=16'd3600;
      39545:data<=16'd3206;
      39546:data<=16'd2974;
      39547:data<=16'd3380;
      39548:data<=16'd3700;
      39549:data<=16'd3709;
      39550:data<=16'd3086;
      39551:data<=16'd3021;
      39552:data<=16'd2907;
      39553:data<=16'd1891;
      39554:data<=16'd1768;
      39555:data<=16'd1556;
      39556:data<=16'd672;
      39557:data<=16'd587;
      39558:data<=16'd693;
      39559:data<=16'd951;
      39560:data<=16'd1005;
      39561:data<=16'd666;
      39562:data<=16'd735;
      39563:data<=16'd297;
      39564:data<=16'd250;
      39565:data<=-16'd5;
      39566:data<=-16'd2171;
      39567:data<=-16'd2622;
      39568:data<=-16'd1897;
      39569:data<=-16'd2491;
      39570:data<=-16'd2144;
      39571:data<=-16'd2162;
      39572:data<=-16'd2261;
      39573:data<=-16'd1339;
      39574:data<=-16'd1797;
      39575:data<=-16'd1055;
      39576:data<=-16'd541;
      39577:data<=-16'd1894;
      39578:data<=-16'd588;
      39579:data<=-16'd5147;
      39580:data<=-16'd16801;
      39581:data<=-16'd19182;
      39582:data<=-16'd15766;
      39583:data<=-16'd16146;
      39584:data<=-16'd15361;
      39585:data<=-16'd14320;
      39586:data<=-16'd14396;
      39587:data<=-16'd13244;
      39588:data<=-16'd12983;
      39589:data<=-16'd12668;
      39590:data<=-16'd12307;
      39591:data<=-16'd13220;
      39592:data<=-16'd12680;
      39593:data<=-16'd11872;
      39594:data<=-16'd11899;
      39595:data<=-16'd10818;
      39596:data<=-16'd9929;
      39597:data<=-16'd9706;
      39598:data<=-16'd9538;
      39599:data<=-16'd9527;
      39600:data<=-16'd8733;
      39601:data<=-16'd7558;
      39602:data<=-16'd7077;
      39603:data<=-16'd7943;
      39604:data<=-16'd9238;
      39605:data<=-16'd8883;
      39606:data<=-16'd7912;
      39607:data<=-16'd7121;
      39608:data<=-16'd6270;
      39609:data<=-16'd6213;
      39610:data<=-16'd5545;
      39611:data<=-16'd4871;
      39612:data<=-16'd5143;
      39613:data<=-16'd3657;
      39614:data<=-16'd2575;
      39615:data<=-16'd3789;
      39616:data<=-16'd4375;
      39617:data<=-16'd4664;
      39618:data<=-16'd4414;
      39619:data<=-16'd3576;
      39620:data<=-16'd3723;
      39621:data<=-16'd2955;
      39622:data<=-16'd2596;
      39623:data<=-16'd3224;
      39624:data<=-16'd2167;
      39625:data<=-16'd2375;
      39626:data<=-16'd2272;
      39627:data<=-16'd740;
      39628:data<=-16'd3239;
      39629:data<=-16'd889;
      39630:data<=16'd10202;
      39631:data<=16'd14064;
      39632:data<=16'd11323;
      39633:data<=16'd11996;
      39634:data<=16'd11905;
      39635:data<=16'd10753;
      39636:data<=16'd11209;
      39637:data<=16'd10749;
      39638:data<=16'd10507;
      39639:data<=16'd10819;
      39640:data<=16'd10040;
      39641:data<=16'd8942;
      39642:data<=16'd7787;
      39643:data<=16'd7485;
      39644:data<=16'd7975;
      39645:data<=16'd7580;
      39646:data<=16'd7150;
      39647:data<=16'd7144;
      39648:data<=16'd7188;
      39649:data<=16'd7500;
      39650:data<=16'd7034;
      39651:data<=16'd6351;
      39652:data<=16'd6648;
      39653:data<=16'd6388;
      39654:data<=16'd5225;
      39655:data<=16'd4731;
      39656:data<=16'd4684;
      39657:data<=16'd4155;
      39658:data<=16'd3882;
      39659:data<=16'd4109;
      39660:data<=16'd3962;
      39661:data<=16'd4099;
      39662:data<=16'd4159;
      39663:data<=16'd3231;
      39664:data<=16'd3287;
      39665:data<=16'd3742;
      39666:data<=16'd3127;
      39667:data<=16'd3269;
      39668:data<=16'd3171;
      39669:data<=16'd2796;
      39670:data<=16'd3874;
      39671:data<=16'd3607;
      39672:data<=16'd2958;
      39673:data<=16'd3923;
      39674:data<=16'd3691;
      39675:data<=16'd3688;
      39676:data<=16'd3589;
      39677:data<=16'd2604;
      39678:data<=16'd5037;
      39679:data<=16'd3401;
      39680:data<=-16'd6646;
      39681:data<=-16'd10845;
      39682:data<=-16'd8296;
      39683:data<=-16'd8549;
      39684:data<=-16'd8492;
      39685:data<=-16'd7413;
      39686:data<=-16'd7843;
      39687:data<=-16'd7336;
      39688:data<=-16'd6790;
      39689:data<=-16'd6801;
      39690:data<=-16'd5723;
      39691:data<=-16'd4114;
      39692:data<=-16'd2746;
      39693:data<=-16'd2783;
      39694:data<=-16'd3307;
      39695:data<=-16'd2726;
      39696:data<=-16'd2525;
      39697:data<=-16'd2205;
      39698:data<=-16'd1706;
      39699:data<=-16'd2478;
      39700:data<=-16'd2235;
      39701:data<=-16'd1202;
      39702:data<=-16'd1345;
      39703:data<=-16'd631;
      39704:data<=16'd572;
      39705:data<=16'd513;
      39706:data<=16'd529;
      39707:data<=16'd1001;
      39708:data<=16'd1037;
      39709:data<=16'd876;
      39710:data<=16'd1262;
      39711:data<=16'd1609;
      39712:data<=16'd1427;
      39713:data<=16'd1767;
      39714:data<=16'd1961;
      39715:data<=16'd2035;
      39716:data<=16'd3579;
      39717:data<=16'd4679;
      39718:data<=16'd4545;
      39719:data<=16'd4367;
      39720:data<=16'd3691;
      39721:data<=16'd3896;
      39722:data<=16'd4447;
      39723:data<=16'd3717;
      39724:data<=16'd3547;
      39725:data<=16'd3353;
      39726:data<=16'd3665;
      39727:data<=16'd4725;
      39728:data<=16'd3445;
      39729:data<=16'd6910;
      39730:data<=16'd17373;
      39731:data<=16'd21171;
      39732:data<=16'd18597;
      39733:data<=16'd18578;
      39734:data<=16'd18413;
      39735:data<=16'd17531;
      39736:data<=16'd16979;
      39737:data<=16'd15435;
      39738:data<=16'd15326;
      39739:data<=16'd15708;
      39740:data<=16'd15077;
      39741:data<=16'd15315;
      39742:data<=16'd15405;
      39743:data<=16'd15124;
      39744:data<=16'd14806;
      39745:data<=16'd13826;
      39746:data<=16'd13596;
      39747:data<=16'd13382;
      39748:data<=16'd12590;
      39749:data<=16'd12413;
      39750:data<=16'd11753;
      39751:data<=16'd10881;
      39752:data<=16'd10399;
      39753:data<=16'd10219;
      39754:data<=16'd11599;
      39755:data<=16'd12323;
      39756:data<=16'd11021;
      39757:data<=16'd10210;
      39758:data<=16'd9558;
      39759:data<=16'd8825;
      39760:data<=16'd8821;
      39761:data<=16'd8393;
      39762:data<=16'd7541;
      39763:data<=16'd6742;
      39764:data<=16'd6425;
      39765:data<=16'd6821;
      39766:data<=16'd7084;
      39767:data<=16'd7498;
      39768:data<=16'd7474;
      39769:data<=16'd6960;
      39770:data<=16'd7232;
      39771:data<=16'd6464;
      39772:data<=16'd5553;
      39773:data<=16'd6238;
      39774:data<=16'd5673;
      39775:data<=16'd5075;
      39776:data<=16'd4881;
      39777:data<=16'd3491;
      39778:data<=16'd4916;
      39779:data<=16'd4272;
      39780:data<=-16'd4639;
      39781:data<=-16'd10909;
      39782:data<=-16'd9931;
      39783:data<=-16'd9406;
      39784:data<=-16'd9644;
      39785:data<=-16'd9186;
      39786:data<=-16'd8994;
      39787:data<=-16'd8396;
      39788:data<=-16'd8238;
      39789:data<=-16'd8533;
      39790:data<=-16'd8272;
      39791:data<=-16'd7524;
      39792:data<=-16'd6344;
      39793:data<=-16'd5850;
      39794:data<=-16'd5888;
      39795:data<=-16'd5474;
      39796:data<=-16'd5591;
      39797:data<=-16'd5727;
      39798:data<=-16'd5325;
      39799:data<=-16'd5442;
      39800:data<=-16'd5506;
      39801:data<=-16'd5184;
      39802:data<=-16'd4801;
      39803:data<=-16'd4173;
      39804:data<=-16'd3920;
      39805:data<=-16'd3733;
      39806:data<=-16'd3124;
      39807:data<=-16'd2787;
      39808:data<=-16'd2625;
      39809:data<=-16'd2648;
      39810:data<=-16'd2826;
      39811:data<=-16'd2598;
      39812:data<=-16'd2529;
      39813:data<=-16'd2540;
      39814:data<=-16'd2346;
      39815:data<=-16'd2528;
      39816:data<=-16'd1924;
      39817:data<=-16'd300;
      39818:data<=16'd362;
      39819:data<=16'd150;
      39820:data<=-16'd36;
      39821:data<=-16'd326;
      39822:data<=-16'd622;
      39823:data<=-16'd801;
      39824:data<=-16'd564;
      39825:data<=-16'd415;
      39826:data<=-16'd769;
      39827:data<=-16'd876;
      39828:data<=-16'd1456;
      39829:data<=16'd247;
      39830:data<=16'd8621;
      39831:data<=16'd16372;
      39832:data<=16'd16304;
      39833:data<=16'd14527;
      39834:data<=16'd14242;
      39835:data<=16'd13283;
      39836:data<=16'd12883;
      39837:data<=16'd12380;
      39838:data<=16'd11577;
      39839:data<=16'd11371;
      39840:data<=16'd9906;
      39841:data<=16'd9377;
      39842:data<=16'd11082;
      39843:data<=16'd10865;
      39844:data<=16'd9382;
      39845:data<=16'd8916;
      39846:data<=16'd8479;
      39847:data<=16'd8238;
      39848:data<=16'd8006;
      39849:data<=16'd7732;
      39850:data<=16'd7673;
      39851:data<=16'd6696;
      39852:data<=16'd5659;
      39853:data<=16'd5780;
      39854:data<=16'd6619;
      39855:data<=16'd7415;
      39856:data<=16'd6959;
      39857:data<=16'd6064;
      39858:data<=16'd5542;
      39859:data<=16'd4795;
      39860:data<=16'd4874;
      39861:data<=16'd5056;
      39862:data<=16'd4258;
      39863:data<=16'd3647;
      39864:data<=16'd2690;
      39865:data<=16'd2032;
      39866:data<=16'd2258;
      39867:data<=16'd1603;
      39868:data<=16'd1072;
      39869:data<=16'd886;
      39870:data<=16'd408;
      39871:data<=16'd625;
      39872:data<=16'd77;
      39873:data<=-16'd425;
      39874:data<=16'd38;
      39875:data<=-16'd704;
      39876:data<=-16'd837;
      39877:data<=-16'd920;
      39878:data<=-16'd1832;
      39879:data<=-16'd1642;
      39880:data<=-16'd7650;
      39881:data<=-16'd18412;
      39882:data<=-16'd20321;
      39883:data<=-16'd17741;
      39884:data<=-16'd18207;
      39885:data<=-16'd17326;
      39886:data<=-16'd16392;
      39887:data<=-16'd16568;
      39888:data<=-16'd15876;
      39889:data<=-16'd15740;
      39890:data<=-16'd15089;
      39891:data<=-16'd14759;
      39892:data<=-16'd16190;
      39893:data<=-16'd16254;
      39894:data<=-16'd15329;
      39895:data<=-16'd14882;
      39896:data<=-16'd14345;
      39897:data<=-16'd14242;
      39898:data<=-16'd13888;
      39899:data<=-16'd13488;
      39900:data<=-16'd13530;
      39901:data<=-16'd13180;
      39902:data<=-16'd13009;
      39903:data<=-16'd12801;
      39904:data<=-16'd12989;
      39905:data<=-16'd13954;
      39906:data<=-16'd13590;
      39907:data<=-16'd12869;
      39908:data<=-16'd12458;
      39909:data<=-16'd11326;
      39910:data<=-16'd11189;
      39911:data<=-16'd10948;
      39912:data<=-16'd10028;
      39913:data<=-16'd10191;
      39914:data<=-16'd9318;
      39915:data<=-16'd8422;
      39916:data<=-16'd9570;
      39917:data<=-16'd10138;
      39918:data<=-16'd9987;
      39919:data<=-16'd9542;
      39920:data<=-16'd9034;
      39921:data<=-16'd9218;
      39922:data<=-16'd8296;
      39923:data<=-16'd7817;
      39924:data<=-16'd8137;
      39925:data<=-16'd7213;
      39926:data<=-16'd7653;
      39927:data<=-16'd7122;
      39928:data<=-16'd5981;
      39929:data<=-16'd9106;
      39930:data<=-16'd5447;
      39931:data<=16'd6590;
      39932:data<=16'd9721;
      39933:data<=16'd6830;
      39934:data<=16'd7514;
      39935:data<=16'd7072;
      39936:data<=16'd6011;
      39937:data<=16'd6191;
      39938:data<=16'd5554;
      39939:data<=16'd5747;
      39940:data<=16'd5958;
      39941:data<=16'd4874;
      39942:data<=16'd3791;
      39943:data<=16'd2711;
      39944:data<=16'd2338;
      39945:data<=16'd2499;
      39946:data<=16'd2499;
      39947:data<=16'd2789;
      39948:data<=16'd2567;
      39949:data<=16'd2382;
      39950:data<=16'd2833;
      39951:data<=16'd2881;
      39952:data<=16'd2893;
      39953:data<=16'd2504;
      39954:data<=16'd1575;
      39955:data<=16'd1011;
      39956:data<=16'd335;
      39957:data<=16'd135;
      39958:data<=16'd384;
      39959:data<=16'd258;
      39960:data<=16'd372;
      39961:data<=16'd26;
      39962:data<=16'd45;
      39963:data<=16'd832;
      39964:data<=16'd100;
      39965:data<=-16'd124;
      39966:data<=16'd89;
      39967:data<=-16'd1967;
      39968:data<=-16'd2940;
      39969:data<=-16'd2685;
      39970:data<=-16'd2993;
      39971:data<=-16'd2127;
      39972:data<=-16'd2087;
      39973:data<=-16'd2399;
      39974:data<=-16'd1650;
      39975:data<=-16'd2123;
      39976:data<=-16'd1497;
      39977:data<=-16'd978;
      39978:data<=-16'd1871;
      39979:data<=-16'd446;
      39980:data<=-16'd5292;
      39981:data<=-16'd17047;
      39982:data<=-16'd19699;
      39983:data<=-16'd16860;
      39984:data<=-16'd17511;
      39985:data<=-16'd16290;
      39986:data<=-16'd14687;
      39987:data<=-16'd14719;
      39988:data<=-16'd13509;
      39989:data<=-16'd13097;
      39990:data<=-16'd12715;
      39991:data<=-16'd11978;
      39992:data<=-16'd12866;
      39993:data<=-16'd12786;
      39994:data<=-16'd11806;
      39995:data<=-16'd11482;
      39996:data<=-16'd10804;
      39997:data<=-16'd10454;
      39998:data<=-16'd10088;
      39999:data<=-16'd9435;
      40000:data<=-16'd9191;
      40001:data<=-16'd8490;
      40002:data<=-16'd7885;
      40003:data<=-16'd7661;
      40004:data<=-16'd7679;
      40005:data<=-16'd8483;
      40006:data<=-16'd8531;
      40007:data<=-16'd8034;
      40008:data<=-16'd7893;
      40009:data<=-16'd7090;
      40010:data<=-16'd6441;
      40011:data<=-16'd5820;
      40012:data<=-16'd5313;
      40013:data<=-16'd5656;
      40014:data<=-16'd4440;
      40015:data<=-16'd3140;
      40016:data<=-16'd4041;
      40017:data<=-16'd4429;
      40018:data<=-16'd4269;
      40019:data<=-16'd3985;
      40020:data<=-16'd3594;
      40021:data<=-16'd4138;
      40022:data<=-16'd3365;
      40023:data<=-16'd2604;
      40024:data<=-16'd2960;
      40025:data<=-16'd1594;
      40026:data<=-16'd1730;
      40027:data<=-16'd2040;
      40028:data<=-16'd176;
      40029:data<=-16'd2067;
      40030:data<=16'd24;
      40031:data<=16'd10715;
      40032:data<=16'd14415;
      40033:data<=16'd11858;
      40034:data<=16'd12774;
      40035:data<=16'd12360;
      40036:data<=16'd11129;
      40037:data<=16'd11543;
      40038:data<=16'd10571;
      40039:data<=16'd10678;
      40040:data<=16'd11596;
      40041:data<=16'd10396;
      40042:data<=16'd9116;
      40043:data<=16'd8479;
      40044:data<=16'd8117;
      40045:data<=16'd7849;
      40046:data<=16'd7288;
      40047:data<=16'd7412;
      40048:data<=16'd7432;
      40049:data<=16'd7040;
      40050:data<=16'd7213;
      40051:data<=16'd7040;
      40052:data<=16'd7081;
      40053:data<=16'd7668;
      40054:data<=16'd6986;
      40055:data<=16'd5573;
      40056:data<=16'd4940;
      40057:data<=16'd5013;
      40058:data<=16'd4936;
      40059:data<=16'd4617;
      40060:data<=16'd4725;
      40061:data<=16'd4687;
      40062:data<=16'd4790;
      40063:data<=16'd5071;
      40064:data<=16'd3941;
      40065:data<=16'd3356;
      40066:data<=16'd4325;
      40067:data<=16'd4341;
      40068:data<=16'd4006;
      40069:data<=16'd3680;
      40070:data<=16'd3353;
      40071:data<=16'd4250;
      40072:data<=16'd4290;
      40073:data<=16'd3744;
      40074:data<=16'd4017;
      40075:data<=16'd3321;
      40076:data<=16'd3506;
      40077:data<=16'd4002;
      40078:data<=16'd3195;
      40079:data<=16'd4977;
      40080:data<=16'd3374;
      40081:data<=-16'd6024;
      40082:data<=-16'd10660;
      40083:data<=-16'd8768;
      40084:data<=-16'd8978;
      40085:data<=-16'd8687;
      40086:data<=-16'd7089;
      40087:data<=-16'd7333;
      40088:data<=-16'd7254;
      40089:data<=-16'd6771;
      40090:data<=-16'd6554;
      40091:data<=-16'd5424;
      40092:data<=-16'd4264;
      40093:data<=-16'd3482;
      40094:data<=-16'd2922;
      40095:data<=-16'd2347;
      40096:data<=-16'd1421;
      40097:data<=-16'd1438;
      40098:data<=-16'd1744;
      40099:data<=-16'd1219;
      40100:data<=-16'd1372;
      40101:data<=-16'd1565;
      40102:data<=-16'd1024;
      40103:data<=-16'd1080;
      40104:data<=-16'd623;
      40105:data<=16'd899;
      40106:data<=16'd1491;
      40107:data<=16'd1327;
      40108:data<=16'd1538;
      40109:data<=16'd1663;
      40110:data<=16'd1633;
      40111:data<=16'd1836;
      40112:data<=16'd1841;
      40113:data<=16'd1839;
      40114:data<=16'd2396;
      40115:data<=16'd2599;
      40116:data<=16'd2599;
      40117:data<=16'd3500;
      40118:data<=16'd4247;
      40119:data<=16'd4608;
      40120:data<=16'd5093;
      40121:data<=16'd4748;
      40122:data<=16'd4237;
      40123:data<=16'd4175;
      40124:data<=16'd4205;
      40125:data<=16'd4772;
      40126:data<=16'd4531;
      40127:data<=16'd3973;
      40128:data<=16'd4414;
      40129:data<=16'd3950;
      40130:data<=16'd7098;
      40131:data<=16'd16524;
      40132:data<=16'd21596;
      40133:data<=16'd20046;
      40134:data<=16'd19541;
      40135:data<=16'd19032;
      40136:data<=16'd17611;
      40137:data<=16'd17475;
      40138:data<=16'd16810;
      40139:data<=16'd16099;
      40140:data<=16'd15935;
      40141:data<=16'd15041;
      40142:data<=16'd15060;
      40143:data<=16'd15797;
      40144:data<=16'd15459;
      40145:data<=16'd14607;
      40146:data<=16'd13641;
      40147:data<=16'd13071;
      40148:data<=16'd12878;
      40149:data<=16'd12339;
      40150:data<=16'd11997;
      40151:data<=16'd11668;
      40152:data<=16'd10907;
      40153:data<=16'd10263;
      40154:data<=16'd10185;
      40155:data<=16'd10863;
      40156:data<=16'd11144;
      40157:data<=16'd10687;
      40158:data<=16'd10466;
      40159:data<=16'd9615;
      40160:data<=16'd8549;
      40161:data<=16'd8475;
      40162:data<=16'd8243;
      40163:data<=16'd7806;
      40164:data<=16'd7344;
      40165:data<=16'd6429;
      40166:data<=16'd6152;
      40167:data<=16'd6813;
      40168:data<=16'd7785;
      40169:data<=16'd7843;
      40170:data<=16'd6775;
      40171:data<=16'd6617;
      40172:data<=16'd6434;
      40173:data<=16'd5677;
      40174:data<=16'd5853;
      40175:data<=16'd4919;
      40176:data<=16'd4303;
      40177:data<=16'd5268;
      40178:data<=16'd3727;
      40179:data<=16'd3497;
      40180:data<=16'd4502;
      40181:data<=-16'd2341;
      40182:data<=-16'd10113;
      40183:data<=-16'd10270;
      40184:data<=-16'd9858;
      40185:data<=-16'd10442;
      40186:data<=-16'd9482;
      40187:data<=-16'd9185;
      40188:data<=-16'd8846;
      40189:data<=-16'd8607;
      40190:data<=-16'd9271;
      40191:data<=-16'd8813;
      40192:data<=-16'd7450;
      40193:data<=-16'd6068;
      40194:data<=-16'd5118;
      40195:data<=-16'd5131;
      40196:data<=-16'd4972;
      40197:data<=-16'd4825;
      40198:data<=-16'd5166;
      40199:data<=-16'd5112;
      40200:data<=-16'd4842;
      40201:data<=-16'd4611;
      40202:data<=-16'd4936;
      40203:data<=-16'd5598;
      40204:data<=-16'd4814;
      40205:data<=-16'd3290;
      40206:data<=-16'd2585;
      40207:data<=-16'd2563;
      40208:data<=-16'd2787;
      40209:data<=-16'd2547;
      40210:data<=-16'd2432;
      40211:data<=-16'd2601;
      40212:data<=-16'd2220;
      40213:data<=-16'd2484;
      40214:data<=-16'd2779;
      40215:data<=-16'd2268;
      40216:data<=-16'd2667;
      40217:data<=-16'd2234;
      40218:data<=-16'd405;
      40219:data<=-16'd77;
      40220:data<=-16'd328;
      40221:data<=-16'd499;
      40222:data<=-16'd920;
      40223:data<=-16'd676;
      40224:data<=-16'd1118;
      40225:data<=-16'd1245;
      40226:data<=-16'd578;
      40227:data<=-16'd1855;
      40228:data<=-16'd2050;
      40229:data<=-16'd879;
      40230:data<=-16'd829;
      40231:data<=16'd5048;
      40232:data<=16'd14486;
      40233:data<=16'd15975;
      40234:data<=16'd13926;
      40235:data<=16'd14320;
      40236:data<=16'd13311;
      40237:data<=16'd11978;
      40238:data<=16'd11782;
      40239:data<=16'd11116;
      40240:data<=16'd10545;
      40241:data<=16'd9535;
      40242:data<=16'd9203;
      40243:data<=16'd10381;
      40244:data<=16'd9932;
      40245:data<=16'd8790;
      40246:data<=16'd8813;
      40247:data<=16'd8370;
      40248:data<=16'd8143;
      40249:data<=16'd7978;
      40250:data<=16'd6772;
      40251:data<=16'd6238;
      40252:data<=16'd6112;
      40253:data<=16'd5442;
      40254:data<=16'd5348;
      40255:data<=16'd5780;
      40256:data<=16'd6029;
      40257:data<=16'd5809;
      40258:data<=16'd5377;
      40259:data<=16'd5178;
      40260:data<=16'd4808;
      40261:data<=16'd4269;
      40262:data<=16'd3562;
      40263:data<=16'd2840;
      40264:data<=16'd2504;
      40265:data<=16'd1754;
      40266:data<=16'd1181;
      40267:data<=16'd1143;
      40268:data<=16'd531;
      40269:data<=16'd629;
      40270:data<=16'd1033;
      40271:data<=16'd509;
      40272:data<=16'd514;
      40273:data<=16'd161;
      40274:data<=-16'd268;
      40275:data<=-16'd94;
      40276:data<=-16'd995;
      40277:data<=-16'd678;
      40278:data<=-16'd531;
      40279:data<=-16'd2083;
      40280:data<=-16'd1268;
      40281:data<=-16'd6055;
      40282:data<=-16'd17734;
      40283:data<=-16'd20298;
      40284:data<=-16'd17437;
      40285:data<=-16'd18624;
      40286:data<=-16'd17728;
      40287:data<=-16'd16457;
      40288:data<=-16'd16933;
      40289:data<=-16'd15854;
      40290:data<=-16'd15998;
      40291:data<=-16'd15796;
      40292:data<=-16'd14836;
      40293:data<=-16'd16251;
      40294:data<=-16'd16163;
      40295:data<=-16'd15109;
      40296:data<=-16'd15591;
      40297:data<=-16'd15000;
      40298:data<=-16'd14316;
      40299:data<=-16'd13925;
      40300:data<=-16'd13332;
      40301:data<=-16'd13295;
      40302:data<=-16'd12425;
      40303:data<=-16'd12198;
      40304:data<=-16'd12771;
      40305:data<=-16'd12399;
      40306:data<=-16'd12847;
      40307:data<=-16'd12757;
      40308:data<=-16'd11849;
      40309:data<=-16'd12152;
      40310:data<=-16'd11567;
      40311:data<=-16'd10866;
      40312:data<=-16'd10613;
      40313:data<=-16'd9373;
      40314:data<=-16'd9488;
      40315:data<=-16'd9652;
      40316:data<=-16'd8442;
      40317:data<=-16'd8508;
      40318:data<=-16'd9539;
      40319:data<=-16'd10716;
      40320:data<=-16'd10470;
      40321:data<=-16'd9015;
      40322:data<=-16'd9106;
      40323:data<=-16'd8654;
      40324:data<=-16'd8384;
      40325:data<=-16'd8983;
      40326:data<=-16'd7476;
      40327:data<=-16'd7908;
      40328:data<=-16'd8308;
      40329:data<=-16'd6182;
      40330:data<=-16'd8643;
      40331:data<=-16'd6294;
      40332:data<=16'd5268;
      40333:data<=16'd8479;
      40334:data<=16'd5974;
      40335:data<=16'd7544;
      40336:data<=16'd7119;
      40337:data<=16'd6213;
      40338:data<=16'd6701;
      40339:data<=16'd5583;
      40340:data<=16'd5770;
      40341:data<=16'd6256;
      40342:data<=16'd5054;
      40343:data<=16'd3689;
      40344:data<=16'd2353;
      40345:data<=16'd2244;
      40346:data<=16'd2431;
      40347:data<=16'd2197;
      40348:data<=16'd2698;
      40349:data<=16'd2211;
      40350:data<=16'd1744;
      40351:data<=16'd2112;
      40352:data<=16'd1554;
      40353:data<=16'd2036;
      40354:data<=16'd2634;
      40355:data<=16'd987;
      40356:data<=-16'd520;
      40357:data<=-16'd836;
      40358:data<=-16'd426;
      40359:data<=-16'd255;
      40360:data<=-16'd534;
      40361:data<=-16'd42;
      40362:data<=-16'd293;
      40363:data<=-16'd708;
      40364:data<=-16'd337;
      40365:data<=-16'd1111;
      40366:data<=-16'd895;
      40367:data<=-16'd693;
      40368:data<=-16'd2801;
      40369:data<=-16'd2861;
      40370:data<=-16'd2237;
      40371:data<=-16'd2869;
      40372:data<=-16'd2023;
      40373:data<=-16'd2027;
      40374:data<=-16'd1870;
      40375:data<=-16'd751;
      40376:data<=-16'd1915;
      40377:data<=-16'd1598;
      40378:data<=-16'd832;
      40379:data<=-16'd1721;
      40380:data<=-16'd325;
      40381:data<=-16'd5045;
      40382:data<=-16'd16342;
      40383:data<=-16'd19053;
      40384:data<=-16'd16797;
      40385:data<=-16'd17294;
      40386:data<=-16'd16193;
      40387:data<=-16'd15315;
      40388:data<=-16'd15206;
      40389:data<=-16'd13556;
      40390:data<=-16'd13253;
      40391:data<=-16'd13066;
      40392:data<=-16'd12149;
      40393:data<=-16'd12598;
      40394:data<=-16'd12333;
      40395:data<=-16'd11297;
      40396:data<=-16'd11169;
      40397:data<=-16'd10998;
      40398:data<=-16'd10358;
      40399:data<=-16'd9367;
      40400:data<=-16'd8831;
      40401:data<=-16'd8875;
      40402:data<=-16'd8436;
      40403:data<=-16'd7867;
      40404:data<=-16'd6954;
      40405:data<=-16'd6426;
      40406:data<=-16'd7556;
      40407:data<=-16'd7884;
      40408:data<=-16'd6889;
      40409:data<=-16'd6361;
      40410:data<=-16'd5755;
      40411:data<=-16'd5468;
      40412:data<=-16'd5380;
      40413:data<=-16'd4626;
      40414:data<=-16'd4249;
      40415:data<=-16'd3776;
      40416:data<=-16'd2971;
      40417:data<=-16'd2889;
      40418:data<=-16'd3398;
      40419:data<=-16'd4396;
      40420:data<=-16'd4360;
      40421:data<=-16'd3359;
      40422:data<=-16'd3435;
      40423:data<=-16'd2901;
      40424:data<=-16'd2334;
      40425:data<=-16'd2943;
      40426:data<=-16'd2100;
      40427:data<=-16'd1835;
      40428:data<=-16'd1882;
      40429:data<=-16'd408;
      40430:data<=-16'd2100;
      40431:data<=-16'd255;
      40432:data<=16'd10363;
      40433:data<=16'd15051;
      40434:data<=16'd12610;
      40435:data<=16'd13453;
      40436:data<=16'd13477;
      40437:data<=16'd11979;
      40438:data<=16'd12204;
      40439:data<=16'd11079;
      40440:data<=16'd10813;
      40441:data<=16'd12075;
      40442:data<=16'd11107;
      40443:data<=16'd9415;
      40444:data<=16'd8329;
      40445:data<=16'd7941;
      40446:data<=16'd8213;
      40447:data<=16'd7790;
      40448:data<=16'd7585;
      40449:data<=16'd7442;
      40450:data<=16'd7157;
      40451:data<=16'd7976;
      40452:data<=16'd7959;
      40453:data<=16'd7551;
      40454:data<=16'd8006;
      40455:data<=16'd6772;
      40456:data<=16'd5335;
      40457:data<=16'd5309;
      40458:data<=16'd4780;
      40459:data<=16'd4535;
      40460:data<=16'd4705;
      40461:data<=16'd4582;
      40462:data<=16'd4789;
      40463:data<=16'd4629;
      40464:data<=16'd4425;
      40465:data<=16'd4463;
      40466:data<=16'd4153;
      40467:data<=16'd4085;
      40468:data<=16'd4027;
      40469:data<=16'd4252;
      40470:data<=16'd4557;
      40471:data<=16'd3873;
      40472:data<=16'd3815;
      40473:data<=16'd4231;
      40474:data<=16'd4278;
      40475:data<=16'd4810;
      40476:data<=16'd4481;
      40477:data<=16'd4510;
      40478:data<=16'd4995;
      40479:data<=16'd3850;
      40480:data<=16'd5233;
      40481:data<=16'd4766;
      40482:data<=-16'd4408;
      40483:data<=-16'd10231;
      40484:data<=-16'd8305;
      40485:data<=-16'd8352;
      40486:data<=-16'd8545;
      40487:data<=-16'd7203;
      40488:data<=-16'd7429;
      40489:data<=-16'd6622;
      40490:data<=-16'd5685;
      40491:data<=-16'd5915;
      40492:data<=-16'd4942;
      40493:data<=-16'd3509;
      40494:data<=-16'd2032;
      40495:data<=-16'd1231;
      40496:data<=-16'd1885;
      40497:data<=-16'd1832;
      40498:data<=-16'd1474;
      40499:data<=-16'd1263;
      40500:data<=-16'd453;
      40501:data<=-16'd629;
      40502:data<=-16'd873;
      40503:data<=-16'd365;
      40504:data<=-16'd393;
      40505:data<=16'd384;
      40506:data<=16'd1727;
      40507:data<=16'd2290;
      40508:data<=16'd2805;
      40509:data<=16'd2740;
      40510:data<=16'd2355;
      40511:data<=16'd2739;
      40512:data<=16'd3283;
      40513:data<=16'd3548;
      40514:data<=16'd3236;
      40515:data<=16'd2989;
      40516:data<=16'd3330;
      40517:data<=16'd3530;
      40518:data<=16'd4434;
      40519:data<=16'd5470;
      40520:data<=16'd5189;
      40521:data<=16'd5009;
      40522:data<=16'd5001;
      40523:data<=16'd4927;
      40524:data<=16'd5007;
      40525:data<=16'd4106;
      40526:data<=16'd3882;
      40527:data<=16'd4540;
      40528:data<=16'd4347;
      40529:data<=16'd4837;
      40530:data<=16'd4937;
      40531:data<=16'd6811;
      40532:data<=16'd15575;
      40533:data<=16'd22692;
      40534:data<=16'd21678;
      40535:data<=16'd20169;
      40536:data<=16'd19898;
      40537:data<=16'd18788;
      40538:data<=16'd18515;
      40539:data<=16'd17737;
      40540:data<=16'd16957;
      40541:data<=16'd17152;
      40542:data<=16'd16228;
      40543:data<=16'd15899;
      40544:data<=16'd16807;
      40545:data<=16'd16460;
      40546:data<=16'd15738;
      40547:data<=16'd15320;
      40548:data<=16'd14639;
      40549:data<=16'd14160;
      40550:data<=16'd13506;
      40551:data<=16'd12895;
      40552:data<=16'd12825;
      40553:data<=16'd12524;
      40554:data<=16'd11897;
      40555:data<=16'd11841;
      40556:data<=16'd12612;
      40557:data<=16'd12687;
      40558:data<=16'd11491;
      40559:data<=16'd10801;
      40560:data<=16'd10433;
      40561:data<=16'd9508;
      40562:data<=16'd9039;
      40563:data<=16'd8801;
      40564:data<=16'd8479;
      40565:data<=16'd8372;
      40566:data<=16'd7652;
      40567:data<=16'd6884;
      40568:data<=16'd7491;
      40569:data<=16'd8895;
      40570:data<=16'd9215;
      40571:data<=16'd8308;
      40572:data<=16'd8178;
      40573:data<=16'd7961;
      40574:data<=16'd6796;
      40575:data<=16'd7000;
      40576:data<=16'd6784;
      40577:data<=16'd5470;
      40578:data<=16'd5758;
      40579:data<=16'd4784;
      40580:data<=16'd4529;
      40581:data<=16'd7133;
      40582:data<=16'd1676;
      40583:data<=-16'd9095;
      40584:data<=-16'd10674;
      40585:data<=-16'd8479;
      40586:data<=-16'd9409;
      40587:data<=-16'd9150;
      40588:data<=-16'd8883;
      40589:data<=-16'd8884;
      40590:data<=-16'd7797;
      40591:data<=-16'd8175;
      40592:data<=-16'd8182;
      40593:data<=-16'd6631;
      40594:data<=-16'd5861;
      40595:data<=-16'd5383;
      40596:data<=-16'd5197;
      40597:data<=-16'd5515;
      40598:data<=-16'd5580;
      40599:data<=-16'd5430;
      40600:data<=-16'd4878;
      40601:data<=-16'd5045;
      40602:data<=-16'd5653;
      40603:data<=-16'd5234;
      40604:data<=-16'd5219;
      40605:data<=-16'd5006;
      40606:data<=-16'd3735;
      40607:data<=-16'd3171;
      40608:data<=-16'd2831;
      40609:data<=-16'd2810;
      40610:data<=-16'd3106;
      40611:data<=-16'd2567;
      40612:data<=-16'd2837;
      40613:data<=-16'd3124;
      40614:data<=-16'd2422;
      40615:data<=-16'd2622;
      40616:data<=-16'd2488;
      40617:data<=-16'd2306;
      40618:data<=-16'd2525;
      40619:data<=-16'd980;
      40620:data<=-16'd312;
      40621:data<=-16'd1202;
      40622:data<=-16'd1363;
      40623:data<=-16'd1812;
      40624:data<=-16'd1554;
      40625:data<=-16'd1483;
      40626:data<=-16'd2375;
      40627:data<=-16'd1559;
      40628:data<=-16'd1673;
      40629:data<=-16'd1908;
      40630:data<=-16'd870;
      40631:data<=-16'd2309;
      40632:data<=16'd2469;
      40633:data<=16'd14001;
      40634:data<=16'd16032;
      40635:data<=16'd12812;
      40636:data<=16'd13479;
      40637:data<=16'd12577;
      40638:data<=16'd11752;
      40639:data<=16'd12113;
      40640:data<=16'd10624;
      40641:data<=16'd9943;
      40642:data<=16'd9329;
      40643:data<=16'd9056;
      40644:data<=16'd10460;
      40645:data<=16'd9800;
      40646:data<=16'd8583;
      40647:data<=16'd8728;
      40648:data<=16'd8208;
      40649:data<=16'd7937;
      40650:data<=16'd7301;
      40651:data<=16'd6237;
      40652:data<=16'd6317;
      40653:data<=16'd5832;
      40654:data<=16'd4893;
      40655:data<=16'd4780;
      40656:data<=16'd5413;
      40657:data<=16'd6191;
      40658:data<=16'd5403;
      40659:data<=16'd4673;
      40660:data<=16'd4828;
      40661:data<=16'd3885;
      40662:data<=16'd3551;
      40663:data<=16'd3284;
      40664:data<=16'd1953;
      40665:data<=16'd1950;
      40666:data<=16'd1635;
      40667:data<=16'd790;
      40668:data<=16'd1078;
      40669:data<=16'd588;
      40670:data<=16'd525;
      40671:data<=16'd893;
      40672:data<=16'd36;
      40673:data<=-16'd18;
      40674:data<=-16'd381;
      40675:data<=-16'd937;
      40676:data<=-16'd358;
      40677:data<=-16'd1281;
      40678:data<=-16'd1876;
      40679:data<=-16'd1941;
      40680:data<=-16'd2663;
      40681:data<=-16'd1521;
      40682:data<=-16'd6502;
      40683:data<=-16'd18146;
      40684:data<=-16'd21133;
      40685:data<=-16'd18404;
      40686:data<=-16'd18826;
      40687:data<=-16'd17987;
      40688:data<=-16'd17262;
      40689:data<=-16'd17960;
      40690:data<=-16'd17129;
      40691:data<=-16'd16707;
      40692:data<=-16'd16111;
      40693:data<=-16'd15916;
      40694:data<=-16'd17608;
      40695:data<=-16'd17406;
      40696:data<=-16'd16460;
      40697:data<=-16'd16841;
      40698:data<=-16'd16283;
      40699:data<=-16'd15793;
      40700:data<=-16'd15471;
      40701:data<=-16'd14524;
      40702:data<=-16'd14343;
      40703:data<=-16'd14340;
      40704:data<=-16'd14052;
      40705:data<=-16'd13697;
      40706:data<=-16'd13773;
      40707:data<=-16'd14613;
      40708:data<=-16'd14223;
      40709:data<=-16'd13458;
      40710:data<=-16'd13374;
      40711:data<=-16'd12205;
      40712:data<=-16'd11732;
      40713:data<=-16'd11914;
      40714:data<=-16'd11000;
      40715:data<=-16'd10922;
      40716:data<=-16'd10646;
      40717:data<=-16'd9875;
      40718:data<=-16'd10533;
      40719:data<=-16'd10992;
      40720:data<=-16'd11418;
      40721:data<=-16'd11703;
      40722:data<=-16'd10921;
      40723:data<=-16'd10883;
      40724:data<=-16'd10345;
      40725:data<=-16'd9644;
      40726:data<=-16'd9935;
      40727:data<=-16'd8916;
      40728:data<=-16'd8828;
      40729:data<=-16'd8408;
      40730:data<=-16'd6599;
      40731:data<=-16'd9306;
      40732:data<=-16'd7480;
      40733:data<=16'd3785;
      40734:data<=16'd7944;
      40735:data<=16'd5430;
      40736:data<=16'd6140;
      40737:data<=16'd5799;
      40738:data<=16'd5344;
      40739:data<=16'd6305;
      40740:data<=16'd5153;
      40741:data<=16'd4469;
      40742:data<=16'd4494;
      40743:data<=16'd3610;
      40744:data<=16'd2761;
      40745:data<=16'd1612;
      40746:data<=16'd1548;
      40747:data<=16'd2170;
      40748:data<=16'd2155;
      40749:data<=16'd2508;
      40750:data<=16'd1973;
      40751:data<=16'd1618;
      40752:data<=16'd2319;
      40753:data<=16'd1579;
      40754:data<=16'd1554;
      40755:data<=16'd2229;
      40756:data<=16'd796;
      40757:data<=-16'd276;
      40758:data<=-16'd420;
      40759:data<=-16'd651;
      40760:data<=-16'd503;
      40761:data<=-16'd781;
      40762:data<=-16'd834;
      40763:data<=-16'd814;
      40764:data<=-16'd1040;
      40765:data<=-16'd823;
      40766:data<=-16'd1366;
      40767:data<=-16'd1002;
      40768:data<=-16'd331;
      40769:data<=-16'd2594;
      40770:data<=-16'd3501;
      40771:data<=-16'd2319;
      40772:data<=-16'd2491;
      40773:data<=-16'd1926;
      40774:data<=-16'd1663;
      40775:data<=-16'd2077;
      40776:data<=-16'd1401;
      40777:data<=-16'd1989;
      40778:data<=-16'd2073;
      40779:data<=-16'd1671;
      40780:data<=-16'd2446;
      40781:data<=-16'd1037;
      40782:data<=-16'd4599;
      40783:data<=-16'd15620;
      40784:data<=-16'd19654;
      40785:data<=-16'd17183;
      40786:data<=-16'd17047;
      40787:data<=-16'd16418;
      40788:data<=-16'd15465;
      40789:data<=-16'd15406;
      40790:data<=-16'd14408;
      40791:data<=-16'd13574;
      40792:data<=-16'd12389;
      40793:data<=-16'd11935;
      40794:data<=-16'd13389;
      40795:data<=-16'd13355;
      40796:data<=-16'd12328;
      40797:data<=-16'd12069;
      40798:data<=-16'd11489;
      40799:data<=-16'd10959;
      40800:data<=-16'd10219;
      40801:data<=-16'd9400;
      40802:data<=-16'd9189;
      40803:data<=-16'd8781;
      40804:data<=-16'd8554;
      40805:data<=-16'd8069;
      40806:data<=-16'd7567;
      40807:data<=-16'd8664;
      40808:data<=-16'd8921;
      40809:data<=-16'd7746;
      40810:data<=-16'd7329;
      40811:data<=-16'd6545;
      40812:data<=-16'd5824;
      40813:data<=-16'd5635;
      40814:data<=-16'd4576;
      40815:data<=-16'd4203;
      40816:data<=-16'd4334;
      40817:data<=-16'd3717;
      40818:data<=-16'd3926;
      40819:data<=-16'd4564;
      40820:data<=-16'd4773;
      40821:data<=-16'd4748;
      40822:data<=-16'd4349;
      40823:data<=-16'd4279;
      40824:data<=-16'd3792;
      40825:data<=-16'd2892;
      40826:data<=-16'd2490;
      40827:data<=-16'd1532;
      40828:data<=-16'd1457;
      40829:data<=-16'd1462;
      40830:data<=16'd83;
      40831:data<=-16'd1538;
      40832:data<=-16'd1093;
      40833:data<=16'd8475;
      40834:data<=16'd14851;
      40835:data<=16'd13104;
      40836:data<=16'd12709;
      40837:data<=16'd12888;
      40838:data<=16'd12182;
      40839:data<=16'd12966;
      40840:data<=16'd12542;
      40841:data<=16'd11705;
      40842:data<=16'd11894;
      40843:data<=16'd11188;
      40844:data<=16'd10334;
      40845:data<=16'd9505;
      40846:data<=16'd8815;
      40847:data<=16'd9007;
      40848:data<=16'd8915;
      40849:data<=16'd9056;
      40850:data<=16'd9210;
      40851:data<=16'd8624;
      40852:data<=16'd8828;
      40853:data<=16'd8880;
      40854:data<=16'd8584;
      40855:data<=16'd9003;
      40856:data<=16'd8047;
      40857:data<=16'd6513;
      40858:data<=16'd6200;
      40859:data<=16'd5821;
      40860:data<=16'd5586;
      40861:data<=16'd5412;
      40862:data<=16'd5021;
      40863:data<=16'd5221;
      40864:data<=16'd5236;
      40865:data<=16'd5222;
      40866:data<=16'd5407;
      40867:data<=16'd5389;
      40868:data<=16'd5839;
      40869:data<=16'd5544;
      40870:data<=16'd4686;
      40871:data<=16'd4977;
      40872:data<=16'd5197;
      40873:data<=16'd5259;
      40874:data<=16'd5121;
      40875:data<=16'd4479;
      40876:data<=16'd4931;
      40877:data<=16'd4904;
      40878:data<=16'd4334;
      40879:data<=16'd4602;
      40880:data<=16'd3929;
      40881:data<=16'd5178;
      40882:data<=16'd5812;
      40883:data<=-16'd2144;
      40884:data<=-16'd9683;
      40885:data<=-16'd8954;
      40886:data<=-16'd8034;
      40887:data<=-16'd8243;
      40888:data<=-16'd7092;
      40889:data<=-16'd6860;
      40890:data<=-16'd6555;
      40891:data<=-16'd5944;
      40892:data<=-16'd5647;
      40893:data<=-16'd4629;
      40894:data<=-16'd3551;
      40895:data<=-16'd2531;
      40896:data<=-16'd1947;
      40897:data<=-16'd1770;
      40898:data<=-16'd1128;
      40899:data<=-16'd1697;
      40900:data<=-16'd2185;
      40901:data<=-16'd867;
      40902:data<=-16'd643;
      40903:data<=-16'd810;
      40904:data<=-16'd244;
      40905:data<=-16'd561;
      40906:data<=16'd229;
      40907:data<=16'd1997;
      40908:data<=16'd2232;
      40909:data<=16'd2209;
      40910:data<=16'd2799;
      40911:data<=16'd3269;
      40912:data<=16'd3178;
      40913:data<=16'd3011;
      40914:data<=16'd3515;
      40915:data<=16'd3513;
      40916:data<=16'd3421;
      40917:data<=16'd3656;
      40918:data<=16'd2969;
      40919:data<=16'd3735;
      40920:data<=16'd5459;
      40921:data<=16'd5140;
      40922:data<=16'd5250;
      40923:data<=16'd5315;
      40924:data<=16'd4287;
      40925:data<=16'd5012;
      40926:data<=16'd5231;
      40927:data<=16'd4683;
      40928:data<=16'd5700;
      40929:data<=16'd5651;
      40930:data<=16'd5551;
      40931:data<=16'd5782;
      40932:data<=16'd6191;
      40933:data<=16'd13524;
      40934:data<=16'd22604;
      40935:data<=16'd22753;
      40936:data<=16'd20316;
      40937:data<=16'd20251;
      40938:data<=16'd19270;
      40939:data<=16'd18694;
      40940:data<=16'd18618;
      40941:data<=16'd17984;
      40942:data<=16'd17258;
      40943:data<=16'd16017;
      40944:data<=16'd16216;
      40945:data<=16'd17382;
      40946:data<=16'd16644;
      40947:data<=16'd15666;
      40948:data<=16'd15314;
      40949:data<=16'd14596;
      40950:data<=16'd14008;
      40951:data<=16'd13271;
      40952:data<=16'd12751;
      40953:data<=16'd12777;
      40954:data<=16'd12260;
      40955:data<=16'd11468;
      40956:data<=16'd11500;
      40957:data<=16'd12490;
      40958:data<=16'd12878;
      40959:data<=16'd12031;
      40960:data<=16'd11427;
      40961:data<=16'd10348;
      40962:data<=16'd8962;
      40963:data<=16'd9157;
      40964:data<=16'd8940;
      40965:data<=16'd7953;
      40966:data<=16'd8025;
      40967:data<=16'd7570;
      40968:data<=16'd6764;
      40969:data<=16'd7345;
      40970:data<=16'd8596;
      40971:data<=16'd8962;
      40972:data<=16'd7797;
      40973:data<=16'd7450;
      40974:data<=16'd7667;
      40975:data<=16'd5959;
      40976:data<=16'd5389;
      40977:data<=16'd5547;
      40978:data<=16'd4255;
      40979:data<=16'd4807;
      40980:data<=16'd4231;
      40981:data<=16'd3137;
      40982:data<=16'd6590;
      40983:data<=16'd3087;
      40984:data<=-16'd8639;
      40985:data<=-16'd11379;
      40986:data<=-16'd8654;
      40987:data<=-16'd9876;
      40988:data<=-16'd9800;
      40989:data<=-16'd9383;
      40990:data<=-16'd10345;
      40991:data<=-16'd9292;
      40992:data<=-16'd8713;
      40993:data<=-16'd9000;
      40994:data<=-16'd7808;
      40995:data<=-16'd6517;
      40996:data<=-16'd5779;
      40997:data<=-16'd5559;
      40998:data<=-16'd5633;
      40999:data<=-16'd5724;
      41000:data<=-16'd6123;
      41001:data<=-16'd5799;
      41002:data<=-16'd5536;
      41003:data<=-16'd6003;
      41004:data<=-16'd5598;
      41005:data<=-16'd5530;
      41006:data<=-16'd5632;
      41007:data<=-16'd4071;
      41008:data<=-16'd3075;
      41009:data<=-16'd3263;
      41010:data<=-16'd3071;
      41011:data<=-16'd2736;
      41012:data<=-16'd2458;
      41013:data<=-16'd2623;
      41014:data<=-16'd2805;
      41015:data<=-16'd2725;
      41016:data<=-16'd3115;
      41017:data<=-16'd3078;
      41018:data<=-16'd3089;
      41019:data<=-16'd3078;
      41020:data<=-16'd1377;
      41021:data<=-16'd461;
      41022:data<=-16'd1042;
      41023:data<=-16'd1245;
      41024:data<=-16'd1542;
      41025:data<=-16'd946;
      41026:data<=-16'd741;
      41027:data<=-16'd1774;
      41028:data<=-16'd1152;
      41029:data<=-16'd1149;
      41030:data<=-16'd1441;
      41031:data<=-16'd657;
      41032:data<=-16'd1936;
      41033:data<=16'd2989;
      41034:data<=16'd14416;
      41035:data<=16'd16348;
      41036:data<=16'd13150;
      41037:data<=16'd14026;
      41038:data<=16'd13004;
      41039:data<=16'd11885;
      41040:data<=16'd12261;
      41041:data<=16'd10942;
      41042:data<=16'd10699;
      41043:data<=16'd10084;
      41044:data<=16'd9265;
      41045:data<=16'd10963;
      41046:data<=16'd10693;
      41047:data<=16'd9007;
      41048:data<=16'd8896;
      41049:data<=16'd8475;
      41050:data<=16'd8200;
      41051:data<=16'd7629;
      41052:data<=16'd6746;
      41053:data<=16'd6678;
      41054:data<=16'd5859;
      41055:data<=16'd5562;
      41056:data<=16'd5683;
      41057:data<=16'd4987;
      41058:data<=16'd5979;
      41059:data<=16'd6523;
      41060:data<=16'd5271;
      41061:data<=16'd5093;
      41062:data<=16'd4579;
      41063:data<=16'd3659;
      41064:data<=16'd3451;
      41065:data<=16'd2968;
      41066:data<=16'd2736;
      41067:data<=16'd2067;
      41068:data<=16'd1710;
      41069:data<=16'd2272;
      41070:data<=16'd1353;
      41071:data<=16'd755;
      41072:data<=16'd914;
      41073:data<=16'd385;
      41074:data<=16'd773;
      41075:data<=16'd58;
      41076:data<=-16'd1257;
      41077:data<=-16'd1199;
      41078:data<=-16'd2187;
      41079:data<=-16'd1911;
      41080:data<=-16'd1609;
      41081:data<=-16'd3162;
      41082:data<=-16'd1952;
      41083:data<=-16'd6329;
      41084:data<=-16'd18063;
      41085:data<=-16'd20985;
      41086:data<=-16'd18111;
      41087:data<=-16'd18516;
      41088:data<=-16'd17873;
      41089:data<=-16'd17581;
      41090:data<=-16'd17898;
      41091:data<=-16'd16774;
      41092:data<=-16'd16903;
      41093:data<=-16'd16154;
      41094:data<=-16'd15494;
      41095:data<=-16'd17224;
      41096:data<=-16'd17077;
      41097:data<=-16'd16251;
      41098:data<=-16'd16536;
      41099:data<=-16'd15843;
      41100:data<=-16'd15438;
      41101:data<=-16'd15151;
      41102:data<=-16'd14650;
      41103:data<=-16'd14516;
      41104:data<=-16'd13778;
      41105:data<=-16'd13486;
      41106:data<=-16'd13160;
      41107:data<=-16'd12848;
      41108:data<=-16'd14131;
      41109:data<=-16'd14095;
      41110:data<=-16'd13345;
      41111:data<=-16'd13840;
      41112:data<=-16'd12700;
      41113:data<=-16'd11693;
      41114:data<=-16'd12061;
      41115:data<=-16'd11462;
      41116:data<=-16'd11335;
      41117:data<=-16'd11124;
      41118:data<=-16'd10311;
      41119:data<=-16'd10904;
      41120:data<=-16'd11403;
      41121:data<=-16'd11312;
      41122:data<=-16'd11238;
      41123:data<=-16'd10916;
      41124:data<=-16'd10803;
      41125:data<=-16'd9662;
      41126:data<=-16'd8781;
      41127:data<=-16'd8843;
      41128:data<=-16'd7696;
      41129:data<=-16'd8108;
      41130:data<=-16'd8399;
      41131:data<=-16'd6728;
      41132:data<=-16'd8969;
      41133:data<=-16'd7248;
      41134:data<=16'd3644;
      41135:data<=16'd7879;
      41136:data<=16'd5045;
      41137:data<=16'd5803;
      41138:data<=16'd5803;
      41139:data<=16'd4575;
      41140:data<=16'd5429;
      41141:data<=16'd5092;
      41142:data<=16'd4488;
      41143:data<=16'd4551;
      41144:data<=16'd3457;
      41145:data<=16'd2331;
      41146:data<=16'd1838;
      41147:data<=16'd2023;
      41148:data<=16'd2159;
      41149:data<=16'd1579;
      41150:data<=16'd1639;
      41151:data<=16'd1707;
      41152:data<=16'd1616;
      41153:data<=16'd1870;
      41154:data<=16'd975;
      41155:data<=16'd861;
      41156:data<=16'd1847;
      41157:data<=16'd473;
      41158:data<=-16'd1077;
      41159:data<=-16'd820;
      41160:data<=-16'd1045;
      41161:data<=-16'd1445;
      41162:data<=-16'd1366;
      41163:data<=-16'd1416;
      41164:data<=-16'd1468;
      41165:data<=-16'd1334;
      41166:data<=-16'd1143;
      41167:data<=-16'd1368;
      41168:data<=-16'd1115;
      41169:data<=-16'd920;
      41170:data<=-16'd2808;
      41171:data<=-16'd4021;
      41172:data<=-16'd3472;
      41173:data<=-16'd3902;
      41174:data<=-16'd3747;
      41175:data<=-16'd2708;
      41176:data<=-16'd2828;
      41177:data<=-16'd3092;
      41178:data<=-16'd3071;
      41179:data<=-16'd2728;
      41180:data<=-16'd2908;
      41181:data<=-16'd3344;
      41182:data<=-16'd1909;
      41183:data<=-16'd5322;
      41184:data<=-16'd15749;
      41185:data<=-16'd20365;
      41186:data<=-16'd18077;
      41187:data<=-16'd17435;
      41188:data<=-16'd16935;
      41189:data<=-16'd15719;
      41190:data<=-16'd15294;
      41191:data<=-16'd14704;
      41192:data<=-16'd14419;
      41193:data<=-16'd13129;
      41194:data<=-16'd11693;
      41195:data<=-16'd12819;
      41196:data<=-16'd13591;
      41197:data<=-16'd12868;
      41198:data<=-16'd12446;
      41199:data<=-16'd11859;
      41200:data<=-16'd11333;
      41201:data<=-16'd10768;
      41202:data<=-16'd10160;
      41203:data<=-16'd10005;
      41204:data<=-16'd9389;
      41205:data<=-16'd8755;
      41206:data<=-16'd8049;
      41207:data<=-16'd7451;
      41208:data<=-16'd8675;
      41209:data<=-16'd9112;
      41210:data<=-16'd7799;
      41211:data<=-16'd7671;
      41212:data<=-16'd7274;
      41213:data<=-16'd6200;
      41214:data<=-16'd6072;
      41215:data<=-16'd5492;
      41216:data<=-16'd4804;
      41217:data<=-16'd4538;
      41218:data<=-16'd4030;
      41219:data<=-16'd4159;
      41220:data<=-16'd4569;
      41221:data<=-16'd4795;
      41222:data<=-16'd4667;
      41223:data<=-16'd3891;
      41224:data<=-16'd3738;
      41225:data<=-16'd3541;
      41226:data<=-16'd2948;
      41227:data<=-16'd2828;
      41228:data<=-16'd1838;
      41229:data<=-16'd1548;
      41230:data<=-16'd1798;
      41231:data<=-16'd267;
      41232:data<=-16'd1444;
      41233:data<=-16'd1577;
      41234:data<=16'd7175;
      41235:data<=16'd14134;
      41236:data<=16'd12778;
      41237:data<=16'd12131;
      41238:data<=16'd12665;
      41239:data<=16'd11512;
      41240:data<=16'd11397;
      41241:data<=16'd11699;
      41242:data<=16'd11295;
      41243:data<=16'd11053;
      41244:data<=16'd10831;
      41245:data<=16'd9837;
      41246:data<=16'd8308;
      41247:data<=16'd8493;
      41248:data<=16'd9274;
      41249:data<=16'd8243;
      41250:data<=16'd7853;
      41251:data<=16'd8185;
      41252:data<=16'd7702;
      41253:data<=16'd7932;
      41254:data<=16'd7968;
      41255:data<=16'd7685;
      41256:data<=16'd8109;
      41257:data<=16'd7227;
      41258:data<=16'd5953;
      41259:data<=16'd5788;
      41260:data<=16'd5501;
      41261:data<=16'd5538;
      41262:data<=16'd5498;
      41263:data<=16'd5180;
      41264:data<=16'd5392;
      41265:data<=16'd5072;
      41266:data<=16'd5281;
      41267:data<=16'd6005;
      41268:data<=16'd5294;
      41269:data<=16'd5313;
      41270:data<=16'd5868;
      41271:data<=16'd5184;
      41272:data<=16'd5201;
      41273:data<=16'd5433;
      41274:data<=16'd5395;
      41275:data<=16'd5753;
      41276:data<=16'd5315;
      41277:data<=16'd5162;
      41278:data<=16'd5228;
      41279:data<=16'd4857;
      41280:data<=16'd5204;
      41281:data<=16'd4584;
      41282:data<=16'd5321;
      41283:data<=16'd7212;
      41284:data<=16'd1143;
      41285:data<=-16'd7368;
      41286:data<=-16'd7509;
      41287:data<=-16'd6159;
      41288:data<=-16'd6792;
      41289:data<=-16'd5369;
      41290:data<=-16'd4602;
      41291:data<=-16'd4842;
      41292:data<=-16'd4176;
      41293:data<=-16'd3779;
      41294:data<=-16'd3203;
      41295:data<=-16'd1924;
      41296:data<=-16'd496;
      41297:data<=16'd303;
      41298:data<=16'd353;
      41299:data<=16'd587;
      41300:data<=16'd453;
      41301:data<=16'd694;
      41302:data<=16'd1626;
      41303:data<=16'd1122;
      41304:data<=16'd1063;
      41305:data<=16'd1871;
      41306:data<=16'd1384;
      41307:data<=16'd2352;
      41308:data<=16'd4225;
      41309:data<=16'd4314;
      41310:data<=16'd4552;
      41311:data<=16'd4443;
      41312:data<=16'd3967;
      41313:data<=16'd4570;
      41314:data<=16'd4710;
      41315:data<=16'd4905;
      41316:data<=16'd4804;
      41317:data<=16'd3938;
      41318:data<=16'd4707;
      41319:data<=16'd5043;
      41320:data<=16'd4949;
      41321:data<=16'd6743;
      41322:data<=16'd6910;
      41323:data<=16'd6256;
      41324:data<=16'd6667;
      41325:data<=16'd5953;
      41326:data<=16'd6325;
      41327:data<=16'd6810;
      41328:data<=16'd5897;
      41329:data<=16'd6672;
      41330:data<=16'd6437;
      41331:data<=16'd5826;
      41332:data<=16'd6825;
      41333:data<=16'd6167;
      41334:data<=16'd11236;
      41335:data<=16'd21631;
      41336:data<=16'd22856;
      41337:data<=16'd19782;
      41338:data<=16'd20525;
      41339:data<=16'd19690;
      41340:data<=16'd18630;
      41341:data<=16'd18318;
      41342:data<=16'd16915;
      41343:data<=16'd17149;
      41344:data<=16'd16882;
      41345:data<=16'd15800;
      41346:data<=16'd16504;
      41347:data<=16'd16277;
      41348:data<=16'd15552;
      41349:data<=16'd15412;
      41350:data<=16'd14387;
      41351:data<=16'd13893;
      41352:data<=16'd13667;
      41353:data<=16'd13141;
      41354:data<=16'd12863;
      41355:data<=16'd11972;
      41356:data<=16'd11558;
      41357:data<=16'd11644;
      41358:data<=16'd11708;
      41359:data<=16'd12325;
      41360:data<=16'd11614;
      41361:data<=16'd10760;
      41362:data<=16'd10944;
      41363:data<=16'd9696;
      41364:data<=16'd8751;
      41365:data<=16'd8563;
      41366:data<=16'd7967;
      41367:data<=16'd8636;
      41368:data<=16'd8160;
      41369:data<=16'd6654;
      41370:data<=16'd7492;
      41371:data<=16'd8282;
      41372:data<=16'd8122;
      41373:data<=16'd7931;
      41374:data<=16'd7688;
      41375:data<=16'd7867;
      41376:data<=16'd6649;
      41377:data<=16'd5782;
      41378:data<=16'd6100;
      41379:data<=16'd4667;
      41380:data<=16'd4675;
      41381:data<=16'd4687;
      41382:data<=16'd3462;
      41383:data<=16'd6437;
      41384:data<=16'd3422;
      41385:data<=-16'd8191;
      41386:data<=-16'd10645;
      41387:data<=-16'd7655;
      41388:data<=-16'd9159;
      41389:data<=-16'd8570;
      41390:data<=-16'd7535;
      41391:data<=-16'd8417;
      41392:data<=-16'd7668;
      41393:data<=-16'd7943;
      41394:data<=-16'd8437;
      41395:data<=-16'd7003;
      41396:data<=-16'd5915;
      41397:data<=-16'd5400;
      41398:data<=-16'd5548;
      41399:data<=-16'd5480;
      41400:data<=-16'd4690;
      41401:data<=-16'd4828;
      41402:data<=-16'd4925;
      41403:data<=-16'd5060;
      41404:data<=-16'd5429;
      41405:data<=-16'd4748;
      41406:data<=-16'd4843;
      41407:data<=-16'd4968;
      41408:data<=-16'd3435;
      41409:data<=-16'd2519;
      41410:data<=-16'd2384;
      41411:data<=-16'd2511;
      41412:data<=-16'd2861;
      41413:data<=-16'd2770;
      41414:data<=-16'd2928;
      41415:data<=-16'd2575;
      41416:data<=-16'd2196;
      41417:data<=-16'd2773;
      41418:data<=-16'd2432;
      41419:data<=-16'd2484;
      41420:data<=-16'd2698;
      41421:data<=-16'd1072;
      41422:data<=-16'd711;
      41423:data<=-16'd1107;
      41424:data<=-16'd892;
      41425:data<=-16'd1645;
      41426:data<=-16'd1242;
      41427:data<=-16'd1069;
      41428:data<=-16'd1765;
      41429:data<=-16'd479;
      41430:data<=-16'd840;
      41431:data<=-16'd1571;
      41432:data<=-16'd1034;
      41433:data<=-16'd2863;
      41434:data<=16'd2137;
      41435:data<=16'd13538;
      41436:data<=16'd15208;
      41437:data<=16'd12135;
      41438:data<=16'd12812;
      41439:data<=16'd11758;
      41440:data<=16'd10654;
      41441:data<=16'd10633;
      41442:data<=16'd9597;
      41443:data<=16'd10003;
      41444:data<=16'd9541;
      41445:data<=16'd7991;
      41446:data<=16'd8909;
      41447:data<=16'd9702;
      41448:data<=16'd9286;
      41449:data<=16'd8874;
      41450:data<=16'd7770;
      41451:data<=16'd6910;
      41452:data<=16'd6589;
      41453:data<=16'd6161;
      41454:data<=16'd5573;
      41455:data<=16'd4983;
      41456:data<=16'd4652;
      41457:data<=16'd3654;
      41458:data<=16'd3580;
      41459:data<=16'd5515;
      41460:data<=16'd5547;
      41461:data<=16'd4246;
      41462:data<=16'd4508;
      41463:data<=16'd4311;
      41464:data<=16'd3327;
      41465:data<=16'd2558;
      41466:data<=16'd2062;
      41467:data<=16'd2238;
      41468:data<=16'd1986;
      41469:data<=16'd1544;
      41470:data<=16'd1347;
      41471:data<=16'd773;
      41472:data<=16'd749;
      41473:data<=16'd331;
      41474:data<=-16'd214;
      41475:data<=16'd328;
      41476:data<=-16'd415;
      41477:data<=-16'd913;
      41478:data<=-16'd585;
      41479:data<=-16'd1994;
      41480:data<=-16'd1624;
      41481:data<=-16'd967;
      41482:data<=-16'd2250;
      41483:data<=-16'd1274;
      41484:data<=-16'd5761;
      41485:data<=-16'd17117;
      41486:data<=-16'd20224;
      41487:data<=-16'd17594;
      41488:data<=-16'd18117;
      41489:data<=-16'd17540;
      41490:data<=-16'd16392;
      41491:data<=-16'd16396;
      41492:data<=-16'd15825;
      41493:data<=-16'd16011;
      41494:data<=-16'd15716;
      41495:data<=-16'd15144;
      41496:data<=-16'd16110;
      41497:data<=-16'd16496;
      41498:data<=-16'd16409;
      41499:data<=-16'd16161;
      41500:data<=-16'd15032;
      41501:data<=-16'd14569;
      41502:data<=-16'd14339;
      41503:data<=-16'd13908;
      41504:data<=-16'd13606;
      41505:data<=-16'd12827;
      41506:data<=-16'd12468;
      41507:data<=-16'd12002;
      41508:data<=-16'd11884;
      41509:data<=-16'd13585;
      41510:data<=-16'd13946;
      41511:data<=-16'd12963;
      41512:data<=-16'd13176;
      41513:data<=-16'd12824;
      41514:data<=-16'd12020;
      41515:data<=-16'd11339;
      41516:data<=-16'd10548;
      41517:data<=-16'd10906;
      41518:data<=-16'd10681;
      41519:data<=-16'd9793;
      41520:data<=-16'd10257;
      41521:data<=-16'd10781;
      41522:data<=-16'd11300;
      41523:data<=-16'd11253;
      41524:data<=-16'd10208;
      41525:data<=-16'd10290;
      41526:data<=-16'd9879;
      41527:data<=-16'd9107;
      41528:data<=-16'd9508;
      41529:data<=-16'd8499;
      41530:data<=-16'd8022;
      41531:data<=-16'd8298;
      41532:data<=-16'd7371;
      41533:data<=-16'd9407;
      41534:data<=-16'd8070;
      41535:data<=16'd2099;
      41536:data<=16'd7403;
      41537:data<=16'd5192;
      41538:data<=16'd5077;
      41539:data<=16'd5292;
      41540:data<=16'd4414;
      41541:data<=16'd4337;
      41542:data<=16'd3929;
      41543:data<=16'd4175;
      41544:data<=16'd4375;
      41545:data<=16'd3353;
      41546:data<=16'd2396;
      41547:data<=16'd1410;
      41548:data<=16'd1259;
      41549:data<=16'd1560;
      41550:data<=16'd846;
      41551:data<=16'd829;
      41552:data<=16'd839;
      41553:data<=16'd214;
      41554:data<=16'd845;
      41555:data<=16'd834;
      41556:data<=-16'd146;
      41557:data<=16'd103;
      41558:data<=-16'd182;
      41559:data<=-16'd1495;
      41560:data<=-16'd1905;
      41561:data<=-16'd1501;
      41562:data<=-16'd1193;
      41563:data<=-16'd1386;
      41564:data<=-16'd1545;
      41565:data<=-16'd1621;
      41566:data<=-16'd1935;
      41567:data<=-16'd1689;
      41568:data<=-16'd1503;
      41569:data<=-16'd1756;
      41570:data<=-16'd1757;
      41571:data<=-16'd2672;
      41572:data<=-16'd3759;
      41573:data<=-16'd3539;
      41574:data<=-16'd3466;
      41575:data<=-16'd3615;
      41576:data<=-16'd3377;
      41577:data<=-16'd3098;
      41578:data<=-16'd2807;
      41579:data<=-16'd3257;
      41580:data<=-16'd3557;
      41581:data<=-16'd3193;
      41582:data<=-16'd2986;
      41583:data<=-16'd2046;
      41584:data<=-16'd4936;
      41585:data<=-16'd14336;
      41586:data<=-16'd19772;
      41587:data<=-16'd18063;
      41588:data<=-16'd17182;
      41589:data<=-16'd16971;
      41590:data<=-16'd15764;
      41591:data<=-16'd15490;
      41592:data<=-16'd14742;
      41593:data<=-16'd13728;
      41594:data<=-16'd13339;
      41595:data<=-16'd12609;
      41596:data<=-16'd12827;
      41597:data<=-16'd13700;
      41598:data<=-16'd13303;
      41599:data<=-16'd12419;
      41600:data<=-16'd11838;
      41601:data<=-16'd11382;
      41602:data<=-16'd10796;
      41603:data<=-16'd9906;
      41604:data<=-16'd9365;
      41605:data<=-16'd9209;
      41606:data<=-16'd8737;
      41607:data<=-16'd7817;
      41608:data<=-16'd7474;
      41609:data<=-16'd8490;
      41610:data<=-16'd9048;
      41611:data<=-16'd8358;
      41612:data<=-16'd7975;
      41613:data<=-16'd7600;
      41614:data<=-16'd7077;
      41615:data<=-16'd6742;
      41616:data<=-16'd5614;
      41617:data<=-16'd4810;
      41618:data<=-16'd5033;
      41619:data<=-16'd4534;
      41620:data<=-16'd3802;
      41621:data<=-16'd4225;
      41622:data<=-16'd5265;
      41623:data<=-16'd5523;
      41624:data<=-16'd4843;
      41625:data<=-16'd4643;
      41626:data<=-16'd4223;
      41627:data<=-16'd3192;
      41628:data<=-16'd3233;
      41629:data<=-16'd2951;
      41630:data<=-16'd2237;
      41631:data<=-16'd2476;
      41632:data<=-16'd1838;
      41633:data<=-16'd2297;
      41634:data<=-16'd2678;
      41635:data<=16'd4316;
      41636:data<=16'd12149;
      41637:data<=16'd12000;
      41638:data<=16'd10780;
      41639:data<=16'd11586;
      41640:data<=16'd10953;
      41641:data<=16'd10828;
      41642:data<=16'd11027;
      41643:data<=16'd10229;
      41644:data<=16'd10392;
      41645:data<=16'd10922;
      41646:data<=16'd10223;
      41647:data<=16'd8675;
      41648:data<=16'd7723;
      41649:data<=16'd7917;
      41650:data<=16'd7483;
      41651:data<=16'd6737;
      41652:data<=16'd6992;
      41653:data<=16'd6904;
      41654:data<=16'd6728;
      41655:data<=16'd6968;
      41656:data<=16'd6498;
      41657:data<=16'd6209;
      41658:data<=16'd6197;
      41659:data<=16'd5307;
      41660:data<=16'd4435;
      41661:data<=16'd4246;
      41662:data<=16'd4411;
      41663:data<=16'd4622;
      41664:data<=16'd4660;
      41665:data<=16'd4555;
      41666:data<=16'd4111;
      41667:data<=16'd3990;
      41668:data<=16'd4425;
      41669:data<=16'd4381;
      41670:data<=16'd4326;
      41671:data<=16'd4481;
      41672:data<=16'd4617;
      41673:data<=16'd5177;
      41674:data<=16'd4925;
      41675:data<=16'd4284;
      41676:data<=16'd4534;
      41677:data<=16'd4363;
      41678:data<=16'd4337;
      41679:data<=16'd4444;
      41680:data<=16'd3899;
      41681:data<=16'd4473;
      41682:data<=16'd4467;
      41683:data<=16'd4684;
      41684:data<=16'd7291;
      41685:data<=16'd3730;
      41686:data<=-16'd5206;
      41687:data<=-16'd6796;
      41688:data<=-16'd4538;
      41689:data<=-16'd5224;
      41690:data<=-16'd4904;
      41691:data<=-16'd4391;
      41692:data<=-16'd4822;
      41693:data<=-16'd3877;
      41694:data<=-16'd3366;
      41695:data<=-16'd3594;
      41696:data<=-16'd2667;
      41697:data<=-16'd966;
      41698:data<=-16'd21;
      41699:data<=-16'd459;
      41700:data<=-16'd112;
      41701:data<=16'd1045;
      41702:data<=16'd767;
      41703:data<=16'd655;
      41704:data<=16'd1154;
      41705:data<=16'd931;
      41706:data<=16'd1215;
      41707:data<=16'd1833;
      41708:data<=16'd2353;
      41709:data<=16'd3482;
      41710:data<=16'd4226;
      41711:data<=16'd4367;
      41712:data<=16'd4554;
      41713:data<=16'd4563;
      41714:data<=16'd4149;
      41715:data<=16'd3720;
      41716:data<=16'd4223;
      41717:data<=16'd4645;
      41718:data<=16'd4170;
      41719:data<=16'd4077;
      41720:data<=16'd4049;
      41721:data<=16'd4696;
      41722:data<=16'd6246;
      41723:data<=16'd6162;
      41724:data<=16'd5853;
      41725:data<=16'd6273;
      41726:data<=16'd5789;
      41727:data<=16'd5900;
      41728:data<=16'd5711;
      41729:data<=16'd5301;
      41730:data<=16'd6434;
      41731:data<=16'd5570;
      41732:data<=16'd4949;
      41733:data<=16'd6328;
      41734:data<=16'd5134;
      41735:data<=16'd9253;
      41736:data<=16'd19387;
      41737:data<=16'd20739;
      41738:data<=16'd17552;
      41739:data<=16'd18240;
      41740:data<=16'd17390;
      41741:data<=16'd16519;
      41742:data<=16'd16838;
      41743:data<=16'd15481;
      41744:data<=16'd15355;
      41745:data<=16'd15462;
      41746:data<=16'd14929;
      41747:data<=16'd15793;
      41748:data<=16'd15602;
      41749:data<=16'd14963;
      41750:data<=16'd14739;
      41751:data<=16'd13280;
      41752:data<=16'd12831;
      41753:data<=16'd12747;
      41754:data<=16'd11767;
      41755:data<=16'd11803;
      41756:data<=16'd11154;
      41757:data<=16'd9947;
      41758:data<=16'd10158;
      41759:data<=16'd10525;
      41760:data<=16'd10994;
      41761:data<=16'd10881;
      41762:data<=16'd9915;
      41763:data<=16'd9897;
      41764:data<=16'd9652;
      41765:data<=16'd8901;
      41766:data<=16'd8545;
      41767:data<=16'd7746;
      41768:data<=16'd7406;
      41769:data<=16'd7275;
      41770:data<=16'd6636;
      41771:data<=16'd7034;
      41772:data<=16'd8128;
      41773:data<=16'd8737;
      41774:data<=16'd8285;
      41775:data<=16'd7536;
      41776:data<=16'd7624;
      41777:data<=16'd6777;
      41778:data<=16'd5909;
      41779:data<=16'd5970;
      41780:data<=16'd4999;
      41781:data<=16'd5433;
      41782:data<=16'd5592;
      41783:data<=16'd4055;
      41784:data<=16'd6448;
      41785:data<=16'd4804;
      41786:data<=-16'd5095;
      41787:data<=-16'd8255;
      41788:data<=-16'd5905;
      41789:data<=-16'd6909;
      41790:data<=-16'd6583;
      41791:data<=-16'd6209;
      41792:data<=-16'd7028;
      41793:data<=-16'd5815;
      41794:data<=-16'd6006;
      41795:data<=-16'd6695;
      41796:data<=-16'd5630;
      41797:data<=-16'd4749;
      41798:data<=-16'd3336;
      41799:data<=-16'd3253;
      41800:data<=-16'd4350;
      41801:data<=-16'd3541;
      41802:data<=-16'd3430;
      41803:data<=-16'd3653;
      41804:data<=-16'd2654;
      41805:data<=-16'd3015;
      41806:data<=-16'd3307;
      41807:data<=-16'd2776;
      41808:data<=-16'd2849;
      41809:data<=-16'd2027;
      41810:data<=-16'd698;
      41811:data<=-16'd185;
      41812:data<=-16'd337;
      41813:data<=-16'd660;
      41814:data<=-16'd550;
      41815:data<=-16'd914;
      41816:data<=-16'd1183;
      41817:data<=-16'd560;
      41818:data<=-16'd699;
      41819:data<=-16'd1130;
      41820:data<=-16'd1181;
      41821:data<=-16'd782;
      41822:data<=16'd506;
      41823:data<=16'd638;
      41824:data<=-16'd18;
      41825:data<=16'd91;
      41826:data<=16'd130;
      41827:data<=16'd561;
      41828:data<=16'd193;
      41829:data<=-16'd394;
      41830:data<=16'd579;
      41831:data<=-16'd367;
      41832:data<=-16'd1010;
      41833:data<=16'd56;
      41834:data<=-16'd1494;
      41835:data<=16'd2455;
      41836:data<=16'd12474;
      41837:data<=16'd14563;
      41838:data<=16'd12430;
      41839:data<=16'd12786;
      41840:data<=16'd11479;
      41841:data<=16'd10975;
      41842:data<=16'd11168;
      41843:data<=16'd9494;
      41844:data<=16'd9292;
      41845:data<=16'd9230;
      41846:data<=16'd8740;
      41847:data<=16'd9661;
      41848:data<=16'd9433;
      41849:data<=16'd8721;
      41850:data<=16'd8702;
      41851:data<=16'd8100;
      41852:data<=16'd7776;
      41853:data<=16'd7089;
      41854:data<=16'd6067;
      41855:data<=16'd5879;
      41856:data<=16'd5324;
      41857:data<=16'd4701;
      41858:data<=16'd4126;
      41859:data<=16'd3539;
      41860:data<=16'd4419;
      41861:data<=16'd5001;
      41862:data<=16'd4378;
      41863:data<=16'd4222;
      41864:data<=16'd3817;
      41865:data<=16'd3233;
      41866:data<=16'd2951;
      41867:data<=16'd2194;
      41868:data<=16'd1656;
      41869:data<=16'd1600;
      41870:data<=16'd1466;
      41871:data<=16'd981;
      41872:data<=16'd376;
      41873:data<=16'd456;
      41874:data<=16'd332;
      41875:data<=-16'd167;
      41876:data<=-16'd287;
      41877:data<=-16'd1030;
      41878:data<=-16'd1497;
      41879:data<=-16'd1422;
      41880:data<=-16'd1855;
      41881:data<=-16'd1318;
      41882:data<=-16'd1563;
      41883:data<=-16'd2692;
      41884:data<=-16'd1838;
      41885:data<=-16'd5553;
      41886:data<=-16'd14832;
      41887:data<=-16'd18490;
      41888:data<=-16'd16917;
      41889:data<=-16'd16477;
      41890:data<=-16'd16157;
      41891:data<=-16'd16160;
      41892:data<=-16'd16222;
      41893:data<=-16'd15135;
      41894:data<=-16'd14786;
      41895:data<=-16'd14791;
      41896:data<=-16'd14875;
      41897:data<=-16'd16022;
      41898:data<=-16'd16290;
      41899:data<=-16'd15550;
      41900:data<=-16'd15362;
      41901:data<=-16'd15218;
      41902:data<=-16'd14800;
      41903:data<=-16'd14069;
      41904:data<=-16'd13195;
      41905:data<=-16'd12778;
      41906:data<=-16'd12660;
      41907:data<=-16'd12377;
      41908:data<=-16'd11579;
      41909:data<=-16'd11411;
      41910:data<=-16'd12515;
      41911:data<=-16'd12572;
      41912:data<=-16'd11655;
      41913:data<=-16'd11623;
      41914:data<=-16'd11549;
      41915:data<=-16'd11262;
      41916:data<=-16'd11042;
      41917:data<=-16'd10225;
      41918:data<=-16'd9838;
      41919:data<=-16'd10000;
      41920:data<=-16'd9682;
      41921:data<=-16'd9489;
      41922:data<=-16'd10079;
      41923:data<=-16'd10903;
      41924:data<=-16'd10658;
      41925:data<=-16'd9855;
      41926:data<=-16'd9799;
      41927:data<=-16'd9157;
      41928:data<=-16'd8251;
      41929:data<=-16'd8220;
      41930:data<=-16'd7785;
      41931:data<=-16'd7958;
      41932:data<=-16'd8193;
      41933:data<=-16'd7322;
      41934:data<=-16'd8821;
      41935:data<=-16'd8326;
      41936:data<=-16'd502;
      41937:data<=16'd5159;
      41938:data<=16'd4196;
      41939:data<=16'd3430;
      41940:data<=16'd3698;
      41941:data<=16'd3821;
      41942:data<=16'd4203;
      41943:data<=16'd3648;
      41944:data<=16'd3243;
      41945:data<=16'd3439;
      41946:data<=16'd3096;
      41947:data<=16'd2449;
      41948:data<=16'd1418;
      41949:data<=16'd842;
      41950:data<=16'd981;
      41951:data<=16'd879;
      41952:data<=16'd1301;
      41953:data<=16'd1310;
      41954:data<=16'd215;
      41955:data<=16'd196;
      41956:data<=16'd497;
      41957:data<=16'd70;
      41958:data<=-16'd83;
      41959:data<=-16'd943;
      41960:data<=-16'd2338;
      41961:data<=-16'd2720;
      41962:data<=-16'd2640;
      41963:data<=-16'd2776;
      41964:data<=-16'd2922;
      41965:data<=-16'd2476;
      41966:data<=-16'd1883;
      41967:data<=-16'd2252;
      41968:data<=-16'd2514;
      41969:data<=-16'd2062;
      41970:data<=-16'd1577;
      41971:data<=-16'd1219;
      41972:data<=-16'd2246;
      41973:data<=-16'd3976;
      41974:data<=-16'd4152;
      41975:data<=-16'd3865;
      41976:data<=-16'd3838;
      41977:data<=-16'd3506;
      41978:data<=-16'd3529;
      41979:data<=-16'd3539;
      41980:data<=-16'd3368;
      41981:data<=-16'd3160;
      41982:data<=-16'd2714;
      41983:data<=-16'd2840;
      41984:data<=-16'd2817;
      41985:data<=-16'd4410;
      41986:data<=-16'd11344;
      41987:data<=-16'd17714;
      41988:data<=-16'd17512;
      41989:data<=-16'd15819;
      41990:data<=-16'd15538;
      41991:data<=-16'd14954;
      41992:data<=-16'd14662;
      41993:data<=-16'd14167;
      41994:data<=-16'd13283;
      41995:data<=-16'd12769;
      41996:data<=-16'd12067;
      41997:data<=-16'd12481;
      41998:data<=-16'd13826;
      41999:data<=-16'd13317;
      42000:data<=-16'd12166;
      42001:data<=-16'd12049;
      42002:data<=-16'd11673;
      42003:data<=-16'd11013;
      42004:data<=-16'd10296;
      42005:data<=-16'd9464;
      42006:data<=-16'd9298;
      42007:data<=-16'd8819;
      42008:data<=-16'd7441;
      42009:data<=-16'd7113;
      42010:data<=-16'd7826;
      42011:data<=-16'd7906;
      42012:data<=-16'd7618;
      42013:data<=-16'd7289;
      42014:data<=-16'd6754;
      42015:data<=-16'd6642;
      42016:data<=-16'd6451;
      42017:data<=-16'd5436;
      42018:data<=-16'd4681;
      42019:data<=-16'd4508;
      42020:data<=-16'd4067;
      42021:data<=-16'd3494;
      42022:data<=-16'd3538;
      42023:data<=-16'd4414;
      42024:data<=-16'd4875;
      42025:data<=-16'd4343;
      42026:data<=-16'd4197;
      42027:data<=-16'd3921;
      42028:data<=-16'd3081;
      42029:data<=-16'd3028;
      42030:data<=-16'd2429;
      42031:data<=-16'd1644;
      42032:data<=-16'd2187;
      42033:data<=-16'd1110;
      42034:data<=-16'd769;
      42035:data<=-16'd3034;
      42036:data<=16'd1424;
      42037:data<=16'd10464;
      42038:data<=16'd11720;
      42039:data<=16'd9667;
      42040:data<=16'd10796;
      42041:data<=16'd10696;
      42042:data<=16'd10160;
      42043:data<=16'd10909;
      42044:data<=16'd10323;
      42045:data<=16'd9838;
      42046:data<=16'd10270;
      42047:data<=16'd9633;
      42048:data<=16'd8411;
      42049:data<=16'd7645;
      42050:data<=16'd7359;
      42051:data<=16'd7274;
      42052:data<=16'd7392;
      42053:data<=16'd7514;
      42054:data<=16'd6863;
      42055:data<=16'd6651;
      42056:data<=16'd7222;
      42057:data<=16'd6863;
      42058:data<=16'd6620;
      42059:data<=16'd6256;
      42060:data<=16'd4238;
      42061:data<=16'd3453;
      42062:data<=16'd4250;
      42063:data<=16'd3950;
      42064:data<=16'd3858;
      42065:data<=16'd4411;
      42066:data<=16'd4225;
      42067:data<=16'd4128;
      42068:data<=16'd4328;
      42069:data<=16'd4219;
      42070:data<=16'd4128;
      42071:data<=16'd4087;
      42072:data<=16'd3779;
      42073:data<=16'd3651;
      42074:data<=16'd4071;
      42075:data<=16'd4111;
      42076:data<=16'd4000;
      42077:data<=16'd4332;
      42078:data<=16'd3977;
      42079:data<=16'd3833;
      42080:data<=16'd4124;
      42081:data<=16'd3630;
      42082:data<=16'd3997;
      42083:data<=16'd3600;
      42084:data<=16'd2789;
      42085:data<=16'd5520;
      42086:data<=16'd3093;
      42087:data<=-16'd6604;
      42088:data<=-16'd8763;
      42089:data<=-16'd5799;
      42090:data<=-16'd6845;
      42091:data<=-16'd6293;
      42092:data<=-16'd5157;
      42093:data<=-16'd6260;
      42094:data<=-16'd5180;
      42095:data<=-16'd4388;
      42096:data<=-16'd4999;
      42097:data<=-16'd3824;
      42098:data<=-16'd2526;
      42099:data<=-16'd1826;
      42100:data<=-16'd1421;
      42101:data<=-16'd1495;
      42102:data<=-16'd1090;
      42103:data<=-16'd839;
      42104:data<=-16'd514;
      42105:data<=-16'd168;
      42106:data<=-16'd517;
      42107:data<=-16'd117;
      42108:data<=16'd212;
      42109:data<=16'd594;
      42110:data<=16'd2729;
      42111:data<=16'd3694;
      42112:data<=16'd3171;
      42113:data<=16'd3527;
      42114:data<=16'd3603;
      42115:data<=16'd3568;
      42116:data<=16'd3686;
      42117:data<=16'd3218;
      42118:data<=16'd3316;
      42119:data<=16'd3838;
      42120:data<=16'd3993;
      42121:data<=16'd3971;
      42122:data<=16'd4451;
      42123:data<=16'd5632;
      42124:data<=16'd5882;
      42125:data<=16'd5592;
      42126:data<=16'd5530;
      42127:data<=16'd4986;
      42128:data<=16'd5319;
      42129:data<=16'd5460;
      42130:data<=16'd4990;
      42131:data<=16'd5841;
      42132:data<=16'd5347;
      42133:data<=16'd5213;
      42134:data<=16'd6692;
      42135:data<=16'd5413;
      42136:data<=16'd9329;
      42137:data<=16'd19649;
      42138:data<=16'd21637;
      42139:data<=16'd18765;
      42140:data<=16'd19273;
      42141:data<=16'd18246;
      42142:data<=16'd17340;
      42143:data<=16'd17638;
      42144:data<=16'd16211;
      42145:data<=16'd15747;
      42146:data<=16'd15673;
      42147:data<=16'd15547;
      42148:data<=16'd16718;
      42149:data<=16'd16486;
      42150:data<=16'd15717;
      42151:data<=16'd15653;
      42152:data<=16'd14871;
      42153:data<=16'd14339;
      42154:data<=16'd13576;
      42155:data<=16'd12616;
      42156:data<=16'd12493;
      42157:data<=16'd12019;
      42158:data<=16'd11539;
      42159:data<=16'd10890;
      42160:data<=16'd10329;
      42161:data<=16'd11391;
      42162:data<=16'd11681;
      42163:data<=16'd10941;
      42164:data<=16'd10806;
      42165:data<=16'd9894;
      42166:data<=16'd9473;
      42167:data<=16'd9670;
      42168:data<=16'd8698;
      42169:data<=16'd8229;
      42170:data<=16'd7752;
      42171:data<=16'd6727;
      42172:data<=16'd7370;
      42173:data<=16'd8792;
      42174:data<=16'd9277;
      42175:data<=16'd8771;
      42176:data<=16'd8476;
      42177:data<=16'd8704;
      42178:data<=16'd7659;
      42179:data<=16'd6862;
      42180:data<=16'd6658;
      42181:data<=16'd5476;
      42182:data<=16'd6021;
      42183:data<=16'd5934;
      42184:data<=16'd4325;
      42185:data<=16'd6672;
      42186:data<=16'd4987;
      42187:data<=-16'd4660;
      42188:data<=-16'd8358;
      42189:data<=-16'd6255;
      42190:data<=-16'd6728;
      42191:data<=-16'd6637;
      42192:data<=-16'd6220;
      42193:data<=-16'd6990;
      42194:data<=-16'd6175;
      42195:data<=-16'd5676;
      42196:data<=-16'd6287;
      42197:data<=-16'd5647;
      42198:data<=-16'd4344;
      42199:data<=-16'd3706;
      42200:data<=-16'd3879;
      42201:data<=-16'd3865;
      42202:data<=-16'd3433;
      42203:data<=-16'd3453;
      42204:data<=-16'd3297;
      42205:data<=-16'd3131;
      42206:data<=-16'd3309;
      42207:data<=-16'd2954;
      42208:data<=-16'd3052;
      42209:data<=-16'd3409;
      42210:data<=-16'd2047;
      42211:data<=-16'd240;
      42212:data<=-16'd55;
      42213:data<=-16'd755;
      42214:data<=-16'd813;
      42215:data<=-16'd599;
      42216:data<=-16'd995;
      42217:data<=-16'd1321;
      42218:data<=-16'd1503;
      42219:data<=-16'd1439;
      42220:data<=-16'd934;
      42221:data<=-16'd1409;
      42222:data<=-16'd1391;
      42223:data<=16'd412;
      42224:data<=16'd1124;
      42225:data<=16'd910;
      42226:data<=16'd660;
      42227:data<=-16'd296;
      42228:data<=-16'd100;
      42229:data<=16'd334;
      42230:data<=16'd49;
      42231:data<=16'd488;
      42232:data<=-16'd174;
      42233:data<=-16'd550;
      42234:data<=16'd196;
      42235:data<=-16'd632;
      42236:data<=16'd3336;
      42237:data<=16'd12555;
      42238:data<=16'd15535;
      42239:data<=16'd13676;
      42240:data<=16'd13338;
      42241:data<=16'd12692;
      42242:data<=16'd12167;
      42243:data<=16'd11726;
      42244:data<=16'd10593;
      42245:data<=16'd10469;
      42246:data<=16'd9955;
      42247:data<=16'd9377;
      42248:data<=16'd10455;
      42249:data<=16'd10980;
      42250:data<=16'd10446;
      42251:data<=16'd9532;
      42252:data<=16'd8320;
      42253:data<=16'd7858;
      42254:data<=16'd7582;
      42255:data<=16'd7036;
      42256:data<=16'd6398;
      42257:data<=16'd5582;
      42258:data<=16'd5328;
      42259:data<=16'd4934;
      42260:data<=16'd4614;
      42261:data<=16'd5347;
      42262:data<=16'd5398;
      42263:data<=16'd5107;
      42264:data<=16'd5031;
      42265:data<=16'd3920;
      42266:data<=16'd3563;
      42267:data<=16'd3909;
      42268:data<=16'd3184;
      42269:data<=16'd2670;
      42270:data<=16'd2244;
      42271:data<=16'd1673;
      42272:data<=16'd1685;
      42273:data<=16'd1431;
      42274:data<=16'd1122;
      42275:data<=16'd789;
      42276:data<=16'd426;
      42277:data<=16'd675;
      42278:data<=16'd294;
      42279:data<=-16'd267;
      42280:data<=-16'd522;
      42281:data<=-16'd1357;
      42282:data<=-16'd1111;
      42283:data<=-16'd1178;
      42284:data<=-16'd2403;
      42285:data<=-16'd1986;
      42286:data<=-16'd5087;
      42287:data<=-16'd13649;
      42288:data<=-16'd18192;
      42289:data<=-16'd17591;
      42290:data<=-16'd17241;
      42291:data<=-16'd16944;
      42292:data<=-16'd16483;
      42293:data<=-16'd16137;
      42294:data<=-16'd15640;
      42295:data<=-16'd15703;
      42296:data<=-16'd15549;
      42297:data<=-16'd15197;
      42298:data<=-16'd15960;
      42299:data<=-16'd16819;
      42300:data<=-16'd16351;
      42301:data<=-16'd15297;
      42302:data<=-16'd14909;
      42303:data<=-16'd14883;
      42304:data<=-16'd14487;
      42305:data<=-16'd13738;
      42306:data<=-16'd12892;
      42307:data<=-16'd12815;
      42308:data<=-16'd12988;
      42309:data<=-16'd12182;
      42310:data<=-16'd11996;
      42311:data<=-16'd12789;
      42312:data<=-16'd12842;
      42313:data<=-16'd12768;
      42314:data<=-16'd12718;
      42315:data<=-16'd12104;
      42316:data<=-16'd11782;
      42317:data<=-16'd11477;
      42318:data<=-16'd10951;
      42319:data<=-16'd10912;
      42320:data<=-16'd10859;
      42321:data<=-16'd10329;
      42322:data<=-16'd9831;
      42323:data<=-16'd10267;
      42324:data<=-16'd11367;
      42325:data<=-16'd11207;
      42326:data<=-16'd10185;
      42327:data<=-16'd10149;
      42328:data<=-16'd10241;
      42329:data<=-16'd9624;
      42330:data<=-16'd8887;
      42331:data<=-16'd8329;
      42332:data<=-16'd8554;
      42333:data<=-16'd8516;
      42334:data<=-16'd7224;
      42335:data<=-16'd7671;
      42336:data<=-16'd8144;
      42337:data<=-16'd2344;
      42338:data<=16'd4723;
      42339:data<=16'd5227;
      42340:data<=16'd3827;
      42341:data<=16'd4261;
      42342:data<=16'd4044;
      42343:data<=16'd4018;
      42344:data<=16'd4358;
      42345:data<=16'd3968;
      42346:data<=16'd4090;
      42347:data<=16'd4099;
      42348:data<=16'd3013;
      42349:data<=16'd1853;
      42350:data<=16'd1392;
      42351:data<=16'd1428;
      42352:data<=16'd1046;
      42353:data<=16'd787;
      42354:data<=16'd987;
      42355:data<=16'd669;
      42356:data<=16'd807;
      42357:data<=16'd917;
      42358:data<=16'd243;
      42359:data<=16'd663;
      42360:data<=16'd193;
      42361:data<=-16'd2082;
      42362:data<=-16'd2485;
      42363:data<=-16'd1798;
      42364:data<=-16'd1724;
      42365:data<=-16'd1571;
      42366:data<=-16'd1844;
      42367:data<=-16'd1842;
      42368:data<=-16'd1378;
      42369:data<=-16'd1272;
      42370:data<=-16'd1290;
      42371:data<=-16'd1618;
      42372:data<=-16'd1630;
      42373:data<=-16'd2221;
      42374:data<=-16'd3967;
      42375:data<=-16'd4055;
      42376:data<=-16'd3683;
      42377:data<=-16'd3902;
      42378:data<=-16'd2943;
      42379:data<=-16'd3297;
      42380:data<=-16'd4043;
      42381:data<=-16'd3184;
      42382:data<=-16'd3410;
      42383:data<=-16'd3262;
      42384:data<=-16'd3206;
      42385:data<=-16'd4696;
      42386:data<=-16'd5168;
      42387:data<=-16'd9947;
      42388:data<=-16'd18195;
      42389:data<=-16'd18971;
      42390:data<=-16'd16510;
      42391:data<=-16'd16953;
      42392:data<=-16'd16187;
      42393:data<=-16'd15245;
      42394:data<=-16'd15059;
      42395:data<=-16'd14270;
      42396:data<=-16'd14032;
      42397:data<=-16'd13341;
      42398:data<=-16'd13286;
      42399:data<=-16'd14587;
      42400:data<=-16'd14219;
      42401:data<=-16'd13029;
      42402:data<=-16'd12320;
      42403:data<=-16'd11677;
      42404:data<=-16'd11508;
      42405:data<=-16'd10707;
      42406:data<=-16'd9779;
      42407:data<=-16'd9553;
      42408:data<=-16'd8887;
      42409:data<=-16'd8489;
      42410:data<=-16'd8508;
      42411:data<=-16'd8651;
      42412:data<=-16'd9144;
      42413:data<=-16'd8646;
      42414:data<=-16'd7917;
      42415:data<=-16'd7799;
      42416:data<=-16'd7221;
      42417:data<=-16'd6869;
      42418:data<=-16'd6490;
      42419:data<=-16'd5917;
      42420:data<=-16'd6043;
      42421:data<=-16'd5453;
      42422:data<=-16'd4432;
      42423:data<=-16'd4582;
      42424:data<=-16'd5532;
      42425:data<=-16'd6235;
      42426:data<=-16'd5353;
      42427:data<=-16'd4696;
      42428:data<=-16'd5219;
      42429:data<=-16'd4261;
      42430:data<=-16'd3644;
      42431:data<=-16'd3688;
      42432:data<=-16'd2481;
      42433:data<=-16'd2696;
      42434:data<=-16'd1856;
      42435:data<=-16'd467;
      42436:data<=-16'd3536;
      42437:data<=-16'd710;
      42438:data<=16'd9800;
      42439:data<=16'd12028;
      42440:data<=16'd9157;
      42441:data<=16'd10607;
      42442:data<=16'd10839;
      42443:data<=16'd9785;
      42444:data<=16'd10282;
      42445:data<=16'd9821;
      42446:data<=16'd9680;
      42447:data<=16'd10260;
      42448:data<=16'd9364;
      42449:data<=16'd7914;
      42450:data<=16'd7259;
      42451:data<=16'd7059;
      42452:data<=16'd6634;
      42453:data<=16'd6689;
      42454:data<=16'd7197;
      42455:data<=16'd6689;
      42456:data<=16'd6340;
      42457:data<=16'd6426;
      42458:data<=16'd5788;
      42459:data<=16'd6006;
      42460:data<=16'd6087;
      42461:data<=16'd4390;
      42462:data<=16'd3427;
      42463:data<=16'd3480;
      42464:data<=16'd3398;
      42465:data<=16'd3850;
      42466:data<=16'd4320;
      42467:data<=16'd4176;
      42468:data<=16'd3797;
      42469:data<=16'd3858;
      42470:data<=16'd4191;
      42471:data<=16'd3965;
      42472:data<=16'd3888;
      42473:data<=16'd3759;
      42474:data<=16'd3439;
      42475:data<=16'd4164;
      42476:data<=16'd4040;
      42477:data<=16'd3351;
      42478:data<=16'd4423;
      42479:data<=16'd4582;
      42480:data<=16'd3917;
      42481:data<=16'd4020;
      42482:data<=16'd3541;
      42483:data<=16'd3993;
      42484:data<=16'd3612;
      42485:data<=16'd2513;
      42486:data<=16'd5338;
      42487:data<=16'd3099;
      42488:data<=-16'd7094;
      42489:data<=-16'd9878;
      42490:data<=-16'd6655;
      42491:data<=-16'd7200;
      42492:data<=-16'd7139;
      42493:data<=-16'd6172;
      42494:data<=-16'd6499;
      42495:data<=-16'd5567;
      42496:data<=-16'd5363;
      42497:data<=-16'd5856;
      42498:data<=-16'd4613;
      42499:data<=-16'd3310;
      42500:data<=-16'd2516;
      42501:data<=-16'd2064;
      42502:data<=-16'd2003;
      42503:data<=-16'd1488;
      42504:data<=-16'd1048;
      42505:data<=-16'd748;
      42506:data<=-16'd464;
      42507:data<=-16'd308;
      42508:data<=16'd285;
      42509:data<=16'd306;
      42510:data<=16'd83;
      42511:data<=16'd1283;
      42512:data<=16'd2728;
      42513:data<=16'd3327;
      42514:data<=16'd3134;
      42515:data<=16'd2634;
      42516:data<=16'd2874;
      42517:data<=16'd3218;
      42518:data<=16'd3186;
      42519:data<=16'd3159;
      42520:data<=16'd3030;
      42521:data<=16'd3037;
      42522:data<=16'd2922;
      42523:data<=16'd3615;
      42524:data<=16'd5256;
      42525:data<=16'd5194;
      42526:data<=16'd4629;
      42527:data<=16'd5010;
      42528:data<=16'd4945;
      42529:data<=16'd5648;
      42530:data<=16'd5861;
      42531:data<=16'd4790;
      42532:data<=16'd5325;
      42533:data<=16'd5583;
      42534:data<=16'd5538;
      42535:data<=16'd5900;
      42536:data<=16'd4581;
      42537:data<=16'd9270;
      42538:data<=16'd19741;
      42539:data<=16'd21813;
      42540:data<=16'd18748;
      42541:data<=16'd19340;
      42542:data<=16'd19202;
      42543:data<=16'd18026;
      42544:data<=16'd17564;
      42545:data<=16'd16606;
      42546:data<=16'd16311;
      42547:data<=16'd15753;
      42548:data<=16'd15432;
      42549:data<=16'd16562;
      42550:data<=16'd16451;
      42551:data<=16'd15528;
      42552:data<=16'd15148;
      42553:data<=16'd14645;
      42554:data<=16'd14422;
      42555:data<=16'd13758;
      42556:data<=16'd12904;
      42557:data<=16'd12516;
      42558:data<=16'd11646;
      42559:data<=16'd11122;
      42560:data<=16'd10915;
      42561:data<=16'd10959;
      42562:data<=16'd12002;
      42563:data<=16'd11820;
      42564:data<=16'd10897;
      42565:data<=16'd11094;
      42566:data<=16'd10728;
      42567:data<=16'd10152;
      42568:data<=16'd9705;
      42569:data<=16'd8868;
      42570:data<=16'd8965;
      42571:data<=16'd8771;
      42572:data<=16'd7797;
      42573:data<=16'd7809;
      42574:data<=16'd8645;
      42575:data<=16'd9709;
      42576:data<=16'd9391;
      42577:data<=16'd8255;
      42578:data<=16'd8428;
      42579:data<=16'd7799;
      42580:data<=16'd7056;
      42581:data<=16'd7348;
      42582:data<=16'd6117;
      42583:data<=16'd5586;
      42584:data<=16'd5350;
      42585:data<=16'd4149;
      42586:data<=16'd6282;
      42587:data<=16'd4737;
      42588:data<=-16'd4607;
      42589:data<=-16'd8420;
      42590:data<=-16'd6200;
      42591:data<=-16'd6933;
      42592:data<=-16'd7535;
      42593:data<=-16'd6769;
      42594:data<=-16'd6889;
      42595:data<=-16'd6482;
      42596:data<=-16'd6328;
      42597:data<=-16'd6584;
      42598:data<=-16'd5803;
      42599:data<=-16'd4454;
      42600:data<=-16'd3377;
      42601:data<=-16'd3300;
      42602:data<=-16'd3560;
      42603:data<=-16'd3339;
      42604:data<=-16'd3169;
      42605:data<=-16'd2863;
      42606:data<=-16'd2869;
      42607:data<=-16'd3228;
      42608:data<=-16'd2719;
      42609:data<=-16'd2434;
      42610:data<=-16'd2922;
      42611:data<=-16'd2417;
      42612:data<=-16'd1052;
      42613:data<=-16'd367;
      42614:data<=-16'd508;
      42615:data<=-16'd628;
      42616:data<=-16'd817;
      42617:data<=-16'd1134;
      42618:data<=-16'd782;
      42619:data<=-16'd654;
      42620:data<=-16'd1086;
      42621:data<=-16'd1054;
      42622:data<=-16'd1230;
      42623:data<=-16'd781;
      42624:data<=16'd846;
      42625:data<=16'd1155;
      42626:data<=16'd679;
      42627:data<=16'd845;
      42628:data<=16'd864;
      42629:data<=16'd958;
      42630:data<=16'd564;
      42631:data<=16'd99;
      42632:data<=16'd725;
      42633:data<=16'd840;
      42634:data<=16'd1090;
      42635:data<=16'd1298;
      42636:data<=16'd77;
      42637:data<=16'd3689;
      42638:data<=16'd12478;
      42639:data<=16'd16004;
      42640:data<=16'd14411;
      42641:data<=16'd14026;
      42642:data<=16'd13673;
      42643:data<=16'd12877;
      42644:data<=16'd12477;
      42645:data<=16'd11494;
      42646:data<=16'd11150;
      42647:data<=16'd11145;
      42648:data<=16'd10204;
      42649:data<=16'd10292;
      42650:data<=16'd10854;
      42651:data<=16'd9961;
      42652:data<=16'd9603;
      42653:data<=16'd9791;
      42654:data<=16'd8619;
      42655:data<=16'd7826;
      42656:data<=16'd7887;
      42657:data<=16'd7138;
      42658:data<=16'd6579;
      42659:data<=16'd6420;
      42660:data<=16'd5677;
      42661:data<=16'd5741;
      42662:data<=16'd6593;
      42663:data<=16'd6401;
      42664:data<=16'd5814;
      42665:data<=16'd5767;
      42666:data<=16'd5391;
      42667:data<=16'd4561;
      42668:data<=16'd4049;
      42669:data<=16'd3880;
      42670:data<=16'd3680;
      42671:data<=16'd3348;
      42672:data<=16'd2784;
      42673:data<=16'd2103;
      42674:data<=16'd1804;
      42675:data<=16'd1818;
      42676:data<=16'd1638;
      42677:data<=16'd1394;
      42678:data<=16'd1098;
      42679:data<=16'd293;
      42680:data<=-16'd417;
      42681:data<=-16'd491;
      42682:data<=-16'd707;
      42683:data<=-16'd1133;
      42684:data<=-16'd1586;
      42685:data<=-16'd1962;
      42686:data<=-16'd1666;
      42687:data<=-16'd4223;
      42688:data<=-16'd12157;
      42689:data<=-16'd17895;
      42690:data<=-16'd17296;
      42691:data<=-16'd16601;
      42692:data<=-16'd17120;
      42693:data<=-16'd16383;
      42694:data<=-16'd15832;
      42695:data<=-16'd15467;
      42696:data<=-16'd15091;
      42697:data<=-16'd15186;
      42698:data<=-16'd14680;
      42699:data<=-16'd14786;
      42700:data<=-16'd15555;
      42701:data<=-16'd14865;
      42702:data<=-16'd14319;
      42703:data<=-16'd14600;
      42704:data<=-16'd14204;
      42705:data<=-16'd13872;
      42706:data<=-16'd13452;
      42707:data<=-16'd12668;
      42708:data<=-16'd12480;
      42709:data<=-16'd12011;
      42710:data<=-16'd11350;
      42711:data<=-16'd11879;
      42712:data<=-16'd12621;
      42713:data<=-16'd12383;
      42714:data<=-16'd11671;
      42715:data<=-16'd11365;
      42716:data<=-16'd11696;
      42717:data<=-16'd12019;
      42718:data<=-16'd11731;
      42719:data<=-16'd10886;
      42720:data<=-16'd10173;
      42721:data<=-16'd9969;
      42722:data<=-16'd9611;
      42723:data<=-16'd9047;
      42724:data<=-16'd9279;
      42725:data<=-16'd10426;
      42726:data<=-16'd10906;
      42727:data<=-16'd10072;
      42728:data<=-16'd9815;
      42729:data<=-16'd9964;
      42730:data<=-16'd8896;
      42731:data<=-16'd8184;
      42732:data<=-16'd8116;
      42733:data<=-16'd7667;
      42734:data<=-16'd7638;
      42735:data<=-16'd7066;
      42736:data<=-16'd7150;
      42737:data<=-16'd8176;
      42738:data<=-16'd3140;
      42739:data<=16'd5210;
      42740:data<=16'd6388;
      42741:data<=16'd4393;
      42742:data<=16'd5116;
      42743:data<=16'd5089;
      42744:data<=16'd4567;
      42745:data<=16'd4937;
      42746:data<=16'd4636;
      42747:data<=16'd4576;
      42748:data<=16'd4863;
      42749:data<=16'd3959;
      42750:data<=16'd2446;
      42751:data<=16'd1770;
      42752:data<=16'd1785;
      42753:data<=16'd1442;
      42754:data<=16'd1365;
      42755:data<=16'd1756;
      42756:data<=16'd1704;
      42757:data<=16'd1836;
      42758:data<=16'd1645;
      42759:data<=16'd928;
      42760:data<=16'd1265;
      42761:data<=16'd1052;
      42762:data<=-16'd417;
      42763:data<=-16'd1130;
      42764:data<=-16'd1463;
      42765:data<=-16'd1401;
      42766:data<=-16'd828;
      42767:data<=-16'd769;
      42768:data<=-16'd513;
      42769:data<=-16'd335;
      42770:data<=-16'd585;
      42771:data<=-16'd494;
      42772:data<=-16'd461;
      42773:data<=-16'd182;
      42774:data<=-16'd657;
      42775:data<=-16'd2237;
      42776:data<=-16'd2388;
      42777:data<=-16'd2478;
      42778:data<=-16'd2874;
      42779:data<=-16'd1924;
      42780:data<=-16'd2455;
      42781:data<=-16'd2989;
      42782:data<=-16'd1747;
      42783:data<=-16'd2185;
      42784:data<=-16'd2332;
      42785:data<=-16'd2017;
      42786:data<=-16'd2863;
      42787:data<=-16'd2272;
      42788:data<=-16'd6631;
      42789:data<=-16'd16466;
      42790:data<=-16'd18628;
      42791:data<=-16'd15575;
      42792:data<=-16'd15696;
      42793:data<=-16'd15267;
      42794:data<=-16'd14037;
      42795:data<=-16'd13809;
      42796:data<=-16'd13355;
      42797:data<=-16'd13355;
      42798:data<=-16'd12900;
      42799:data<=-16'd12326;
      42800:data<=-16'd12860;
      42801:data<=-16'd12757;
      42802:data<=-16'd12410;
      42803:data<=-16'd12125;
      42804:data<=-16'd10965;
      42805:data<=-16'd10210;
      42806:data<=-16'd9888;
      42807:data<=-16'd9483;
      42808:data<=-16'd9171;
      42809:data<=-16'd8464;
      42810:data<=-16'd7888;
      42811:data<=-16'd7705;
      42812:data<=-16'd8061;
      42813:data<=-16'd8718;
      42814:data<=-16'd8173;
      42815:data<=-16'd7459;
      42816:data<=-16'd7307;
      42817:data<=-16'd6811;
      42818:data<=-16'd6895;
      42819:data<=-16'd6589;
      42820:data<=-16'd5527;
      42821:data<=-16'd5650;
      42822:data<=-16'd5407;
      42823:data<=-16'd4543;
      42824:data<=-16'd4977;
      42825:data<=-16'd5785;
      42826:data<=-16'd6091;
      42827:data<=-16'd5379;
      42828:data<=-16'd4570;
      42829:data<=-16'd4661;
      42830:data<=-16'd3651;
      42831:data<=-16'd3011;
      42832:data<=-16'd3577;
      42833:data<=-16'd2857;
      42834:data<=-16'd2757;
      42835:data<=-16'd2071;
      42836:data<=-16'd746;
      42837:data<=-16'd3469;
      42838:data<=-16'd1221;
      42839:data<=16'd9371;
      42840:data<=16'd12646;
      42841:data<=16'd9482;
      42842:data<=16'd10205;
      42843:data<=16'd10489;
      42844:data<=16'd9398;
      42845:data<=16'd9858;
      42846:data<=16'd9552;
      42847:data<=16'd9453;
      42848:data<=16'd9996;
      42849:data<=16'd8927;
      42850:data<=16'd7025;
      42851:data<=16'd6026;
      42852:data<=16'd6296;
      42853:data<=16'd6467;
      42854:data<=16'd6187;
      42855:data<=16'd6269;
      42856:data<=16'd5899;
      42857:data<=16'd5821;
      42858:data<=16'd6141;
      42859:data<=16'd5398;
      42860:data<=16'd5416;
      42861:data<=16'd5702;
      42862:data<=16'd4141;
      42863:data<=16'd3005;
      42864:data<=16'd2978;
      42865:data<=16'd2922;
      42866:data<=16'd2943;
      42867:data<=16'd2922;
      42868:data<=16'd3381;
      42869:data<=16'd3535;
      42870:data<=16'd3087;
      42871:data<=16'd3371;
      42872:data<=16'd3383;
      42873:data<=16'd3292;
      42874:data<=16'd3428;
      42875:data<=16'd2754;
      42876:data<=16'd3019;
      42877:data<=16'd3424;
      42878:data<=16'd2848;
      42879:data<=16'd3297;
      42880:data<=16'd3042;
      42881:data<=16'd2540;
      42882:data<=16'd3140;
      42883:data<=16'd2467;
      42884:data<=16'd2784;
      42885:data<=16'd2946;
      42886:data<=16'd1563;
      42887:data<=16'd4291;
      42888:data<=16'd3112;
      42889:data<=-16'd6951;
      42890:data<=-16'd10489;
      42891:data<=-16'd7420;
      42892:data<=-16'd7814;
      42893:data<=-16'd7744;
      42894:data<=-16'd6868;
      42895:data<=-16'd7397;
      42896:data<=-16'd6646;
      42897:data<=-16'd6302;
      42898:data<=-16'd6763;
      42899:data<=-16'd5882;
      42900:data<=-16'd4234;
      42901:data<=-16'd2945;
      42902:data<=-16'd2846;
      42903:data<=-16'd2629;
      42904:data<=-16'd1920;
      42905:data<=-16'd1941;
      42906:data<=-16'd1406;
      42907:data<=-16'd1301;
      42908:data<=-16'd2152;
      42909:data<=-16'd1533;
      42910:data<=-16'd1257;
      42911:data<=-16'd1604;
      42912:data<=-16'd35;
      42913:data<=16'd1542;
      42914:data<=16'd1745;
      42915:data<=16'd1642;
      42916:data<=16'd1736;
      42917:data<=16'd1952;
      42918:data<=16'd1870;
      42919:data<=16'd2079;
      42920:data<=16'd1885;
      42921:data<=16'd1166;
      42922:data<=16'd1694;
      42923:data<=16'd1950;
      42924:data<=16'd2361;
      42925:data<=16'd4220;
      42926:data<=16'd4250;
      42927:data<=16'd3776;
      42928:data<=16'd4508;
      42929:data<=16'd4308;
      42930:data<=16'd4846;
      42931:data<=16'd5142;
      42932:data<=16'd4190;
      42933:data<=16'd4507;
      42934:data<=16'd4081;
      42935:data<=16'd4444;
      42936:data<=16'd5789;
      42937:data<=16'd3873;
      42938:data<=16'd7438;
      42939:data<=16'd17711;
      42940:data<=16'd20334;
      42941:data<=16'd17744;
      42942:data<=16'd17851;
      42943:data<=16'd17415;
      42944:data<=16'd16697;
      42945:data<=16'd16298;
      42946:data<=16'd15399;
      42947:data<=16'd15453;
      42948:data<=16'd15154;
      42949:data<=16'd14985;
      42950:data<=16'd15760;
      42951:data<=16'd15427;
      42952:data<=16'd14798;
      42953:data<=16'd14234;
      42954:data<=16'd13295;
      42955:data<=16'd12928;
      42956:data<=16'd12331;
      42957:data<=16'd11771;
      42958:data<=16'd11673;
      42959:data<=16'd11206;
      42960:data<=16'd10853;
      42961:data<=16'd10041;
      42962:data<=16'd9721;
      42963:data<=16'd11018;
      42964:data<=16'd10953;
      42965:data<=16'd10016;
      42966:data<=16'd10117;
      42967:data<=16'd9697;
      42968:data<=16'd9483;
      42969:data<=16'd9277;
      42970:data<=16'd7982;
      42971:data<=16'd7815;
      42972:data<=16'd8214;
      42973:data<=16'd7523;
      42974:data<=16'd7138;
      42975:data<=16'd7715;
      42976:data<=16'd8475;
      42977:data<=16'd8081;
      42978:data<=16'd7306;
      42979:data<=16'd7435;
      42980:data<=16'd6737;
      42981:data<=16'd6014;
      42982:data<=16'd6184;
      42983:data<=16'd5556;
      42984:data<=16'd5580;
      42985:data<=16'd5010;
      42986:data<=16'd3348;
      42987:data<=16'd5198;
      42988:data<=16'd4334;
      42989:data<=-16'd4103;
      42990:data<=-16'd8798;
      42991:data<=-16'd7488;
      42992:data<=-16'd7656;
      42993:data<=-16'd7967;
      42994:data<=-16'd7371;
      42995:data<=-16'd7350;
      42996:data<=-16'd6780;
      42997:data<=-16'd6613;
      42998:data<=-16'd7169;
      42999:data<=-16'd7030;
      43000:data<=-16'd6253;
      43001:data<=-16'd5113;
      43002:data<=-16'd4313;
      43003:data<=-16'd4108;
      43004:data<=-16'd4090;
      43005:data<=-16'd4237;
      43006:data<=-16'd3874;
      43007:data<=-16'd3642;
      43008:data<=-16'd4184;
      43009:data<=-16'd4021;
      43010:data<=-16'd3573;
      43011:data<=-16'd3609;
      43012:data<=-16'd3068;
      43013:data<=-16'd2144;
      43014:data<=-16'd1495;
      43015:data<=-16'd1357;
      43016:data<=-16'd1701;
      43017:data<=-16'd1914;
      43018:data<=-16'd2076;
      43019:data<=-16'd1956;
      43020:data<=-16'd1491;
      43021:data<=-16'd1459;
      43022:data<=-16'd1565;
      43023:data<=-16'd1941;
      43024:data<=-16'd2181;
      43025:data<=-16'd807;
      43026:data<=16'd669;
      43027:data<=16'd980;
      43028:data<=16'd967;
      43029:data<=16'd470;
      43030:data<=16'd302;
      43031:data<=16'd839;
      43032:data<=16'd937;
      43033:data<=16'd839;
      43034:data<=16'd585;
      43035:data<=16'd584;
      43036:data<=16'd658;
      43037:data<=-16'd274;
      43038:data<=16'd2397;
      43039:data<=16'd10564;
      43040:data<=16'd15550;
      43041:data<=16'd14460;
      43042:data<=16'd13379;
      43043:data<=16'd13415;
      43044:data<=16'd12756;
      43045:data<=16'd12237;
      43046:data<=16'd12022;
      43047:data<=16'd11342;
      43048:data<=16'd10537;
      43049:data<=16'd10349;
      43050:data<=16'd10759;
      43051:data<=16'd11220;
      43052:data<=16'd11018;
      43053:data<=16'd10011;
      43054:data<=16'd9229;
      43055:data<=16'd8968;
      43056:data<=16'd8455;
      43057:data<=16'd7799;
      43058:data<=16'd7468;
      43059:data<=16'd7298;
      43060:data<=16'd6620;
      43061:data<=16'd5513;
      43062:data<=16'd5767;
      43063:data<=16'd7244;
      43064:data<=16'd7515;
      43065:data<=16'd6813;
      43066:data<=16'd6434;
      43067:data<=16'd5961;
      43068:data<=16'd5692;
      43069:data<=16'd5609;
      43070:data<=16'd4814;
      43071:data<=16'd4275;
      43072:data<=16'd4382;
      43073:data<=16'd3961;
      43074:data<=16'd3597;
      43075:data<=16'd3595;
      43076:data<=16'd3045;
      43077:data<=16'd2464;
      43078:data<=16'd2120;
      43079:data<=16'd1841;
      43080:data<=16'd1642;
      43081:data<=16'd772;
      43082:data<=16'd185;
      43083:data<=16'd478;
      43084:data<=16'd14;
      43085:data<=-16'd616;
      43086:data<=-16'd728;
      43087:data<=-16'd843;
      43088:data<=-16'd2247;
      43089:data<=-16'd8755;
      43090:data<=-16'd16346;
      43091:data<=-16'd16800;
      43092:data<=-16'd14979;
      43093:data<=-16'd15747;
      43094:data<=-16'd15383;
      43095:data<=-16'd14915;
      43096:data<=-16'd15000;
      43097:data<=-16'd13864;
      43098:data<=-16'd13620;
      43099:data<=-16'd13714;
      43100:data<=-16'd13602;
      43101:data<=-16'd14921;
      43102:data<=-16'd15136;
      43103:data<=-16'd13769;
      43104:data<=-16'd13353;
      43105:data<=-16'd13215;
      43106:data<=-16'd12736;
      43107:data<=-16'd12287;
      43108:data<=-16'd11864;
      43109:data<=-16'd11661;
      43110:data<=-16'd11264;
      43111:data<=-16'd10746;
      43112:data<=-16'd10933;
      43113:data<=-16'd12093;
      43114:data<=-16'd13021;
      43115:data<=-16'd12440;
      43116:data<=-16'd11649;
      43117:data<=-16'd11376;
      43118:data<=-16'd10947;
      43119:data<=-16'd10854;
      43120:data<=-16'd10489;
      43121:data<=-16'd9837;
      43122:data<=-16'd10026;
      43123:data<=-16'd9905;
      43124:data<=-16'd9373;
      43125:data<=-16'd9662;
      43126:data<=-16'd10516;
      43127:data<=-16'd10913;
      43128:data<=-16'd10066;
      43129:data<=-16'd9650;
      43130:data<=-16'd9694;
      43131:data<=-16'd8470;
      43132:data<=-16'd8469;
      43133:data<=-16'd8660;
      43134:data<=-16'd7062;
      43135:data<=-16'd7236;
      43136:data<=-16'd6902;
      43137:data<=-16'd6328;
      43138:data<=-16'd9218;
      43139:data<=-16'd5494;
      43140:data<=16'd4752;
      43141:data<=16'd6761;
      43142:data<=16'd4513;
      43143:data<=16'd5513;
      43144:data<=16'd5071;
      43145:data<=16'd4358;
      43146:data<=16'd5002;
      43147:data<=16'd4440;
      43148:data<=16'd4150;
      43149:data<=16'd4558;
      43150:data<=16'd4026;
      43151:data<=16'd2605;
      43152:data<=16'd1653;
      43153:data<=16'd1912;
      43154:data<=16'd1710;
      43155:data<=16'd1221;
      43156:data<=16'd1439;
      43157:data<=16'd1101;
      43158:data<=16'd1077;
      43159:data<=16'd1497;
      43160:data<=16'd1022;
      43161:data<=16'd892;
      43162:data<=16'd634;
      43163:data<=-16'd408;
      43164:data<=-16'd672;
      43165:data<=-16'd563;
      43166:data<=-16'd748;
      43167:data<=-16'd1246;
      43168:data<=-16'd1568;
      43169:data<=-16'd996;
      43170:data<=-16'd1025;
      43171:data<=-16'd1198;
      43172:data<=-16'd607;
      43173:data<=-16'd878;
      43174:data<=-16'd698;
      43175:data<=-16'd588;
      43176:data<=-16'd2591;
      43177:data<=-16'd3386;
      43178:data<=-16'd2807;
      43179:data<=-16'd2960;
      43180:data<=-16'd2842;
      43181:data<=-16'd3272;
      43182:data<=-16'd3275;
      43183:data<=-16'd2557;
      43184:data<=-16'd3203;
      43185:data<=-16'd2949;
      43186:data<=-16'd2954;
      43187:data<=-16'd3770;
      43188:data<=-16'd2305;
      43189:data<=-16'd6551;
      43190:data<=-16'd16569;
      43191:data<=-16'd18710;
      43192:data<=-16'd16504;
      43193:data<=-16'd17021;
      43194:data<=-16'd15810;
      43195:data<=-16'd14598;
      43196:data<=-16'd14389;
      43197:data<=-16'd13082;
      43198:data<=-16'd13251;
      43199:data<=-16'd13192;
      43200:data<=-16'd12443;
      43201:data<=-16'd13597;
      43202:data<=-16'd13462;
      43203:data<=-16'd12058;
      43204:data<=-16'd11991;
      43205:data<=-16'd11593;
      43206:data<=-16'd10892;
      43207:data<=-16'd10296;
      43208:data<=-16'd9435;
      43209:data<=-16'd9165;
      43210:data<=-16'd8801;
      43211:data<=-16'd8070;
      43212:data<=-16'd7618;
      43213:data<=-16'd7858;
      43214:data<=-16'd8997;
      43215:data<=-16'd9195;
      43216:data<=-16'd8251;
      43217:data<=-16'd7694;
      43218:data<=-16'd7016;
      43219:data<=-16'd6554;
      43220:data<=-16'd6372;
      43221:data<=-16'd5744;
      43222:data<=-16'd5645;
      43223:data<=-16'd5497;
      43224:data<=-16'd4730;
      43225:data<=-16'd4719;
      43226:data<=-16'd5501;
      43227:data<=-16'd6102;
      43228:data<=-16'd5764;
      43229:data<=-16'd5520;
      43230:data<=-16'd5576;
      43231:data<=-16'd4206;
      43232:data<=-16'd3541;
      43233:data<=-16'd3698;
      43234:data<=-16'd2634;
      43235:data<=-16'd3019;
      43236:data<=-16'd2291;
      43237:data<=-16'd247;
      43238:data<=-16'd2875;
      43239:data<=-16'd890;
      43240:data<=16'd9094;
      43241:data<=16'd11909;
      43242:data<=16'd9699;
      43243:data<=16'd10945;
      43244:data<=16'd10501;
      43245:data<=16'd9646;
      43246:data<=16'd10360;
      43247:data<=16'd9403;
      43248:data<=16'd9359;
      43249:data<=16'd10082;
      43250:data<=16'd9201;
      43251:data<=16'd8146;
      43252:data<=16'd7063;
      43253:data<=16'd6631;
      43254:data<=16'd6757;
      43255:data<=16'd6384;
      43256:data<=16'd6611;
      43257:data<=16'd6579;
      43258:data<=16'd6291;
      43259:data<=16'd6758;
      43260:data<=16'd6434;
      43261:data<=16'd6354;
      43262:data<=16'd6534;
      43263:data<=16'd4942;
      43264:data<=16'd3915;
      43265:data<=16'd4203;
      43266:data<=16'd4094;
      43267:data<=16'd3961;
      43268:data<=16'd3712;
      43269:data<=16'd3595;
      43270:data<=16'd3651;
      43271:data<=16'd3515;
      43272:data<=16'd3911;
      43273:data<=16'd3862;
      43274:data<=16'd3454;
      43275:data<=16'd3879;
      43276:data<=16'd3883;
      43277:data<=16'd3583;
      43278:data<=16'd3385;
      43279:data<=16'd3236;
      43280:data<=16'd3839;
      43281:data<=16'd3641;
      43282:data<=16'd3206;
      43283:data<=16'd3606;
      43284:data<=16'd3102;
      43285:data<=16'd3347;
      43286:data<=16'd3365;
      43287:data<=16'd2108;
      43288:data<=16'd3979;
      43289:data<=16'd2836;
      43290:data<=-16'd5535;
      43291:data<=-16'd9606;
      43292:data<=-16'd8502;
      43293:data<=-16'd8746;
      43294:data<=-16'd7730;
      43295:data<=-16'd6534;
      43296:data<=-16'd6875;
      43297:data<=-16'd6272;
      43298:data<=-16'd5888;
      43299:data<=-16'd5741;
      43300:data<=-16'd4971;
      43301:data<=-16'd4208;
      43302:data<=-16'd2883;
      43303:data<=-16'd2256;
      43304:data<=-16'd2426;
      43305:data<=-16'd2094;
      43306:data<=-16'd2143;
      43307:data<=-16'd1668;
      43308:data<=-16'd884;
      43309:data<=-16'd1268;
      43310:data<=-16'd972;
      43311:data<=-16'd394;
      43312:data<=-16'd614;
      43313:data<=16'd341;
      43314:data<=16'd1823;
      43315:data<=16'd1932;
      43316:data<=16'd1415;
      43317:data<=16'd1670;
      43318:data<=16'd2234;
      43319:data<=16'd2024;
      43320:data<=16'd2200;
      43321:data<=16'd2669;
      43322:data<=16'd2343;
      43323:data<=16'd2531;
      43324:data<=16'd2578;
      43325:data<=16'd2500;
      43326:data<=16'd4094;
      43327:data<=16'd5049;
      43328:data<=16'd4740;
      43329:data<=16'd4726;
      43330:data<=16'd4229;
      43331:data<=16'd4241;
      43332:data<=16'd4742;
      43333:data<=16'd4792;
      43334:data<=16'd5043;
      43335:data<=16'd4467;
      43336:data<=16'd4684;
      43337:data<=16'd5488;
      43338:data<=16'd4284;
      43339:data<=16'd8084;
      43340:data<=16'd17059;
      43341:data<=16'd20048;
      43342:data<=16'd19123;
      43343:data<=16'd19414;
      43344:data<=16'd17929;
      43345:data<=16'd16519;
      43346:data<=16'd16428;
      43347:data<=16'd15826;
      43348:data<=16'd15700;
      43349:data<=16'd15297;
      43350:data<=16'd14697;
      43351:data<=16'd15361;
      43352:data<=16'd15706;
      43353:data<=16'd15057;
      43354:data<=16'd14257;
      43355:data<=16'd13722;
      43356:data<=16'd13265;
      43357:data<=16'd12310;
      43358:data<=16'd11808;
      43359:data<=16'd11737;
      43360:data<=16'd11174;
      43361:data<=16'd10666;
      43362:data<=16'd9791;
      43363:data<=16'd9480;
      43364:data<=16'd10884;
      43365:data<=16'd11298;
      43366:data<=16'd10445;
      43367:data<=16'd10201;
      43368:data<=16'd9643;
      43369:data<=16'd8730;
      43370:data<=16'd8085;
      43371:data<=16'd7527;
      43372:data<=16'd7447;
      43373:data<=16'd7235;
      43374:data<=16'd6513;
      43375:data<=16'd6384;
      43376:data<=16'd7332;
      43377:data<=16'd8231;
      43378:data<=16'd7653;
      43379:data<=16'd6818;
      43380:data<=16'd7033;
      43381:data<=16'd6733;
      43382:data<=16'd5877;
      43383:data<=16'd5366;
      43384:data<=16'd4901;
      43385:data<=16'd5012;
      43386:data<=16'd4469;
      43387:data<=16'd3175;
      43388:data<=16'd4250;
      43389:data<=16'd3780;
      43390:data<=-16'd3090;
      43391:data<=-16'd9138;
      43392:data<=-16'd9100;
      43393:data<=-16'd8129;
      43394:data<=-16'd8288;
      43395:data<=-16'd8100;
      43396:data<=-16'd8173;
      43397:data<=-16'd7932;
      43398:data<=-16'd7544;
      43399:data<=-16'd8040;
      43400:data<=-16'd7776;
      43401:data<=-16'd6408;
      43402:data<=-16'd5486;
      43403:data<=-16'd5081;
      43404:data<=-16'd4877;
      43405:data<=-16'd4710;
      43406:data<=-16'd4764;
      43407:data<=-16'd4919;
      43408:data<=-16'd4493;
      43409:data<=-16'd4256;
      43410:data<=-16'd4134;
      43411:data<=-16'd3744;
      43412:data<=-16'd4329;
      43413:data<=-16'd4038;
      43414:data<=-16'd1971;
      43415:data<=-16'd1650;
      43416:data<=-16'd2491;
      43417:data<=-16'd2029;
      43418:data<=-16'd1538;
      43419:data<=-16'd1615;
      43420:data<=-16'd1902;
      43421:data<=-16'd2331;
      43422:data<=-16'd2325;
      43423:data<=-16'd1936;
      43424:data<=-16'd1741;
      43425:data<=-16'd1923;
      43426:data<=-16'd1400;
      43427:data<=-16'd217;
      43428:data<=-16'd91;
      43429:data<=-16'd77;
      43430:data<=16'd162;
      43431:data<=-16'd411;
      43432:data<=-16'd165;
      43433:data<=16'd162;
      43434:data<=-16'd567;
      43435:data<=-16'd381;
      43436:data<=-16'd58;
      43437:data<=-16'd188;
      43438:data<=16'd0;
      43439:data<=16'd1554;
      43440:data<=16'd7756;
      43441:data<=16'd14222;
      43442:data<=16'd14612;
      43443:data<=16'd13750;
      43444:data<=16'd13749;
      43445:data<=16'd12225;
      43446:data<=16'd11429;
      43447:data<=16'd11127;
      43448:data<=16'd10759;
      43449:data<=16'd10815;
      43450:data<=16'd9588;
      43451:data<=16'd9451;
      43452:data<=16'd10956;
      43453:data<=16'd10593;
      43454:data<=16'd9865;
      43455:data<=16'd9699;
      43456:data<=16'd8901;
      43457:data<=16'd8416;
      43458:data<=16'd7749;
      43459:data<=16'd6980;
      43460:data<=16'd6678;
      43461:data<=16'd5927;
      43462:data<=16'd5360;
      43463:data<=16'd5238;
      43464:data<=16'd5595;
      43465:data<=16'd6602;
      43466:data<=16'd6592;
      43467:data<=16'd6049;
      43468:data<=16'd5836;
      43469:data<=16'd4975;
      43470:data<=16'd4449;
      43471:data<=16'd4434;
      43472:data<=16'd4222;
      43473:data<=16'd4087;
      43474:data<=16'd3169;
      43475:data<=16'd2244;
      43476:data<=16'd2326;
      43477:data<=16'd2253;
      43478:data<=16'd1999;
      43479:data<=16'd1538;
      43480:data<=16'd1348;
      43481:data<=16'd1674;
      43482:data<=16'd748;
      43483:data<=-16'd41;
      43484:data<=16'd59;
      43485:data<=-16'd493;
      43486:data<=-16'd138;
      43487:data<=-16'd550;
      43488:data<=-16'd2191;
      43489:data<=-16'd1988;
      43490:data<=-16'd6205;
      43491:data<=-16'd14929;
      43492:data<=-16'd16895;
      43493:data<=-16'd15068;
      43494:data<=-16'd15805;
      43495:data<=-16'd15151;
      43496:data<=-16'd13955;
      43497:data<=-16'd14019;
      43498:data<=-16'd13687;
      43499:data<=-16'd13684;
      43500:data<=-16'd13109;
      43501:data<=-16'd12718;
      43502:data<=-16'd14190;
      43503:data<=-16'd14387;
      43504:data<=-16'd13280;
      43505:data<=-16'd13063;
      43506:data<=-16'd12669;
      43507:data<=-16'd12251;
      43508:data<=-16'd11949;
      43509:data<=-16'd11203;
      43510:data<=-16'd10778;
      43511:data<=-16'd10473;
      43512:data<=-16'd10125;
      43513:data<=-16'd10176;
      43514:data<=-16'd10683;
      43515:data<=-16'd11338;
      43516:data<=-16'd11136;
      43517:data<=-16'd10569;
      43518:data<=-16'd10316;
      43519:data<=-16'd9617;
      43520:data<=-16'd9088;
      43521:data<=-16'd8786;
      43522:data<=-16'd8346;
      43523:data<=-16'd8540;
      43524:data<=-16'd8175;
      43525:data<=-16'd7254;
      43526:data<=-16'd7958;
      43527:data<=-16'd9508;
      43528:data<=-16'd9688;
      43529:data<=-16'd8366;
      43530:data<=-16'd7861;
      43531:data<=-16'd8328;
      43532:data<=-16'd7316;
      43533:data<=-16'd6584;
      43534:data<=-16'd6678;
      43535:data<=-16'd5858;
      43536:data<=-16'd6366;
      43537:data<=-16'd6044;
      43538:data<=-16'd4866;
      43539:data<=-16'd7571;
      43540:data<=-16'd5037;
      43541:data<=16'd5056;
      43542:data<=16'd7783;
      43543:data<=16'd5668;
      43544:data<=16'd7074;
      43545:data<=16'd6402;
      43546:data<=16'd5143;
      43547:data<=16'd6093;
      43548:data<=16'd5248;
      43549:data<=16'd5021;
      43550:data<=16'd6126;
      43551:data<=16'd4877;
      43552:data<=16'd2957;
      43553:data<=16'd2537;
      43554:data<=16'd2902;
      43555:data<=16'd2890;
      43556:data<=16'd2485;
      43557:data<=16'd2461;
      43558:data<=16'd2011;
      43559:data<=16'd1488;
      43560:data<=16'd1665;
      43561:data<=16'd1569;
      43562:data<=16'd1776;
      43563:data<=16'd1760;
      43564:data<=16'd308;
      43565:data<=-16'd640;
      43566:data<=-16'd663;
      43567:data<=-16'd705;
      43568:data<=-16'd534;
      43569:data<=-16'd629;
      43570:data<=-16'd741;
      43571:data<=-16'd619;
      43572:data<=-16'd846;
      43573:data<=-16'd1222;
      43574:data<=-16'd1293;
      43575:data<=-16'd529;
      43576:data<=-16'd494;
      43577:data<=-16'd2379;
      43578:data<=-16'd3237;
      43579:data<=-16'd2913;
      43580:data<=-16'd3143;
      43581:data<=-16'd2931;
      43582:data<=-16'd2911;
      43583:data<=-16'd2857;
      43584:data<=-16'd2378;
      43585:data<=-16'd3016;
      43586:data<=-16'd2971;
      43587:data<=-16'd2711;
      43588:data<=-16'd3160;
      43589:data<=-16'd2309;
      43590:data<=-16'd6599;
      43591:data<=-16'd16060;
      43592:data<=-16'd18289;
      43593:data<=-16'd16137;
      43594:data<=-16'd16927;
      43595:data<=-16'd15908;
      43596:data<=-16'd14026;
      43597:data<=-16'd14308;
      43598:data<=-16'd14360;
      43599:data<=-16'd14085;
      43600:data<=-16'd12932;
      43601:data<=-16'd12057;
      43602:data<=-16'd13333;
      43603:data<=-16'd13573;
      43604:data<=-16'd12656;
      43605:data<=-16'd12320;
      43606:data<=-16'd11421;
      43607:data<=-16'd10662;
      43608:data<=-16'd9967;
      43609:data<=-16'd8915;
      43610:data<=-16'd8642;
      43611:data<=-16'd8351;
      43612:data<=-16'd7720;
      43613:data<=-16'd7166;
      43614:data<=-16'd7292;
      43615:data<=-16'd8627;
      43616:data<=-16'd8610;
      43617:data<=-16'd7600;
      43618:data<=-16'd7885;
      43619:data<=-16'd7453;
      43620:data<=-16'd6714;
      43621:data<=-16'd6399;
      43622:data<=-16'd5131;
      43623:data<=-16'd5109;
      43624:data<=-16'd5401;
      43625:data<=-16'd4046;
      43626:data<=-16'd4340;
      43627:data<=-16'd5799;
      43628:data<=-16'd5735;
      43629:data<=-16'd5051;
      43630:data<=-16'd4681;
      43631:data<=-16'd4595;
      43632:data<=-16'd3973;
      43633:data<=-16'd3583;
      43634:data<=-16'd3601;
      43635:data<=-16'd2487;
      43636:data<=-16'd2519;
      43637:data<=-16'd2458;
      43638:data<=-16'd890;
      43639:data<=-16'd2710;
      43640:data<=-16'd1001;
      43641:data<=16'd8619;
      43642:data<=16'd11981;
      43643:data<=16'd9395;
      43644:data<=16'd10499;
      43645:data<=16'd10569;
      43646:data<=16'd9533;
      43647:data<=16'd10434;
      43648:data<=16'd10034;
      43649:data<=16'd9797;
      43650:data<=16'd10144;
      43651:data<=16'd9060;
      43652:data<=16'd7849;
      43653:data<=16'd6975;
      43654:data<=16'd7130;
      43655:data<=16'd7251;
      43656:data<=16'd6150;
      43657:data<=16'd6328;
      43658:data<=16'd6454;
      43659:data<=16'd5733;
      43660:data<=16'd6291;
      43661:data<=16'd5862;
      43662:data<=16'd5033;
      43663:data<=16'd5603;
      43664:data<=16'd4863;
      43665:data<=16'd3648;
      43666:data<=16'd3412;
      43667:data<=16'd3259;
      43668:data<=16'd3504;
      43669:data<=16'd3319;
      43670:data<=16'd3201;
      43671:data<=16'd3709;
      43672:data<=16'd3301;
      43673:data<=16'd3122;
      43674:data<=16'd3236;
      43675:data<=16'd2611;
      43676:data<=16'd2796;
      43677:data<=16'd3236;
      43678:data<=16'd3295;
      43679:data<=16'd3610;
      43680:data<=16'd3407;
      43681:data<=16'd3090;
      43682:data<=16'd3058;
      43683:data<=16'd3374;
      43684:data<=16'd3811;
      43685:data<=16'd3297;
      43686:data<=16'd3312;
      43687:data<=16'd3162;
      43688:data<=16'd2326;
      43689:data<=16'd4252;
      43690:data<=16'd2964;
      43691:data<=-16'd5318;
      43692:data<=-16'd9409;
      43693:data<=-16'd8113;
      43694:data<=-16'd8366;
      43695:data<=-16'd7688;
      43696:data<=-16'd6197;
      43697:data<=-16'd6285;
      43698:data<=-16'd6284;
      43699:data<=-16'd6548;
      43700:data<=-16'd6505;
      43701:data<=-16'd5330;
      43702:data<=-16'd3971;
      43703:data<=-16'd2417;
      43704:data<=-16'd2155;
      43705:data<=-16'd2645;
      43706:data<=-16'd2012;
      43707:data<=-16'd1848;
      43708:data<=-16'd1439;
      43709:data<=-16'd553;
      43710:data<=-16'd1121;
      43711:data<=-16'd892;
      43712:data<=16'd3;
      43713:data<=-16'd431;
      43714:data<=16'd214;
      43715:data<=16'd1727;
      43716:data<=16'd2238;
      43717:data<=16'd2461;
      43718:data<=16'd2376;
      43719:data<=16'd2241;
      43720:data<=16'd2366;
      43721:data<=16'd2607;
      43722:data<=16'd3174;
      43723:data<=16'd3098;
      43724:data<=16'd2725;
      43725:data<=16'd2940;
      43726:data<=16'd3257;
      43727:data<=16'd4349;
      43728:data<=16'd5190;
      43729:data<=16'd4601;
      43730:data<=16'd4541;
      43731:data<=16'd4911;
      43732:data<=16'd4986;
      43733:data<=16'd5184;
      43734:data<=16'd4746;
      43735:data<=16'd4405;
      43736:data<=16'd4404;
      43737:data<=16'd4306;
      43738:data<=16'd4531;
      43739:data<=16'd4170;
      43740:data<=16'd7162;
      43741:data<=16'd15561;
      43742:data<=16'd19946;
      43743:data<=16'd18609;
      43744:data<=16'd18647;
      43745:data<=16'd18390;
      43746:data<=16'd16769;
      43747:data<=16'd16601;
      43748:data<=16'd16357;
      43749:data<=16'd15834;
      43750:data<=16'd15553;
      43751:data<=16'd14777;
      43752:data<=16'd14819;
      43753:data<=16'd15286;
      43754:data<=16'd14942;
      43755:data<=16'd14468;
      43756:data<=16'd13982;
      43757:data<=16'd13423;
      43758:data<=16'd12504;
      43759:data<=16'd11351;
      43760:data<=16'd11036;
      43761:data<=16'd10974;
      43762:data<=16'd10248;
      43763:data<=16'd9518;
      43764:data<=16'd9946;
      43765:data<=16'd11035;
      43766:data<=16'd10516;
      43767:data<=16'd9448;
      43768:data<=16'd9823;
      43769:data<=16'd9530;
      43770:data<=16'd8373;
      43771:data<=16'd7865;
      43772:data<=16'd7172;
      43773:data<=16'd6719;
      43774:data<=16'd6692;
      43775:data<=16'd6100;
      43776:data<=16'd5768;
      43777:data<=16'd6329;
      43778:data<=16'd7351;
      43779:data<=16'd7655;
      43780:data<=16'd6828;
      43781:data<=16'd6328;
      43782:data<=16'd5829;
      43783:data<=16'd5254;
      43784:data<=16'd5416;
      43785:data<=16'd4871;
      43786:data<=16'd4679;
      43787:data<=16'd5075;
      43788:data<=16'd3707;
      43789:data<=16'd4047;
      43790:data<=16'd4604;
      43791:data<=-16'd1815;
      43792:data<=-16'd8586;
      43793:data<=-16'd8598;
      43794:data<=-16'd8085;
      43795:data<=-16'd8986;
      43796:data<=-16'd8396;
      43797:data<=-16'd7965;
      43798:data<=-16'd8032;
      43799:data<=-16'd7765;
      43800:data<=-16'd8029;
      43801:data<=-16'd8296;
      43802:data<=-16'd7274;
      43803:data<=-16'd5567;
      43804:data<=-16'd5119;
      43805:data<=-16'd5538;
      43806:data<=-16'd5084;
      43807:data<=-16'd4801;
      43808:data<=-16'd5025;
      43809:data<=-16'd4696;
      43810:data<=-16'd4690;
      43811:data<=-16'd4614;
      43812:data<=-16'd4023;
      43813:data<=-16'd4335;
      43814:data<=-16'd4293;
      43815:data<=-16'd2931;
      43816:data<=-16'd2161;
      43817:data<=-16'd2223;
      43818:data<=-16'd2305;
      43819:data<=-16'd2262;
      43820:data<=-16'd2290;
      43821:data<=-16'd2347;
      43822:data<=-16'd1750;
      43823:data<=-16'd1556;
      43824:data<=-16'd2064;
      43825:data<=-16'd1807;
      43826:data<=-16'd1997;
      43827:data<=-16'd1949;
      43828:data<=-16'd293;
      43829:data<=-16'd265;
      43830:data<=-16'd990;
      43831:data<=-16'd30;
      43832:data<=16'd79;
      43833:data<=-16'd446;
      43834:data<=-16'd723;
      43835:data<=-16'd1016;
      43836:data<=-16'd335;
      43837:data<=-16'd678;
      43838:data<=-16'd1225;
      43839:data<=-16'd270;
      43840:data<=16'd466;
      43841:data<=16'd5600;
      43842:data<=16'd13497;
      43843:data<=16'd14228;
      43844:data<=16'd12411;
      43845:data<=16'd13133;
      43846:data<=16'd12022;
      43847:data<=16'd11182;
      43848:data<=16'd11169;
      43849:data<=16'd9962;
      43850:data<=16'd9902;
      43851:data<=16'd9544;
      43852:data<=16'd9013;
      43853:data<=16'd10260;
      43854:data<=16'd10340;
      43855:data<=16'd9520;
      43856:data<=16'd9183;
      43857:data<=16'd8405;
      43858:data<=16'd7884;
      43859:data<=16'd7072;
      43860:data<=16'd6297;
      43861:data<=16'd6166;
      43862:data<=16'd5328;
      43863:data<=16'd5128;
      43864:data<=16'd5890;
      43865:data<=16'd6458;
      43866:data<=16'd6883;
      43867:data<=16'd5935;
      43868:data<=16'd5289;
      43869:data<=16'd5949;
      43870:data<=16'd5238;
      43871:data<=16'd4314;
      43872:data<=16'd3598;
      43873:data<=16'd2513;
      43874:data<=16'd2840;
      43875:data<=16'd2775;
      43876:data<=16'd2253;
      43877:data<=16'd2672;
      43878:data<=16'd2003;
      43879:data<=16'd1639;
      43880:data<=16'd1738;
      43881:data<=16'd795;
      43882:data<=16'd876;
      43883:data<=16'd634;
      43884:data<=-16'd68;
      43885:data<=16'd39;
      43886:data<=-16'd1222;
      43887:data<=-16'd1242;
      43888:data<=-16'd376;
      43889:data<=-16'd1489;
      43890:data<=-16'd1469;
      43891:data<=-16'd5709;
      43892:data<=-16'd15150;
      43893:data<=-16'd17320;
      43894:data<=-16'd15126;
      43895:data<=-16'd15954;
      43896:data<=-16'd15484;
      43897:data<=-16'd14800;
      43898:data<=-16'd15114;
      43899:data<=-16'd14254;
      43900:data<=-16'd13966;
      43901:data<=-16'd13490;
      43902:data<=-16'd13220;
      43903:data<=-16'd14563;
      43904:data<=-16'd14879;
      43905:data<=-16'd14424;
      43906:data<=-16'd13888;
      43907:data<=-16'd12862;
      43908:data<=-16'd12704;
      43909:data<=-16'd12367;
      43910:data<=-16'd11734;
      43911:data<=-16'd11565;
      43912:data<=-16'd10684;
      43913:data<=-16'd10231;
      43914:data<=-16'd10569;
      43915:data<=-16'd11113;
      43916:data<=-16'd12019;
      43917:data<=-16'd11479;
      43918:data<=-16'd10616;
      43919:data<=-16'd10590;
      43920:data<=-16'd9652;
      43921:data<=-16'd9538;
      43922:data<=-16'd9900;
      43923:data<=-16'd8830;
      43924:data<=-16'd8560;
      43925:data<=-16'd8432;
      43926:data<=-16'd7703;
      43927:data<=-16'd8405;
      43928:data<=-16'd9585;
      43929:data<=-16'd10040;
      43930:data<=-16'd9365;
      43931:data<=-16'd8379;
      43932:data<=-16'd8196;
      43933:data<=-16'd7303;
      43934:data<=-16'd7228;
      43935:data<=-16'd7870;
      43936:data<=-16'd6322;
      43937:data<=-16'd6137;
      43938:data<=-16'd6437;
      43939:data<=-16'd5304;
      43940:data<=-16'd7498;
      43941:data<=-16'd5385;
      43942:data<=16'd4475;
      43943:data<=16'd7659;
      43944:data<=16'd5453;
      43945:data<=16'd6540;
      43946:data<=16'd6144;
      43947:data<=16'd5007;
      43948:data<=16'd5855;
      43949:data<=16'd5498;
      43950:data<=16'd5315;
      43951:data<=16'd5645;
      43952:data<=16'd4569;
      43953:data<=16'd3283;
      43954:data<=16'd2541;
      43955:data<=16'd2560;
      43956:data<=16'd2561;
      43957:data<=16'd2079;
      43958:data<=16'd2264;
      43959:data<=16'd2158;
      43960:data<=16'd1889;
      43961:data<=16'd2367;
      43962:data<=16'd2176;
      43963:data<=16'd2106;
      43964:data<=16'd2319;
      43965:data<=16'd1128;
      43966:data<=-16'd42;
      43967:data<=-16'd396;
      43968:data<=-16'd596;
      43969:data<=-16'd425;
      43970:data<=-16'd320;
      43971:data<=-16'd215;
      43972:data<=-16'd35;
      43973:data<=-16'd141;
      43974:data<=-16'd232;
      43975:data<=-16'd165;
      43976:data<=16'd300;
      43977:data<=-16'd118;
      43978:data<=-16'd1785;
      43979:data<=-16'd1883;
      43980:data<=-16'd1400;
      43981:data<=-16'd2118;
      43982:data<=-16'd2174;
      43983:data<=-16'd2064;
      43984:data<=-16'd1973;
      43985:data<=-16'd1598;
      43986:data<=-16'd2043;
      43987:data<=-16'd1647;
      43988:data<=-16'd1583;
      43989:data<=-16'd2262;
      43990:data<=-16'd1037;
      43991:data<=-16'd5028;
      43992:data<=-16'd14716;
      43993:data<=-16'd17273;
      43994:data<=-16'd14979;
      43995:data<=-16'd15418;
      43996:data<=-16'd14816;
      43997:data<=-16'd13571;
      43998:data<=-16'd13399;
      43999:data<=-16'd12469;
      44000:data<=-16'd11981;
      44001:data<=-16'd11571;
      44002:data<=-16'd11350;
      44003:data<=-16'd12266;
      44004:data<=-16'd11984;
      44005:data<=-16'd11124;
      44006:data<=-16'd10840;
      44007:data<=-16'd9934;
      44008:data<=-16'd9409;
      44009:data<=-16'd9074;
      44010:data<=-16'd8272;
      44011:data<=-16'd7961;
      44012:data<=-16'd7644;
      44013:data<=-16'd7238;
      44014:data<=-16'd6716;
      44015:data<=-16'd6428;
      44016:data<=-16'd7338;
      44017:data<=-16'd7304;
      44018:data<=-16'd6376;
      44019:data<=-16'd6687;
      44020:data<=-16'd6373;
      44021:data<=-16'd5509;
      44022:data<=-16'd5321;
      44023:data<=-16'd4390;
      44024:data<=-16'd3768;
      44025:data<=-16'd4106;
      44026:data<=-16'd3823;
      44027:data<=-16'd3501;
      44028:data<=-16'd4252;
      44029:data<=-16'd5251;
      44030:data<=-16'd4772;
      44031:data<=-16'd3883;
      44032:data<=-16'd3933;
      44033:data<=-16'd2857;
      44034:data<=-16'd2077;
      44035:data<=-16'd2766;
      44036:data<=-16'd1944;
      44037:data<=-16'd1407;
      44038:data<=-16'd1105;
      44039:data<=-16'd5;
      44040:data<=-16'd2193;
      44041:data<=-16'd805;
      44042:data<=16'd8335;
      44043:data<=16'd11981;
      44044:data<=16'd9797;
      44045:data<=16'd10712;
      44046:data<=16'd11132;
      44047:data<=16'd10235;
      44048:data<=16'd10257;
      44049:data<=16'd9362;
      44050:data<=16'd9098;
      44051:data<=16'd9388;
      44052:data<=16'd8575;
      44053:data<=16'd7642;
      44054:data<=16'd6351;
      44055:data<=16'd5591;
      44056:data<=16'd5935;
      44057:data<=16'd5949;
      44058:data<=16'd5839;
      44059:data<=16'd5576;
      44060:data<=16'd5750;
      44061:data<=16'd6385;
      44062:data<=16'd5630;
      44063:data<=16'd5298;
      44064:data<=16'd5891;
      44065:data<=16'd4816;
      44066:data<=16'd3579;
      44067:data<=16'd3277;
      44068:data<=16'd2995;
      44069:data<=16'd3128;
      44070:data<=16'd3256;
      44071:data<=16'd3363;
      44072:data<=16'd3466;
      44073:data<=16'd3230;
      44074:data<=16'd3479;
      44075:data<=16'd3647;
      44076:data<=16'd3425;
      44077:data<=16'd3334;
      44078:data<=16'd3240;
      44079:data<=16'd3865;
      44080:data<=16'd4088;
      44081:data<=16'd3720;
      44082:data<=16'd4479;
      44083:data<=16'd4255;
      44084:data<=16'd3582;
      44085:data<=16'd4270;
      44086:data<=16'd3680;
      44087:data<=16'd3277;
      44088:data<=16'd3303;
      44089:data<=16'd2127;
      44090:data<=16'd3899;
      44091:data<=16'd3657;
      44092:data<=-16'd4121;
      44093:data<=-16'd8818;
      44094:data<=-16'd7609;
      44095:data<=-16'd7639;
      44096:data<=-16'd7507;
      44097:data<=-16'd6448;
      44098:data<=-16'd6199;
      44099:data<=-16'd5526;
      44100:data<=-16'd5019;
      44101:data<=-16'd4965;
      44102:data<=-16'd4654;
      44103:data<=-16'd3930;
      44104:data<=-16'd2390;
      44105:data<=-16'd1424;
      44106:data<=-16'd1216;
      44107:data<=-16'd767;
      44108:data<=-16'd958;
      44109:data<=-16'd987;
      44110:data<=-16'd490;
      44111:data<=-16'd881;
      44112:data<=-16'd884;
      44113:data<=-16'd80;
      44114:data<=16'd38;
      44115:data<=16'd320;
      44116:data<=16'd1525;
      44117:data<=16'd2479;
      44118:data<=16'd2491;
      44119:data<=16'd2387;
      44120:data<=16'd2705;
      44121:data<=16'd2608;
      44122:data<=16'd2414;
      44123:data<=16'd2980;
      44124:data<=16'd3435;
      44125:data<=16'd3459;
      44126:data<=16'd3242;
      44127:data<=16'd2895;
      44128:data<=16'd3600;
      44129:data<=16'd4807;
      44130:data<=16'd4951;
      44131:data<=16'd4769;
      44132:data<=16'd4778;
      44133:data<=16'd4752;
      44134:data<=16'd4889;
      44135:data<=16'd4640;
      44136:data<=16'd4261;
      44137:data<=16'd4440;
      44138:data<=16'd4877;
      44139:data<=16'd5201;
      44140:data<=16'd4670;
      44141:data<=16'd6443;
      44142:data<=16'd14034;
      44143:data<=16'd19926;
      44144:data<=16'd19030;
      44145:data<=16'd18268;
      44146:data<=16'd18289;
      44147:data<=16'd16521;
      44148:data<=16'd16451;
      44149:data<=16'd16345;
      44150:data<=16'd14827;
      44151:data<=16'd14684;
      44152:data<=16'd13928;
      44153:data<=16'd13424;
      44154:data<=16'd14675;
      44155:data<=16'd13928;
      44156:data<=16'd12792;
      44157:data<=16'd13051;
      44158:data<=16'd12149;
      44159:data<=16'd11321;
      44160:data<=16'd11051;
      44161:data<=16'd10671;
      44162:data<=16'd10904;
      44163:data<=16'd10129;
      44164:data<=16'd8862;
      44165:data<=16'd8971;
      44166:data<=16'd9688;
      44167:data<=16'd10361;
      44168:data<=16'd9920;
      44169:data<=16'd9036;
      44170:data<=16'd8922;
      44171:data<=16'd8034;
      44172:data<=16'd7526;
      44173:data<=16'd7787;
      44174:data<=16'd6702;
      44175:data<=16'd6235;
      44176:data<=16'd6343;
      44177:data<=16'd5250;
      44178:data<=16'd5595;
      44179:data<=16'd7297;
      44180:data<=16'd7498;
      44181:data<=16'd6581;
      44182:data<=16'd6156;
      44183:data<=16'd6169;
      44184:data<=16'd5771;
      44185:data<=16'd5761;
      44186:data<=16'd5706;
      44187:data<=16'd4658;
      44188:data<=16'd4364;
      44189:data<=16'd3756;
      44190:data<=16'd3548;
      44191:data<=16'd5247;
      44192:data<=16'd933;
      44193:data<=-16'd7753;
      44194:data<=-16'd9030;
      44195:data<=-16'd7271;
      44196:data<=-16'd8150;
      44197:data<=-16'd7530;
      44198:data<=-16'd6912;
      44199:data<=-16'd7056;
      44200:data<=-16'd6422;
      44201:data<=-16'd6890;
      44202:data<=-16'd7335;
      44203:data<=-16'd6686;
      44204:data<=-16'd5503;
      44205:data<=-16'd4262;
      44206:data<=-16'd4678;
      44207:data<=-16'd4827;
      44208:data<=-16'd4009;
      44209:data<=-16'd4575;
      44210:data<=-16'd4548;
      44211:data<=-16'd4035;
      44212:data<=-16'd4648;
      44213:data<=-16'd4352;
      44214:data<=-16'd4020;
      44215:data<=-16'd4049;
      44216:data<=-16'd2652;
      44217:data<=-16'd1677;
      44218:data<=-16'd2150;
      44219:data<=-16'd2549;
      44220:data<=-16'd2061;
      44221:data<=-16'd1481;
      44222:data<=-16'd1892;
      44223:data<=-16'd1894;
      44224:data<=-16'd1369;
      44225:data<=-16'd1621;
      44226:data<=-16'd1883;
      44227:data<=-16'd2346;
      44228:data<=-16'd1851;
      44229:data<=16'd52;
      44230:data<=-16'd61;
      44231:data<=-16'd864;
      44232:data<=-16'd525;
      44233:data<=-16'd758;
      44234:data<=-16'd434;
      44235:data<=-16'd567;
      44236:data<=-16'd1436;
      44237:data<=-16'd814;
      44238:data<=-16'd1222;
      44239:data<=-16'd1286;
      44240:data<=-16'd223;
      44241:data<=-16'd1260;
      44242:data<=16'd3303;
      44243:data<=16'd12953;
      44244:data<=16'd14243;
      44245:data<=16'd11500;
      44246:data<=16'd12137;
      44247:data<=16'd11377;
      44248:data<=16'd10414;
      44249:data<=16'd10827;
      44250:data<=16'd10082;
      44251:data<=16'd9433;
      44252:data<=16'd9066;
      44253:data<=16'd9098;
      44254:data<=16'd9875;
      44255:data<=16'd9462;
      44256:data<=16'd8630;
      44257:data<=16'd8410;
      44258:data<=16'd8175;
      44259:data<=16'd7971;
      44260:data<=16'd7282;
      44261:data<=16'd6645;
      44262:data<=16'd6308;
      44263:data<=16'd5544;
      44264:data<=16'd5236;
      44265:data<=16'd5169;
      44266:data<=16'd5339;
      44267:data<=16'd6211;
      44268:data<=16'd5959;
      44269:data<=16'd4869;
      44270:data<=16'd4306;
      44271:data<=16'd3979;
      44272:data<=16'd4026;
      44273:data<=16'd3583;
      44274:data<=16'd2861;
      44275:data<=16'd2701;
      44276:data<=16'd2184;
      44277:data<=16'd2270;
      44278:data<=16'd2340;
      44279:data<=16'd1313;
      44280:data<=16'd1506;
      44281:data<=16'd1466;
      44282:data<=16'd582;
      44283:data<=16'd1021;
      44284:data<=16'd502;
      44285:data<=-16'd114;
      44286:data<=16'd435;
      44287:data<=-16'd268;
      44288:data<=-16'd249;
      44289:data<=-16'd690;
      44290:data<=-16'd1982;
      44291:data<=-16'd591;
      44292:data<=-16'd4821;
      44293:data<=-16'd15083;
      44294:data<=-16'd17776;
      44295:data<=-16'd16167;
      44296:data<=-16'd16738;
      44297:data<=-16'd15702;
      44298:data<=-16'd15224;
      44299:data<=-16'd15531;
      44300:data<=-16'd14539;
      44301:data<=-16'd14575;
      44302:data<=-16'd14237;
      44303:data<=-16'd14211;
      44304:data<=-16'd15571;
      44305:data<=-16'd14701;
      44306:data<=-16'd13640;
      44307:data<=-16'd13943;
      44308:data<=-16'd13294;
      44309:data<=-16'd13057;
      44310:data<=-16'd12563;
      44311:data<=-16'd11301;
      44312:data<=-16'd11315;
      44313:data<=-16'd11256;
      44314:data<=-16'd10869;
      44315:data<=-16'd10739;
      44316:data<=-16'd10414;
      44317:data<=-16'd11113;
      44318:data<=-16'd11600;
      44319:data<=-16'd10804;
      44320:data<=-16'd10266;
      44321:data<=-16'd9937;
      44322:data<=-16'd10076;
      44323:data<=-16'd10079;
      44324:data<=-16'd9086;
      44325:data<=-16'd8724;
      44326:data<=-16'd8619;
      44327:data<=-16'd8445;
      44328:data<=-16'd8780;
      44329:data<=-16'd8887;
      44330:data<=-16'd9744;
      44331:data<=-16'd10091;
      44332:data<=-16'd8987;
      44333:data<=-16'd9235;
      44334:data<=-16'd9000;
      44335:data<=-16'd7824;
      44336:data<=-16'd8111;
      44337:data<=-16'd7647;
      44338:data<=-16'd7330;
      44339:data<=-16'd6907;
      44340:data<=-16'd5160;
      44341:data<=-16'd7121;
      44342:data<=-16'd6132;
      44343:data<=16'd3351;
      44344:data<=16'd7203;
      44345:data<=16'd4645;
      44346:data<=16'd5767;
      44347:data<=16'd6220;
      44348:data<=16'd5313;
      44349:data<=16'd6182;
      44350:data<=16'd5564;
      44351:data<=16'd4881;
      44352:data<=16'd5251;
      44353:data<=16'd4593;
      44354:data<=16'd3747;
      44355:data<=16'd2552;
      44356:data<=16'd1428;
      44357:data<=16'd1327;
      44358:data<=16'd1381;
      44359:data<=16'd1718;
      44360:data<=16'd1550;
      44361:data<=16'd937;
      44362:data<=16'd1084;
      44363:data<=16'd931;
      44364:data<=16'd1377;
      44365:data<=16'd2347;
      44366:data<=16'd942;
      44367:data<=-16'd966;
      44368:data<=-16'd1039;
      44369:data<=-16'd789;
      44370:data<=-16'd837;
      44371:data<=-16'd785;
      44372:data<=-16'd344;
      44373:data<=-16'd2;
      44374:data<=-16'd384;
      44375:data<=-16'd839;
      44376:data<=-16'd796;
      44377:data<=-16'd30;
      44378:data<=-16'd161;
      44379:data<=-16'd2047;
      44380:data<=-16'd2804;
      44381:data<=-16'd2582;
      44382:data<=-16'd2564;
      44383:data<=-16'd1600;
      44384:data<=-16'd1723;
      44385:data<=-16'd2564;
      44386:data<=-16'd1992;
      44387:data<=-16'd2009;
      44388:data<=-16'd2164;
      44389:data<=-16'd2446;
      44390:data<=-16'd2813;
      44391:data<=-16'd1181;
      44392:data<=-16'd4623;
      44393:data<=-16'd14135;
      44394:data<=-16'd17490;
      44395:data<=-16'd15838;
      44396:data<=-16'd15711;
      44397:data<=-16'd14598;
      44398:data<=-16'd14008;
      44399:data<=-16'd14431;
      44400:data<=-16'd13092;
      44401:data<=-16'd11972;
      44402:data<=-16'd11367;
      44403:data<=-16'd11053;
      44404:data<=-16'd11926;
      44405:data<=-16'd11890;
      44406:data<=-16'd10836;
      44407:data<=-16'd9950;
      44408:data<=-16'd8865;
      44409:data<=-16'd7685;
      44410:data<=-16'd6613;
      44411:data<=-16'd6272;
      44412:data<=-16'd5868;
      44413:data<=-16'd5028;
      44414:data<=-16'd5328;
      44415:data<=-16'd5030;
      44416:data<=-16'd4444;
      44417:data<=-16'd5858;
      44418:data<=-16'd5850;
      44419:data<=-16'd4548;
      44420:data<=-16'd4814;
      44421:data<=-16'd4447;
      44422:data<=-16'd3876;
      44423:data<=-16'd3882;
      44424:data<=-16'd2992;
      44425:data<=-16'd2593;
      44426:data<=-16'd2272;
      44427:data<=-16'd1527;
      44428:data<=-16'd1944;
      44429:data<=-16'd2610;
      44430:data<=-16'd3221;
      44431:data<=-16'd3395;
      44432:data<=-16'd2611;
      44433:data<=-16'd2678;
      44434:data<=-16'd2500;
      44435:data<=-16'd1512;
      44436:data<=-16'd1428;
      44437:data<=-16'd1036;
      44438:data<=-16'd496;
      44439:data<=16'd117;
      44440:data<=16'd796;
      44441:data<=-16'd1277;
      44442:data<=-16'd1033;
      44443:data<=16'd5682;
      44444:data<=16'd9917;
      44445:data<=16'd8990;
      44446:data<=16'd8866;
      44447:data<=16'd9188;
      44448:data<=16'd8743;
      44449:data<=16'd8798;
      44450:data<=16'd8887;
      44451:data<=16'd8416;
      44452:data<=16'd7759;
      44453:data<=16'd7539;
      44454:data<=16'd6739;
      44455:data<=16'd5131;
      44456:data<=16'd4843;
      44457:data<=16'd4984;
      44458:data<=16'd4326;
      44459:data<=16'd4355;
      44460:data<=16'd4487;
      44461:data<=16'd4314;
      44462:data<=16'd4675;
      44463:data<=16'd4723;
      44464:data<=16'd4610;
      44465:data<=16'd4693;
      44466:data<=16'd4194;
      44467:data<=16'd3526;
      44468:data<=16'd3021;
      44469:data<=16'd2761;
      44470:data<=16'd2958;
      44471:data<=16'd3019;
      44472:data<=16'd3075;
      44473:data<=16'd3289;
      44474:data<=16'd3298;
      44475:data<=16'd3457;
      44476:data<=16'd3397;
      44477:data<=16'd2805;
      44478:data<=16'd2610;
      44479:data<=16'd2995;
      44480:data<=16'd3472;
      44481:data<=16'd3486;
      44482:data<=16'd3087;
      44483:data<=16'd3222;
      44484:data<=16'd3515;
      44485:data<=16'd3301;
      44486:data<=16'd3046;
      44487:data<=16'd3002;
      44488:data<=16'd3391;
      44489:data<=16'd3109;
      44490:data<=16'd2118;
      44491:data<=16'd3574;
      44492:data<=16'd4482;
      44493:data<=-16'd610;
      44494:data<=-16'd5855;
      44495:data<=-16'd5785;
      44496:data<=-16'd4887;
      44497:data<=-16'd5002;
      44498:data<=-16'd4669;
      44499:data<=-16'd4613;
      44500:data<=-16'd4238;
      44501:data<=-16'd3374;
      44502:data<=-16'd3260;
      44503:data<=-16'd3272;
      44504:data<=-16'd2384;
      44505:data<=-16'd940;
      44506:data<=-16'd221;
      44507:data<=-16'd305;
      44508:data<=16'd61;
      44509:data<=16'd387;
      44510:data<=16'd378;
      44511:data<=16'd813;
      44512:data<=16'd1069;
      44513:data<=16'd1110;
      44514:data<=16'd958;
      44515:data<=16'd249;
      44516:data<=16'd546;
      44517:data<=16'd2011;
      44518:data<=16'd3096;
      44519:data<=16'd3253;
      44520:data<=16'd2604;
      44521:data<=16'd2952;
      44522:data<=16'd4052;
      44523:data<=16'd3521;
      44524:data<=16'd2958;
      44525:data<=16'd3300;
      44526:data<=16'd3290;
      44527:data<=16'd3383;
      44528:data<=16'd2980;
      44529:data<=16'd3207;
      44530:data<=16'd4990;
      44531:data<=16'd5059;
      44532:data<=16'd4513;
      44533:data<=16'd5081;
      44534:data<=16'd4440;
      44535:data<=16'd4293;
      44536:data<=16'd4924;
      44537:data<=16'd4065;
      44538:data<=16'd3651;
      44539:data<=16'd3983;
      44540:data<=16'd4243;
      44541:data<=16'd4516;
      44542:data<=16'd5357;
      44543:data<=16'd10578;
      44544:data<=16'd16698;
      44545:data<=16'd16736;
      44546:data<=16'd15343;
      44547:data<=16'd15470;
      44548:data<=16'd14528;
      44549:data<=16'd14210;
      44550:data<=16'd13813;
      44551:data<=16'd13106;
      44552:data<=16'd13406;
      44553:data<=16'd12066;
      44554:data<=16'd11580;
      44555:data<=16'd13796;
      44556:data<=16'd13555;
      44557:data<=16'd11988;
      44558:data<=16'd11846;
      44559:data<=16'd11166;
      44560:data<=16'd10557;
      44561:data<=16'd10002;
      44562:data<=16'd9033;
      44563:data<=16'd9309;
      44564:data<=16'd9545;
      44565:data<=16'd8611;
      44566:data<=16'd8299;
      44567:data<=16'd9050;
      44568:data<=16'd9453;
      44569:data<=16'd8727;
      44570:data<=16'd8099;
      44571:data<=16'd7906;
      44572:data<=16'd7036;
      44573:data<=16'd6438;
      44574:data<=16'd6654;
      44575:data<=16'd6448;
      44576:data<=16'd5689;
      44577:data<=16'd4986;
      44578:data<=16'd4993;
      44579:data<=16'd5583;
      44580:data<=16'd6419;
      44581:data<=16'd7450;
      44582:data<=16'd7336;
      44583:data<=16'd6391;
      44584:data<=16'd6011;
      44585:data<=16'd5565;
      44586:data<=16'd5500;
      44587:data<=16'd5476;
      44588:data<=16'd4857;
      44589:data<=16'd5031;
      44590:data<=16'd4009;
      44591:data<=16'd2886;
      44592:data<=16'd4993;
      44593:data<=16'd3001;
      44594:data<=-16'd4341;
      44595:data<=-16'd6417;
      44596:data<=-16'd4726;
      44597:data<=-16'd5468;
      44598:data<=-16'd6008;
      44599:data<=-16'd5736;
      44600:data<=-16'd5817;
      44601:data<=-16'd5918;
      44602:data<=-16'd6479;
      44603:data<=-16'd6319;
      44604:data<=-16'd5300;
      44605:data<=-16'd4319;
      44606:data<=-16'd2996;
      44607:data<=-16'd2306;
      44608:data<=-16'd2458;
      44609:data<=-16'd2870;
      44610:data<=-16'd3818;
      44611:data<=-16'd3668;
      44612:data<=-16'd2334;
      44613:data<=-16'd2440;
      44614:data<=-16'd3676;
      44615:data<=-16'd3815;
      44616:data<=-16'd2773;
      44617:data<=-16'd1989;
      44618:data<=-16'd1525;
      44619:data<=-16'd1115;
      44620:data<=-16'd1770;
      44621:data<=-16'd2302;
      44622:data<=-16'd1762;
      44623:data<=-16'd1941;
      44624:data<=-16'd2408;
      44625:data<=-16'd2435;
      44626:data<=-16'd2275;
      44627:data<=-16'd1914;
      44628:data<=-16'd2946;
      44629:data<=-16'd3221;
      44630:data<=-16'd960;
      44631:data<=-16'd493;
      44632:data<=-16'd890;
      44633:data<=-16'd253;
      44634:data<=-16'd1292;
      44635:data<=-16'd1742;
      44636:data<=-16'd1262;
      44637:data<=-16'd1673;
      44638:data<=-16'd1178;
      44639:data<=-16'd1850;
      44640:data<=-16'd2234;
      44641:data<=-16'd475;
      44642:data<=-16'd1037;
      44643:data<=16'd2199;
      44644:data<=16'd10372;
      44645:data<=16'd11262;
      44646:data<=16'd8907;
      44647:data<=16'd9382;
      44648:data<=16'd7908;
      44649:data<=16'd7567;
      44650:data<=16'd8278;
      44651:data<=16'd7230;
      44652:data<=16'd8009;
      44653:data<=16'd7645;
      44654:data<=16'd6011;
      44655:data<=16'd7177;
      44656:data<=16'd7216;
      44657:data<=16'd6501;
      44658:data<=16'd6889;
      44659:data<=16'd5688;
      44660:data<=16'd5162;
      44661:data<=16'd5454;
      44662:data<=16'd4589;
      44663:data<=16'd4454;
      44664:data<=16'd4408;
      44665:data<=16'd4115;
      44666:data<=16'd4370;
      44667:data<=16'd4297;
      44668:data<=16'd4319;
      44669:data<=16'd4076;
      44670:data<=16'd3748;
      44671:data<=16'd3742;
      44672:data<=16'd2581;
      44673:data<=16'd1718;
      44674:data<=16'd1701;
      44675:data<=16'd1084;
      44676:data<=16'd708;
      44677:data<=16'd96;
      44678:data<=-16'd77;
      44679:data<=16'd883;
      44680:data<=16'd870;
      44681:data<=16'd787;
      44682:data<=16'd337;
      44683:data<=-16'd775;
      44684:data<=-16'd185;
      44685:data<=-16'd619;
      44686:data<=-16'd1609;
      44687:data<=-16'd669;
      44688:data<=-16'd1309;
      44689:data<=-16'd1506;
      44690:data<=-16'd816;
      44691:data<=-16'd2220;
      44692:data<=-16'd1607;
      44693:data<=-16'd3994;
      44694:data<=-16'd12754;
      44695:data<=-16'd15578;
      44696:data<=-16'd13441;
      44697:data<=-16'd14076;
      44698:data<=-16'd13931;
      44699:data<=-16'd13832;
      44700:data<=-16'd14736;
      44701:data<=-16'd14104;
      44702:data<=-16'd13653;
      44703:data<=-16'd12922;
      44704:data<=-16'd12536;
      44705:data<=-16'd13806;
      44706:data<=-16'd13650;
      44707:data<=-16'd12985;
      44708:data<=-16'd13273;
      44709:data<=-16'd12977;
      44710:data<=-16'd12695;
      44711:data<=-16'd11897;
      44712:data<=-16'd10916;
      44713:data<=-16'd11386;
      44714:data<=-16'd11953;
      44715:data<=-16'd11703;
      44716:data<=-16'd10668;
      44717:data<=-16'd10387;
      44718:data<=-16'd11694;
      44719:data<=-16'd11467;
      44720:data<=-16'd11163;
      44721:data<=-16'd12472;
      44722:data<=-16'd11165;
      44723:data<=-16'd9157;
      44724:data<=-16'd9723;
      44725:data<=-16'd9932;
      44726:data<=-16'd9597;
      44727:data<=-16'd9257;
      44728:data<=-16'd8558;
      44729:data<=-16'd8965;
      44730:data<=-16'd9565;
      44731:data<=-16'd9867;
      44732:data<=-16'd10561;
      44733:data<=-16'd10383;
      44734:data<=-16'd9570;
      44735:data<=-16'd9088;
      44736:data<=-16'd8937;
      44737:data<=-16'd8625;
      44738:data<=-16'd7700;
      44739:data<=-16'd7706;
      44740:data<=-16'd7536;
      44741:data<=-16'd6173;
      44742:data<=-16'd7166;
      44743:data<=-16'd6663;
      44744:data<=-16'd678;
      44745:data<=16'd2601;
      44746:data<=16'd1832;
      44747:data<=16'd2736;
      44748:data<=16'd2820;
      44749:data<=16'd2202;
      44750:data<=16'd3347;
      44751:data<=16'd3130;
      44752:data<=16'd2676;
      44753:data<=16'd3580;
      44754:data<=16'd2253;
      44755:data<=-16'd387;
      44756:data<=-16'd1647;
      44757:data<=-16'd1958;
      44758:data<=-16'd1002;
      44759:data<=-16'd205;
      44760:data<=-16'd878;
      44761:data<=-16'd678;
      44762:data<=16'd94;
      44763:data<=-16'd397;
      44764:data<=-16'd482;
      44765:data<=16'd355;
      44766:data<=16'd485;
      44767:data<=-16'd537;
      44768:data<=-16'd2099;
      44769:data<=-16'd2520;
      44770:data<=-16'd1903;
      44771:data<=-16'd2231;
      44772:data<=-16'd2385;
      44773:data<=-16'd1685;
      44774:data<=-16'd1639;
      44775:data<=-16'd989;
      44776:data<=-16'd24;
      44777:data<=-16'd775;
      44778:data<=-16'd1221;
      44779:data<=-16'd1107;
      44780:data<=-16'd2343;
      44781:data<=-16'd3011;
      44782:data<=-16'd1980;
      44783:data<=-16'd926;
      44784:data<=-16'd823;
      44785:data<=-16'd769;
      44786:data<=16'd293;
      44787:data<=16'd70;
      44788:data<=-16'd1246;
      44789:data<=-16'd226;
      44790:data<=16'd256;
      44791:data<=-16'd711;
      44792:data<=-16'd296;
      44793:data<=-16'd3650;
      44794:data<=-16'd10543;
      44795:data<=-16'd12707;
      44796:data<=-16'd11881;
      44797:data<=-16'd11744;
      44798:data<=-16'd10947;
      44799:data<=-16'd10363;
      44800:data<=-16'd9970;
      44801:data<=-16'd9905;
      44802:data<=-16'd10399;
      44803:data<=-16'd9277;
      44804:data<=-16'd8229;
      44805:data<=-16'd8514;
      44806:data<=-16'd8191;
      44807:data<=-16'd8348;
      44808:data<=-16'd8440;
      44809:data<=-16'd7228;
      44810:data<=-16'd6601;
      44811:data<=-16'd6273;
      44812:data<=-16'd5996;
      44813:data<=-16'd6122;
      44814:data<=-16'd5477;
      44815:data<=-16'd4745;
      44816:data<=-16'd4152;
      44817:data<=-16'd4041;
      44818:data<=-16'd5098;
      44819:data<=-16'd4493;
      44820:data<=-16'd3016;
      44821:data<=-16'd3606;
      44822:data<=-16'd3621;
      44823:data<=-16'd2416;
      44824:data<=-16'd1930;
      44825:data<=-16'd1967;
      44826:data<=-16'd2658;
      44827:data<=-16'd2864;
      44828:data<=-16'd2099;
      44829:data<=-16'd1821;
      44830:data<=-16'd1764;
      44831:data<=-16'd2276;
      44832:data<=-16'd2905;
      44833:data<=-16'd2308;
      44834:data<=-16'd2056;
      44835:data<=-16'd1795;
      44836:data<=-16'd854;
      44837:data<=-16'd908;
      44838:data<=-16'd884;
      44839:data<=-16'd698;
      44840:data<=-16'd1142;
      44841:data<=-16'd1413;
      44842:data<=-16'd2990;
      44843:data<=-16'd2372;
      44844:data<=16'd4407;
      44845:data<=16'd9245;
      44846:data<=16'd8296;
      44847:data<=16'd7982;
      44848:data<=16'd8913;
      44849:data<=16'd9051;
      44850:data<=16'd9270;
      44851:data<=16'd9397;
      44852:data<=16'd9221;
      44853:data<=16'd8745;
      44854:data<=16'd8692;
      44855:data<=16'd8360;
      44856:data<=16'd5729;
      44857:data<=16'd4517;
      44858:data<=16'd6103;
      44859:data<=16'd5773;
      44860:data<=16'd5286;
      44861:data<=16'd5990;
      44862:data<=16'd4977;
      44863:data<=16'd4998;
      44864:data<=16'd6038;
      44865:data<=16'd5688;
      44866:data<=16'd5927;
      44867:data<=16'd4758;
      44868:data<=16'd2880;
      44869:data<=16'd3965;
      44870:data<=16'd3770;
      44871:data<=16'd2463;
      44872:data<=16'd3492;
      44873:data<=16'd3732;
      44874:data<=16'd3268;
      44875:data<=16'd2734;
      44876:data<=16'd2209;
      44877:data<=16'd3996;
      44878:data<=16'd4179;
      44879:data<=16'd2943;
      44880:data<=16'd4387;
      44881:data<=16'd4288;
      44882:data<=16'd3803;
      44883:data<=16'd5225;
      44884:data<=16'd4193;
      44885:data<=16'd3771;
      44886:data<=16'd4736;
      44887:data<=16'd3231;
      44888:data<=16'd2740;
      44889:data<=16'd3991;
      44890:data<=16'd4946;
      44891:data<=16'd5165;
      44892:data<=16'd4454;
      44893:data<=16'd4726;
      44894:data<=16'd1629;
      44895:data<=-16'd4942;
      44896:data<=-16'd5741;
      44897:data<=-16'd4258;
      44898:data<=-16'd5042;
      44899:data<=-16'd4664;
      44900:data<=-16'd5181;
      44901:data<=-16'd4901;
      44902:data<=-16'd3456;
      44903:data<=-16'd4705;
      44904:data<=-16'd4091;
      44905:data<=-16'd2005;
      44906:data<=-16'd1098;
      44907:data<=16'd817;
      44908:data<=16'd555;
      44909:data<=16'd494;
      44910:data<=16'd2106;
      44911:data<=16'd74;
      44912:data<=-16'd563;
      44913:data<=16'd966;
      44914:data<=16'd411;
      44915:data<=16'd999;
      44916:data<=16'd146;
      44917:data<=-16'd429;
      44918:data<=16'd3068;
      44919:data<=16'd3535;
      44920:data<=16'd3559;
      44921:data<=16'd5435;
      44922:data<=16'd3092;
      44923:data<=16'd2191;
      44924:data<=16'd4347;
      44925:data<=16'd4137;
      44926:data<=16'd3991;
      44927:data<=16'd4196;
      44928:data<=16'd3714;
      44929:data<=16'd2757;
      44930:data<=16'd2118;
      44931:data<=16'd4479;
      44932:data<=16'd5570;
      44933:data<=16'd4074;
      44934:data<=16'd4273;
      44935:data<=16'd3938;
      44936:data<=16'd4264;
      44937:data<=16'd5635;
      44938:data<=16'd4099;
      44939:data<=16'd3651;
      44940:data<=16'd4737;
      44941:data<=16'd4099;
      44942:data<=16'd3200;
      44943:data<=16'd3274;
      44944:data<=16'd8583;
      44945:data<=16'd15335;
      44946:data<=16'd15242;
      44947:data<=16'd14898;
      44948:data<=16'd15699;
      44949:data<=16'd13162;
      44950:data<=16'd12912;
      44951:data<=16'd13540;
      44952:data<=16'd11934;
      44953:data<=16'd12067;
      44954:data<=16'd12601;
      44955:data<=16'd13006;
      44956:data<=16'd13517;
      44957:data<=16'd12386;
      44958:data<=16'd12000;
      44959:data<=16'd11230;
      44960:data<=16'd8854;
      44961:data<=16'd9163;
      44962:data<=16'd11188;
      44963:data<=16'd11345;
      44964:data<=16'd10956;
      44965:data<=16'd11330;
      44966:data<=16'd10681;
      44967:data<=16'd9407;
      44968:data<=16'd9662;
      44969:data<=16'd9081;
      44970:data<=16'd8031;
      44971:data<=16'd9051;
      44972:data<=16'd8580;
      44973:data<=16'd7460;
      44974:data<=16'd7598;
      44975:data<=16'd6296;
      44976:data<=16'd6484;
      44977:data<=16'd7065;
      44978:data<=16'd4864;
      44979:data<=16'd4519;
      44980:data<=16'd5460;
      44981:data<=16'd6519;
      44982:data<=16'd8055;
      44983:data<=16'd7203;
      44984:data<=16'd7840;
      44985:data<=16'd8457;
      44986:data<=16'd5507;
      44987:data<=16'd6064;
      44988:data<=16'd6698;
      44989:data<=16'd4428;
      44990:data<=16'd5711;
      44991:data<=16'd5594;
      44992:data<=16'd4707;
      44993:data<=16'd7221;
      44994:data<=16'd4168;
      44995:data<=-16'd2487;
      44996:data<=-16'd4361;
      44997:data<=-16'd4026;
      44998:data<=-16'd4147;
      44999:data<=-16'd4798;
      45000:data<=-16'd4796;
      45001:data<=-16'd4470;
      45002:data<=-16'd4487;
      45003:data<=-16'd3812;
      45004:data<=-16'd5430;
      45005:data<=-16'd5937;
      45006:data<=-16'd2531;
      45007:data<=-16'd3086;
      45008:data<=-16'd4046;
      45009:data<=-16'd2303;
      45010:data<=-16'd3832;
      45011:data<=-16'd3744;
      45012:data<=-16'd2763;
      45013:data<=-16'd4077;
      45014:data<=-16'd2670;
      45015:data<=-16'd3209;
      45016:data<=-16'd4411;
      45017:data<=-16'd2114;
      45018:data<=-16'd2740;
      45019:data<=-16'd1798;
      45020:data<=16'd55;
      45021:data<=-16'd3385;
      45022:data<=-16'd2990;
      45023:data<=-16'd1154;
      45024:data<=-16'd2743;
      45025:data<=-16'd967;
      45026:data<=-16'd802;
      45027:data<=-16'd2267;
      45028:data<=-16'd224;
      45029:data<=-16'd1004;
      45030:data<=-16'd2359;
      45031:data<=-16'd673;
      45032:data<=-16'd634;
      45033:data<=-16'd1906;
      45034:data<=-16'd2384;
      45035:data<=-16'd399;
      45036:data<=16'd949;
      45037:data<=-16'd1152;
      45038:data<=-16'd414;
      45039:data<=16'd159;
      45040:data<=-16'd2746;
      45041:data<=-16'd749;
      45042:data<=16'd1218;
      45043:data<=-16'd2017;
      45044:data<=16'd708;
      45045:data<=16'd9420;
      45046:data<=16'd12519;
      45047:data<=16'd9846;
      45048:data<=16'd9467;
      45049:data<=16'd11079;
      45050:data<=16'd9226;
      45051:data<=16'd6971;
      45052:data<=16'd7700;
      45053:data<=16'd8185;
      45054:data<=16'd7186;
      45055:data<=16'd6320;
      45056:data<=16'd7051;
      45057:data<=16'd7928;
      45058:data<=16'd7815;
      45059:data<=16'd8137;
      45060:data<=16'd7012;
      45061:data<=16'd6044;
      45062:data<=16'd6874;
      45063:data<=16'd4983;
      45064:data<=16'd4272;
      45065:data<=16'd5735;
      45066:data<=16'd3400;
      45067:data<=16'd3008;
      45068:data<=16'd5002;
      45069:data<=16'd3915;
      45070:data<=16'd3283;
      45071:data<=16'd2432;
      45072:data<=16'd1767;
      45073:data<=16'd2270;
      45074:data<=-16'd156;
      45075:data<=-16'd781;
      45076:data<=16'd177;
      45077:data<=-16'd1604;
      45078:data<=-16'd707;
      45079:data<=16'd264;
      45080:data<=-16'd576;
      45081:data<=16'd881;
      45082:data<=16'd842;
      45083:data<=-16'd221;
      45084:data<=-16'd2300;
      45085:data<=-16'd5645;
      45086:data<=-16'd3946;
      45087:data<=-16'd2710;
      45088:data<=-16'd3882;
      45089:data<=-16'd2541;
      45090:data<=-16'd5059;
      45091:data<=-16'd6893;
      45092:data<=-16'd3494;
      45093:data<=-16'd4162;
      45094:data<=-16'd8337;
      45095:data<=-16'd14862;
      45096:data<=-16'd19443;
      45097:data<=-16'd15907;
      45098:data<=-16'd17697;
      45099:data<=-16'd24924;
      45100:data<=-16'd24667;
      45101:data<=-16'd23892;
      45102:data<=-16'd24535;
      45103:data<=-16'd22398;
      45104:data<=-16'd21695;
      45105:data<=-16'd21889;
      45106:data<=-16'd22400;
      45107:data<=-16'd21570;
      45108:data<=-16'd18698;
      45109:data<=-16'd21191;
      45110:data<=-16'd25913;
      45111:data<=-16'd23234;
      45112:data<=-16'd15870;
      45113:data<=-16'd13082;
      45114:data<=-16'd15725;
      45115:data<=-16'd14722;
      45116:data<=-16'd12704;
      45117:data<=-16'd15740;
      45118:data<=-16'd13894;
      45119:data<=-16'd8125;
      45120:data<=-16'd8099;
      45121:data<=-16'd10602;
      45122:data<=-16'd12471;
      45123:data<=-16'd11779;
      45124:data<=-16'd10383;
      45125:data<=-16'd10975;
      45126:data<=-16'd8156;
      45127:data<=-16'd6417;
      45128:data<=-16'd7191;
      45129:data<=-16'd5539;
      45130:data<=-16'd9172;
      45131:data<=-16'd6015;
      45132:data<=16'd9841;
      45133:data<=16'd5694;
      45134:data<=-16'd13188;
      45135:data<=-16'd15370;
      45136:data<=-16'd10085;
      45137:data<=-16'd4957;
      45138:data<=16'd1204;
      45139:data<=-16'd4784;
      45140:data<=-16'd12011;
      45141:data<=-16'd402;
      45142:data<=16'd15658;
      45143:data<=16'd17617;
      45144:data<=16'd11194;
      45145:data<=16'd6752;
      45146:data<=16'd8163;
      45147:data<=16'd12869;
      45148:data<=16'd12734;
      45149:data<=16'd9602;
      45150:data<=16'd9430;
      45151:data<=16'd9406;
      45152:data<=16'd11803;
      45153:data<=16'd11835;
      45154:data<=16'd162;
      45155:data<=-16'd5815;
      45156:data<=16'd2108;
      45157:data<=16'd5594;
      45158:data<=16'd2561;
      45159:data<=-16'd854;
      45160:data<=-16'd4326;
      45161:data<=-16'd4522;
      45162:data<=-16'd1462;
      45163:data<=16'd1438;
      45164:data<=-16'd3573;
      45165:data<=-16'd11485;
      45166:data<=-16'd7418;
      45167:data<=-16'd3867;
      45168:data<=-16'd5990;
      45169:data<=-16'd2237;
      45170:data<=-16'd6948;
      45171:data<=-16'd12834;
      45172:data<=-16'd1574;
      45173:data<=-16'd2156;
      45174:data<=-16'd16393;
      45175:data<=-16'd13013;
      45176:data<=-16'd7175;
      45177:data<=-16'd13515;
      45178:data<=-16'd14392;
      45179:data<=-16'd11615;
      45180:data<=-16'd12628;
      45181:data<=-16'd8887;
      45182:data<=-16'd7991;
      45183:data<=-16'd18948;
      45184:data<=-16'd23725;
      45185:data<=-16'd18700;
      45186:data<=-16'd19973;
      45187:data<=-16'd22660;
      45188:data<=-16'd22262;
      45189:data<=-16'd24726;
      45190:data<=-16'd25945;
      45191:data<=-16'd23240;
      45192:data<=-16'd16659;
      45193:data<=-16'd14991;
      45194:data<=-16'd24024;
      45195:data<=-16'd23217;
      45196:data<=-16'd15787;
      45197:data<=-16'd21094;
      45198:data<=-16'd22900;
      45199:data<=-16'd17807;
      45200:data<=-16'd16233;
      45201:data<=-16'd11412;
      45202:data<=-16'd9150;
      45203:data<=-16'd11194;
      45204:data<=-16'd12337;
      45205:data<=-16'd13467;
      45206:data<=-16'd7274;
      45207:data<=-16'd5227;
      45208:data<=-16'd10865;
      45209:data<=-16'd6100;
      45210:data<=-16'd6617;
      45211:data<=-16'd9646;
      45212:data<=16'd6099;
      45213:data<=16'd10003;
      45214:data<=-16'd3509;
      45215:data<=-16'd4294;
      45216:data<=-16'd808;
      45217:data<=16'd165;
      45218:data<=16'd5216;
      45219:data<=16'd4135;
      45220:data<=-16'd5921;
      45221:data<=-16'd9545;
      45222:data<=-16'd1189;
      45223:data<=16'd6;
      45224:data<=-16'd2362;
      45225:data<=16'd11829;
      45226:data<=16'd19516;
      45227:data<=16'd15814;
      45228:data<=16'd24498;
      45229:data<=16'd26837;
      45230:data<=16'd19952;
      45231:data<=16'd23875;
      45232:data<=16'd26585;
      45233:data<=16'd26063;
      45234:data<=16'd26326;
      45235:data<=16'd22312;
      45236:data<=16'd20742;
      45237:data<=16'd20316;
      45238:data<=16'd22125;
      45239:data<=16'd23352;
      45240:data<=16'd12301;
      45241:data<=16'd8505;
      45242:data<=16'd17855;
      45243:data<=16'd19872;
      45244:data<=16'd19032;
      45245:data<=16'd16785;
      45246:data<=16'd13982;
      45247:data<=16'd18675;
      45248:data<=16'd19828;
      45249:data<=16'd18483;
      45250:data<=16'd17249;
      45251:data<=16'd13565;
      45252:data<=16'd21452;
      45253:data<=16'd24579;
      45254:data<=16'd12336;
      45255:data<=16'd13876;
      45256:data<=16'd19584;
      45257:data<=16'd13967;
      45258:data<=16'd13982;
      45259:data<=16'd14860;
      45260:data<=16'd11065;
      45261:data<=16'd8202;
      45262:data<=16'd4751;
      45263:data<=16'd5612;
      45264:data<=16'd7081;
      45265:data<=16'd5964;
      45266:data<=16'd7659;
      45267:data<=16'd2682;
      45268:data<=-16'd8022;
      45269:data<=-16'd10916;
      45270:data<=-16'd8445;
      45271:data<=-16'd6960;
      45272:data<=-16'd9491;
      45273:data<=-16'd12419;
      45274:data<=-16'd8308;
      45275:data<=-16'd2995;
      45276:data<=-16'd4654;
      45277:data<=-16'd7550;
      45278:data<=-16'd2490;
      45279:data<=-16'd635;
      45280:data<=-16'd10727;
      45281:data<=-16'd9197;
      45282:data<=16'd723;
      45283:data<=-16'd4893;
      45284:data<=-16'd4423;
      45285:data<=16'd6413;
      45286:data<=16'd5046;
      45287:data<=16'd4027;
      45288:data<=16'd4884;
      45289:data<=16'd140;
      45290:data<=16'd1060;
      45291:data<=16'd1612;
      45292:data<=16'd1892;
      45293:data<=16'd5254;
      45294:data<=-16'd1080;
      45295:data<=-16'd6605;
      45296:data<=-16'd2472;
      45297:data<=16'd2241;
      45298:data<=16'd5009;
      45299:data<=16'd1565;
      45300:data<=16'd2247;
      45301:data<=16'd8175;
      45302:data<=16'd2917;
      45303:data<=16'd5407;
      45304:data<=16'd14231;
      45305:data<=16'd4331;
      45306:data<=-16'd613;
      45307:data<=16'd2475;
      45308:data<=-16'd943;
      45309:data<=16'd11793;
      45310:data<=16'd25775;
      45311:data<=16'd21604;
      45312:data<=16'd26080;
      45313:data<=16'd32761;
      45314:data<=16'd26233;
      45315:data<=16'd25629;
      45316:data<=16'd31616;
      45317:data<=16'd31492;
      45318:data<=16'd29543;
      45319:data<=16'd30970;
      45320:data<=16'd28746;
      45321:data<=16'd22204;
      45322:data<=16'd24513;
      45323:data<=16'd27372;
      45324:data<=16'd20521;
      45325:data<=16'd21585;
      45326:data<=16'd23484;
      45327:data<=16'd13054;
      45328:data<=16'd13847;
      45329:data<=16'd23758;
      45330:data<=16'd19572;
      45331:data<=16'd12490;
      45332:data<=16'd15515;
      45333:data<=16'd18553;
      45334:data<=16'd11514;
      45335:data<=16'd4502;
      45336:data<=16'd10683;
      45337:data<=16'd12593;
      45338:data<=16'd1447;
      45339:data<=16'd974;
      45340:data<=16'd9756;
      45341:data<=16'd8479;
      45342:data<=16'd1283;
      45343:data<=-16'd916;
      45344:data<=16'd4896;
      45345:data<=16'd6721;
      45346:data<=-16'd3594;
      45347:data<=-16'd7914;
      45348:data<=-16'd5269;
      45349:data<=-16'd8235;
      45350:data<=-16'd4739;
      45351:data<=-16'd2473;
      45352:data<=-16'd17690;
      45353:data<=-16'd26488;
      45354:data<=-16'd21105;
      45355:data<=-16'd20983;
      45356:data<=-16'd23554;
      45357:data<=-16'd24685;
      45358:data<=-16'd25787;
      45359:data<=-16'd22532;
      45360:data<=-16'd20491;
      45361:data<=-16'd22093;
      45362:data<=-16'd24665;
      45363:data<=-16'd29654;
      45364:data<=-16'd29122;
      45365:data<=-16'd22973;
      45366:data<=-16'd22974;
      45367:data<=-16'd26376;
      45368:data<=-16'd27442;
      45369:data<=-16'd27108;
      45370:data<=-16'd25150;
      45371:data<=-16'd23681;
      45372:data<=-16'd23355;
      45373:data<=-16'd23790;
      45374:data<=-16'd24967;
      45375:data<=-16'd23871;
      45376:data<=-16'd20930;
      45377:data<=-16'd19259;
      45378:data<=-16'd20760;
      45379:data<=-16'd21601;
      45380:data<=-16'd18477;
      45381:data<=-16'd21823;
      45382:data<=-16'd25924;
      45383:data<=-16'd16007;
      45384:data<=-16'd12960;
      45385:data<=-16'd21993;
      45386:data<=-16'd19623;
      45387:data<=-16'd15967;
      45388:data<=-16'd18448;
      45389:data<=-16'd15300;
      45390:data<=-16'd13323;
      45391:data<=-16'd12625;
      45392:data<=-16'd12231;
      45393:data<=-16'd13599;
      45394:data<=-16'd1997;
      45395:data<=16'd8032;
      45396:data<=16'd462;
      45397:data<=16'd133;
      45398:data<=16'd5177;
      45399:data<=16'd21;
      45400:data<=-16'd634;
      45401:data<=16'd4064;
      45402:data<=16'd6232;
      45403:data<=16'd7436;
      45404:data<=16'd3664;
      45405:data<=-16'd802;
      45406:data<=-16'd214;
      45407:data<=16'd1083;
      45408:data<=16'd343;
      45409:data<=-16'd1010;
      45410:data<=16'd1368;
      45411:data<=16'd2334;
      45412:data<=16'd1172;
      45413:data<=16'd9388;
      45414:data<=16'd12094;
      45415:data<=16'd2917;
      45416:data<=16'd5530;
      45417:data<=16'd9317;
      45418:data<=16'd3098;
      45419:data<=16'd3606;
      45420:data<=16'd3827;
      45421:data<=16'd1535;
      45422:data<=16'd3394;
      45423:data<=16'd1444;
      45424:data<=16'd4654;
      45425:data<=16'd6705;
      45426:data<=-16'd4356;
      45427:data<=-16'd2246;
      45428:data<=16'd7151;
      45429:data<=16'd2510;
      45430:data<=16'd3366;
      45431:data<=16'd6933;
      45432:data<=16'd3861;
      45433:data<=16'd8592;
      45434:data<=16'd10665;
      45435:data<=16'd732;
      45436:data<=-16'd9016;
      45437:data<=-16'd11097;
      45438:data<=-16'd6205;
      45439:data<=-16'd7790;
      45440:data<=-16'd11336;
      45441:data<=-16'd2736;
      45442:data<=-16'd1345;
      45443:data<=-16'd6987;
      45444:data<=-16'd1882;
      45445:data<=-16'd3741;
      45446:data<=-16'd11794;
      45447:data<=-16'd5924;
      45448:data<=16'd523;
      45449:data<=-16'd3839;
      45450:data<=-16'd7645;
      45451:data<=-16'd3262;
      45452:data<=16'd2710;
      45453:data<=16'd2258;
      45454:data<=16'd1770;
      45455:data<=16'd2889;
      45456:data<=-16'd1259;
      45457:data<=-16'd5912;
      45458:data<=-16'd6536;
      45459:data<=-16'd3362;
      45460:data<=16'd111;
      45461:data<=-16'd2645;
      45462:data<=-16'd6032;
      45463:data<=-16'd6617;
      45464:data<=-16'd7274;
      45465:data<=-16'd3110;
      45466:data<=16'd535;
      45467:data<=-16'd1865;
      45468:data<=-16'd74;
      45469:data<=16'd5216;
      45470:data<=16'd2275;
      45471:data<=-16'd6088;
      45472:data<=-16'd4143;
      45473:data<=16'd5119;
      45474:data<=16'd3730;
      45475:data<=16'd180;
      45476:data<=16'd2834;
      45477:data<=16'd2726;
      45478:data<=16'd9826;
      45479:data<=16'd19866;
      45480:data<=16'd17520;
      45481:data<=16'd19418;
      45482:data<=16'd23156;
      45483:data<=16'd15635;
      45484:data<=16'd15238;
      45485:data<=16'd21352;
      45486:data<=16'd21629;
      45487:data<=16'd20580;
      45488:data<=16'd15261;
      45489:data<=16'd10847;
      45490:data<=16'd15394;
      45491:data<=16'd18791;
      45492:data<=16'd17925;
      45493:data<=16'd17142;
      45494:data<=16'd18116;
      45495:data<=16'd19611;
      45496:data<=16'd14672;
      45497:data<=16'd9379;
      45498:data<=16'd12199;
      45499:data<=16'd13392;
      45500:data<=16'd12061;
      45501:data<=16'd16745;
      45502:data<=16'd21231;
      45503:data<=16'd19790;
      45504:data<=16'd15361;
      45505:data<=16'd9033;
      45506:data<=16'd8608;
      45507:data<=16'd15414;
      45508:data<=16'd12809;
      45509:data<=16'd7285;
      45510:data<=16'd12085;
      45511:data<=16'd9347;
      45512:data<=16'd6270;
      45513:data<=16'd17619;
      45514:data<=16'd18779;
      45515:data<=16'd17133;
      45516:data<=16'd24750;
      45517:data<=16'd16903;
      45518:data<=16'd11634;
      45519:data<=16'd16557;
      45520:data<=16'd1087;
      45521:data<=-16'd9711;
      45522:data<=-16'd2611;
      45523:data<=-16'd4786;
      45524:data<=-16'd5036;
      45525:data<=-16'd1039;
      45526:data<=-16'd4557;
      45527:data<=-16'd5949;
      45528:data<=-16'd7785;
      45529:data<=-16'd6384;
      45530:data<=-16'd385;
      45531:data<=-16'd4996;
      45532:data<=-16'd7386;
      45533:data<=-16'd3004;
      45534:data<=-16'd6996;
      45535:data<=-16'd10006;
      45536:data<=-16'd9752;
      45537:data<=-16'd10611;
      45538:data<=-16'd7282;
      45539:data<=-16'd7523;
      45540:data<=-16'd9471;
      45541:data<=-16'd5703;
      45542:data<=-16'd6540;
      45543:data<=-16'd12052;
      45544:data<=-16'd13250;
      45545:data<=-16'd12170;
      45546:data<=-16'd13409;
      45547:data<=-16'd12983;
      45548:data<=-16'd7312;
      45549:data<=-16'd6984;
      45550:data<=-16'd11069;
      45551:data<=-16'd8296;
      45552:data<=-16'd7433;
      45553:data<=-16'd8314;
      45554:data<=-16'd6734;
      45555:data<=-16'd13103;
      45556:data<=-16'd13999;
      45557:data<=-16'd4605;
      45558:data<=-16'd7028;
      45559:data<=-16'd16543;
      45560:data<=-16'd21643;
      45561:data<=-16'd16318;
      45562:data<=16'd1190;
      45563:data<=16'd1811;
      45564:data<=-16'd11590;
      45565:data<=-16'd5529;
      45566:data<=16'd1929;
      45567:data<=-16'd2349;
      45568:data<=-16'd832;
      45569:data<=-16'd1083;
      45570:data<=-16'd1897;
      45571:data<=16'd3239;
      45572:data<=-16'd3048;
      45573:data<=-16'd13947;
      45574:data<=-16'd12348;
      45575:data<=-16'd7327;
      45576:data<=-16'd4096;
      45577:data<=-16'd3547;
      45578:data<=-16'd8560;
      45579:data<=-16'd10161;
      45580:data<=-16'd7538;
      45581:data<=-16'd8980;
      45582:data<=-16'd10311;
      45583:data<=-16'd8831;
      45584:data<=-16'd6931;
      45585:data<=-16'd2361;
      45586:data<=-16'd2416;
      45587:data<=-16'd11515;
      45588:data<=-16'd15177;
      45589:data<=-16'd9782;
      45590:data<=-16'd5186;
      45591:data<=-16'd4672;
      45592:data<=-16'd8971;
      45593:data<=-16'd10000;
      45594:data<=-16'd5392;
      45595:data<=-16'd9388;
      45596:data<=-16'd13864;
      45597:data<=-16'd6579;
      45598:data<=-16'd3462;
      45599:data<=-16'd7373;
      45600:data<=-16'd9391;
      45601:data<=-16'd9787;
      45602:data<=-16'd4258;
      45603:data<=-16'd3372;
      45604:data<=-16'd18224;
      45605:data<=-16'd29214;
      45606:data<=-16'd27181;
      45607:data<=-16'd24755;
      45608:data<=-16'd26271;
      45609:data<=-16'd28517;
      45610:data<=-16'd26348;
      45611:data<=-16'd21913;
      45612:data<=-16'd19992;
      45613:data<=-16'd16274;
      45614:data<=-16'd13367;
      45615:data<=-16'd13973;
      45616:data<=-16'd12008;
      45617:data<=-16'd10525;
      45618:data<=-16'd11524;
      45619:data<=-16'd10601;
      45620:data<=-16'd9567;
      45621:data<=-16'd9856;
      45622:data<=-16'd9988;
      45623:data<=-16'd7535;
      45624:data<=-16'd5098;
      45625:data<=-16'd7764;
      45626:data<=-16'd7982;
      45627:data<=-16'd5935;
      45628:data<=-16'd8417;
      45629:data<=-16'd5134;
      45630:data<=-16'd162;
      45631:data<=-16'd3551;
      45632:data<=-16'd3547;
      45633:data<=-16'd1804;
      45634:data<=-16'd613;
      45635:data<=16'd6552;
      45636:data<=16'd5051;
      45637:data<=-16'd450;
      45638:data<=16'd5333;
      45639:data<=16'd5056;
      45640:data<=16'd220;
      45641:data<=16'd4601;
      45642:data<=16'd6822;
      45643:data<=16'd7344;
      45644:data<=16'd8392;
      45645:data<=16'd7498;
      45646:data<=16'd16841;
      45647:data<=16'd26884;
      45648:data<=16'd24838;
      45649:data<=16'd23316;
      45650:data<=16'd21610;
      45651:data<=16'd19731;
      45652:data<=16'd24668;
      45653:data<=16'd23241;
      45654:data<=16'd16625;
      45655:data<=16'd18503;
      45656:data<=16'd22711;
      45657:data<=16'd23933;
      45658:data<=16'd20912;
      45659:data<=16'd15556;
      45660:data<=16'd17713;
      45661:data<=16'd22318;
      45662:data<=16'd19042;
      45663:data<=16'd11453;
      45664:data<=16'd8818;
      45665:data<=16'd14671;
      45666:data<=16'd15576;
      45667:data<=16'd9333;
      45668:data<=16'd12689;
      45669:data<=16'd16198;
      45670:data<=16'd10563;
      45671:data<=16'd10745;
      45672:data<=16'd14035;
      45673:data<=16'd14973;
      45674:data<=16'd16810;
      45675:data<=16'd11802;
      45676:data<=16'd5213;
      45677:data<=16'd7006;
      45678:data<=16'd11009;
      45679:data<=16'd12784;
      45680:data<=16'd9875;
      45681:data<=16'd7228;
      45682:data<=16'd12035;
      45683:data<=16'd13121;
      45684:data<=16'd7762;
      45685:data<=16'd9130;
      45686:data<=16'd14248;
      45687:data<=16'd8530;
      45688:data<=-16'd5277;
      45689:data<=-16'd8924;
      45690:data<=-16'd7830;
      45691:data<=-16'd14380;
      45692:data<=-16'd10950;
      45693:data<=-16'd3137;
      45694:data<=-16'd8887;
      45695:data<=-16'd7368;
      45696:data<=-16'd3609;
      45697:data<=-16'd11674;
      45698:data<=-16'd5856;
      45699:data<=16'd3386;
      45700:data<=-16'd2748;
      45701:data<=-16'd1986;
      45702:data<=16'd2014;
      45703:data<=16'd917;
      45704:data<=16'd2275;
      45705:data<=-16'd4111;
      45706:data<=-16'd6196;
      45707:data<=16'd4855;
      45708:data<=16'd3621;
      45709:data<=-16'd2006;
      45710:data<=16'd1563;
      45711:data<=-16'd481;
      45712:data<=16'd1560;
      45713:data<=16'd10813;
      45714:data<=16'd8813;
      45715:data<=16'd7955;
      45716:data<=16'd14819;
      45717:data<=16'd13298;
      45718:data<=16'd9884;
      45719:data<=16'd9306;
      45720:data<=16'd6369;
      45721:data<=16'd8699;
      45722:data<=16'd10361;
      45723:data<=16'd6091;
      45724:data<=16'd6573;
      45725:data<=16'd5515;
      45726:data<=16'd3498;
      45727:data<=16'd8699;
      45728:data<=16'd8146;
      45729:data<=16'd8945;
      45730:data<=16'd18780;
      45731:data<=16'd18647;
      45732:data<=16'd18848;
      45733:data<=16'd26671;
      45734:data<=16'd23629;
      45735:data<=16'd19996;
      45736:data<=16'd19884;
      45737:data<=16'd14942;
      45738:data<=16'd17126;
      45739:data<=16'd19259;
      45740:data<=16'd15144;
      45741:data<=16'd15823;
      45742:data<=16'd11872;
      45743:data<=16'd4949;
      45744:data<=16'd5870;
      45745:data<=16'd8548;
      45746:data<=16'd14642;
      45747:data<=16'd15274;
      45748:data<=16'd4124;
      45749:data<=16'd2972;
      45750:data<=16'd7418;
      45751:data<=16'd3189;
      45752:data<=16'd2726;
      45753:data<=16'd2135;
      45754:data<=-16'd3174;
      45755:data<=-16'd121;
      45756:data<=16'd3412;
      45757:data<=16'd209;
      45758:data<=-16'd1525;
      45759:data<=-16'd7594;
      45760:data<=-16'd13450;
      45761:data<=-16'd5222;
      45762:data<=-16'd1530;
      45763:data<=-16'd9952;
      45764:data<=-16'd8091;
      45765:data<=-16'd5084;
      45766:data<=-16'd12666;
      45767:data<=-16'd13527;
      45768:data<=-16'd11600;
      45769:data<=-16'd10927;
      45770:data<=-16'd4734;
      45771:data<=-16'd11943;
      45772:data<=-16'd28656;
      45773:data<=-16'd29974;
      45774:data<=-16'd27388;
      45775:data<=-16'd31235;
      45776:data<=-16'd32479;
      45777:data<=-16'd28959;
      45778:data<=-16'd24557;
      45779:data<=-16'd28197;
      45780:data<=-16'd33860;
      45781:data<=-16'd30523;
      45782:data<=-16'd28702;
      45783:data<=-16'd28169;
      45784:data<=-16'd23689;
      45785:data<=-16'd23182;
      45786:data<=-16'd20836;
      45787:data<=-16'd18801;
      45788:data<=-16'd27407;
      45789:data<=-16'd31360;
      45790:data<=-16'd26040;
      45791:data<=-16'd24157;
      45792:data<=-16'd21382;
      45793:data<=-16'd18545;
      45794:data<=-16'd23778;
      45795:data<=-16'd24623;
      45796:data<=-16'd15300;
      45797:data<=-16'd13386;
      45798:data<=-16'd18459;
      45799:data<=-16'd16266;
      45800:data<=-16'd15027;
      45801:data<=-16'd17091;
      45802:data<=-16'd10740;
      45803:data<=-16'd6217;
      45804:data<=-16'd11726;
      45805:data<=-16'd14574;
      45806:data<=-16'd11752;
      45807:data<=-16'd11585;
      45808:data<=-16'd17039;
      45809:data<=-16'd20234;
      45810:data<=-16'd15279;
      45811:data<=-16'd11505;
      45812:data<=-16'd10945;
      45813:data<=-16'd2588;
      45814:data<=16'd11791;
      45815:data<=16'd18457;
      45816:data<=16'd14803;
      45817:data<=16'd13391;
      45818:data<=16'd13993;
      45819:data<=16'd9576;
      45820:data<=16'd12589;
      45821:data<=16'd18151;
      45822:data<=16'd10863;
      45823:data<=16'd7697;
      45824:data<=16'd10378;
      45825:data<=16'd6094;
      45826:data<=16'd9831;
      45827:data<=16'd16213;
      45828:data<=16'd8056;
      45829:data<=16'd5121;
      45830:data<=16'd15461;
      45831:data<=16'd18258;
      45832:data<=16'd12342;
      45833:data<=16'd10434;
      45834:data<=16'd10416;
      45835:data<=16'd10308;
      45836:data<=16'd14292;
      45837:data<=16'd14549;
      45838:data<=16'd11019;
      45839:data<=16'd14169;
      45840:data<=16'd14871;
      45841:data<=16'd11044;
      45842:data<=16'd12881;
      45843:data<=16'd11523;
      45844:data<=16'd6135;
      45845:data<=16'd6387;
      45846:data<=16'd8469;
      45847:data<=16'd9972;
      45848:data<=16'd9453;
      45849:data<=16'd6868;
      45850:data<=16'd6736;
      45851:data<=16'd8002;
      45852:data<=16'd9981;
      45853:data<=16'd9594;
      45854:data<=16'd9351;
      45855:data<=16'd12000;
      45856:data<=16'd1542;
      45857:data<=-16'd9858;
      45858:data<=-16'd2783;
      45859:data<=-16'd5049;
      45860:data<=-16'd14774;
      45861:data<=-16'd6633;
      45862:data<=-16'd1624;
      45863:data<=-16'd7915;
      45864:data<=-16'd11629;
      45865:data<=-16'd13192;
      45866:data<=-16'd10906;
      45867:data<=-16'd9824;
      45868:data<=-16'd9856;
      45869:data<=-16'd6253;
      45870:data<=-16'd9870;
      45871:data<=-16'd13057;
      45872:data<=-16'd7454;
      45873:data<=-16'd6228;
      45874:data<=-16'd8229;
      45875:data<=-16'd10824;
      45876:data<=-16'd12234;
      45877:data<=-16'd6956;
      45878:data<=-16'd5755;
      45879:data<=-16'd5521;
      45880:data<=16'd1130;
      45881:data<=16'd1324;
      45882:data<=-16'd707;
      45883:data<=16'd1515;
      45884:data<=16'd425;
      45885:data<=-16'd961;
      45886:data<=-16'd594;
      45887:data<=16'd2033;
      45888:data<=16'd4595;
      45889:data<=16'd39;
      45890:data<=16'd197;
      45891:data<=16'd7138;
      45892:data<=16'd3533;
      45893:data<=-16'd2795;
      45894:data<=16'd370;
      45895:data<=16'd3037;
      45896:data<=16'd705;
      45897:data<=16'd2634;
      45898:data<=16'd14055;
      45899:data<=16'd25029;
      45900:data<=16'd23887;
      45901:data<=16'd16116;
      45902:data<=16'd14416;
      45903:data<=16'd19080;
      45904:data<=16'd20263;
      45905:data<=16'd17719;
      45906:data<=16'd17379;
      45907:data<=16'd16628;
      45908:data<=16'd15576;
      45909:data<=16'd16363;
      45910:data<=16'd17581;
      45911:data<=16'd19813;
      45912:data<=16'd18882;
      45913:data<=16'd17873;
      45914:data<=16'd23710;
      45915:data<=16'd27338;
      45916:data<=16'd27599;
      45917:data<=16'd27678;
      45918:data<=16'd25244;
      45919:data<=16'd27887;
      45920:data<=16'd25755;
      45921:data<=16'd13852;
      45922:data<=16'd14007;
      45923:data<=16'd16581;
      45924:data<=16'd12690;
      45925:data<=16'd17637;
      45926:data<=16'd17091;
      45927:data<=16'd10501;
      45928:data<=16'd12933;
      45929:data<=16'd10851;
      45930:data<=16'd10107;
      45931:data<=16'd15253;
      45932:data<=16'd9359;
      45933:data<=16'd6052;
      45934:data<=16'd10038;
      45935:data<=16'd6922;
      45936:data<=16'd3862;
      45937:data<=16'd97;
      45938:data<=-16'd3729;
      45939:data<=-16'd726;
      45940:data<=-16'd7141;
      45941:data<=-16'd20422;
      45942:data<=-16'd21258;
      45943:data<=-16'd17584;
      45944:data<=-16'd16766;
      45945:data<=-16'd16260;
      45946:data<=-16'd17666;
      45947:data<=-16'd16678;
      45948:data<=-16'd13577;
      45949:data<=-16'd13916;
      45950:data<=-16'd14622;
      45951:data<=-16'd15047;
      45952:data<=-16'd17544;
      45953:data<=-16'd18042;
      45954:data<=-16'd16841;
      45955:data<=-16'd17159;
      45956:data<=-16'd16214;
      45957:data<=-16'd18040;
      45958:data<=-16'd22908;
      45959:data<=-16'd19221;
      45960:data<=-16'd16390;
      45961:data<=-16'd21828;
      45962:data<=-16'd18472;
      45963:data<=-16'd16236;
      45964:data<=-16'd24385;
      45965:data<=-16'd22463;
      45966:data<=-16'd21787;
      45967:data<=-16'd29379;
      45968:data<=-16'd22709;
      45969:data<=-16'd18295;
      45970:data<=-16'd24480;
      45971:data<=-16'd18022;
      45972:data<=-16'd15239;
      45973:data<=-16'd25417;
      45974:data<=-16'd24212;
      45975:data<=-16'd17538;
      45976:data<=-16'd19569;
      45977:data<=-16'd22589;
      45978:data<=-16'd21748;
      45979:data<=-16'd18871;
      45980:data<=-16'd17838;
      45981:data<=-16'd16589;
      45982:data<=-16'd7996;
      45983:data<=16'd1101;
      45984:data<=16'd294;
      45985:data<=-16'd3227;
      45986:data<=-16'd2046;
      45987:data<=-16'd4980;
      45988:data<=-16'd8710;
      45989:data<=-16'd38;
      45990:data<=16'd4090;
      45991:data<=-16'd6172;
      45992:data<=-16'd8261;
      45993:data<=-16'd2532;
      45994:data<=-16'd707;
      45995:data<=16'd103;
      45996:data<=-16'd3334;
      45997:data<=-16'd4129;
      45998:data<=16'd1544;
      45999:data<=16'd963;
      46000:data<=-16'd2017;
      46001:data<=-16'd3947;
      46002:data<=-16'd3368;
      46003:data<=16'd3576;
      46004:data<=-16'd1119;
      46005:data<=-16'd8220;
      46006:data<=16'd1172;
      46007:data<=-16'd303;
      46008:data<=-16'd8343;
      46009:data<=-16'd723;
      46010:data<=16'd234;
      46011:data<=-16'd3480;
      46012:data<=-16'd1014;
      46013:data<=-16'd5661;
      46014:data<=-16'd4902;
      46015:data<=16'd3401;
      46016:data<=16'd4522;
      46017:data<=16'd6299;
      46018:data<=16'd4927;
      46019:data<=-16'd796;
      46020:data<=16'd3140;
      46021:data<=16'd6857;
      46022:data<=16'd3542;
      46023:data<=16'd1586;
      46024:data<=-16'd2861;
      46025:data<=-16'd12082;
      46026:data<=-16'd17743;
      46027:data<=-16'd13778;
      46028:data<=-16'd8725;
      46029:data<=-16'd11000;
      46030:data<=-16'd8664;
      46031:data<=-16'd1595;
      46032:data<=-16'd3980;
      46033:data<=-16'd9377;
      46034:data<=-16'd9524;
      46035:data<=-16'd5997;
      46036:data<=-16'd1683;
      46037:data<=-16'd3803;
      46038:data<=-16'd5882;
      46039:data<=-16'd682;
      46040:data<=-16'd1227;
      46041:data<=-16'd6710;
      46042:data<=-16'd4470;
      46043:data<=-16'd2108;
      46044:data<=-16'd3924;
      46045:data<=16'd1894;
      46046:data<=16'd10859;
      46047:data<=16'd8975;
      46048:data<=16'd5618;
      46049:data<=16'd10707;
      46050:data<=16'd13019;
      46051:data<=16'd10378;
      46052:data<=16'd10031;
      46053:data<=16'd10194;
      46054:data<=16'd11075;
      46055:data<=16'd11997;
      46056:data<=16'd10839;
      46057:data<=16'd11606;
      46058:data<=16'd11634;
      46059:data<=16'd8907;
      46060:data<=16'd8987;
      46061:data<=16'd9782;
      46062:data<=16'd10026;
      46063:data<=16'd10795;
      46064:data<=16'd5930;
      46065:data<=16'd337;
      46066:data<=16'd6866;
      46067:data<=16'd19637;
      46068:data<=16'd24318;
      46069:data<=16'd21420;
      46070:data<=16'd19288;
      46071:data<=16'd19212;
      46072:data<=16'd19000;
      46073:data<=16'd18624;
      46074:data<=16'd18145;
      46075:data<=16'd18224;
      46076:data<=16'd18683;
      46077:data<=16'd17807;
      46078:data<=16'd16619;
      46079:data<=16'd17083;
      46080:data<=16'd17857;
      46081:data<=16'd16399;
      46082:data<=16'd14462;
      46083:data<=16'd15162;
      46084:data<=16'd15432;
      46085:data<=16'd14210;
      46086:data<=16'd15597;
      46087:data<=16'd16732;
      46088:data<=16'd14283;
      46089:data<=16'd12930;
      46090:data<=16'd14421;
      46091:data<=16'd14942;
      46092:data<=16'd13599;
      46093:data<=16'd12988;
      46094:data<=16'd12771;
      46095:data<=16'd11502;
      46096:data<=16'd10724;
      46097:data<=16'd9700;
      46098:data<=16'd9229;
      46099:data<=16'd11570;
      46100:data<=16'd11935;
      46101:data<=16'd10604;
      46102:data<=16'd11217;
      46103:data<=16'd10316;
      46104:data<=16'd10035;
      46105:data<=16'd10314;
      46106:data<=16'd8334;
      46107:data<=16'd10154;
      46108:data<=16'd7100;
      46109:data<=-16'd6683;
      46110:data<=-16'd10981;
      46111:data<=-16'd6285;
      46112:data<=-16'd7210;
      46113:data<=-16'd5753;
      46114:data<=-16'd364;
      46115:data<=16'd1213;
      46116:data<=16'd2181;
      46117:data<=16'd3698;
      46118:data<=16'd4020;
      46119:data<=16'd4137;
      46120:data<=16'd3927;
      46121:data<=16'd2931;
      46122:data<=16'd1967;
      46123:data<=16'd2608;
      46124:data<=16'd2434;
      46125:data<=16'd629;
      46126:data<=16'd980;
      46127:data<=16'd1104;
      46128:data<=16'd306;
      46129:data<=16'd826;
      46130:data<=-16'd743;
      46131:data<=-16'd2027;
      46132:data<=-16'd1858;
      46133:data<=-16'd3921;
      46134:data<=-16'd3700;
      46135:data<=-16'd3037;
      46136:data<=-16'd5656;
      46137:data<=-16'd5156;
      46138:data<=-16'd4196;
      46139:data<=-16'd5463;
      46140:data<=-16'd4143;
      46141:data<=-16'd3783;
      46142:data<=-16'd6096;
      46143:data<=-16'd7517;
      46144:data<=-16'd7145;
      46145:data<=-16'd6264;
      46146:data<=-16'd7602;
      46147:data<=-16'd6548;
      46148:data<=-16'd4402;
      46149:data<=-16'd8721;
      46150:data<=-16'd5084;
      46151:data<=16'd9265;
      46152:data<=16'd11632;
      46153:data<=16'd6746;
      46154:data<=16'd8003;
      46155:data<=16'd7780;
      46156:data<=16'd6138;
      46157:data<=16'd5169;
      46158:data<=16'd2376;
      46159:data<=16'd2961;
      46160:data<=16'd4664;
      46161:data<=16'd2165;
      46162:data<=16'd174;
      46163:data<=-16'd914;
      46164:data<=-16'd4320;
      46165:data<=-16'd7054;
      46166:data<=-16'd7656;
      46167:data<=-16'd8722;
      46168:data<=-16'd9597;
      46169:data<=-16'd9320;
      46170:data<=-16'd9812;
      46171:data<=-16'd9100;
      46172:data<=-16'd7259;
      46173:data<=-16'd9213;
      46174:data<=-16'd11053;
      46175:data<=-16'd9283;
      46176:data<=-16'd9116;
      46177:data<=-16'd9917;
      46178:data<=-16'd10140;
      46179:data<=-16'd11505;
      46180:data<=-16'd11188;
      46181:data<=-16'd9746;
      46182:data<=-16'd10290;
      46183:data<=-16'd11232;
      46184:data<=-16'd10686;
      46185:data<=-16'd9100;
      46186:data<=-16'd9632;
      46187:data<=-16'd10860;
      46188:data<=-16'd9335;
      46189:data<=-16'd10295;
      46190:data<=-16'd11485;
      46191:data<=-16'd8530;
      46192:data<=-16'd14446;
      46193:data<=-16'd27660;
      46194:data<=-16'd30327;
      46195:data<=-16'd27429;
      46196:data<=-16'd28004;
      46197:data<=-16'd26793;
      46198:data<=-16'd25029;
      46199:data<=-16'd25131;
      46200:data<=-16'd23737;
      46201:data<=-16'd22905;
      46202:data<=-16'd23940;
      46203:data<=-16'd23096;
      46204:data<=-16'd21776;
      46205:data<=-16'd22621;
      46206:data<=-16'd21776;
      46207:data<=-16'd19047;
      46208:data<=-16'd18504;
      46209:data<=-16'd17599;
      46210:data<=-16'd15850;
      46211:data<=-16'd16672;
      46212:data<=-16'd17058;
      46213:data<=-16'd16368;
      46214:data<=-16'd14888;
      46215:data<=-16'd8856;
      46216:data<=-16'd4748;
      46217:data<=-16'd7627;
      46218:data<=-16'd9541;
      46219:data<=-16'd8778;
      46220:data<=-16'd7753;
      46221:data<=-16'd5806;
      46222:data<=-16'd5774;
      46223:data<=-16'd6361;
      46224:data<=-16'd5010;
      46225:data<=-16'd4704;
      46226:data<=-16'd4866;
      46227:data<=-16'd4077;
      46228:data<=-16'd3758;
      46229:data<=-16'd4178;
      46230:data<=-16'd3823;
      46231:data<=16'd8;
      46232:data<=16'd1809;
      46233:data<=-16'd1670;
      46234:data<=16'd3497;
      46235:data<=16'd16803;
      46236:data<=16'd20803;
      46237:data<=16'd19103;
      46238:data<=16'd20528;
      46239:data<=16'd20525;
      46240:data<=16'd19281;
      46241:data<=16'd18850;
      46242:data<=16'd18630;
      46243:data<=16'd19332;
      46244:data<=16'd19014;
      46245:data<=16'd18158;
      46246:data<=16'd18089;
      46247:data<=16'd17155;
      46248:data<=16'd17499;
      46249:data<=16'd18844;
      46250:data<=16'd17233;
      46251:data<=16'd15109;
      46252:data<=16'd15482;
      46253:data<=16'd15594;
      46254:data<=16'd13687;
      46255:data<=16'd13591;
      46256:data<=16'd16506;
      46257:data<=16'd17098;
      46258:data<=16'd15797;
      46259:data<=16'd15594;
      46260:data<=16'd14046;
      46261:data<=16'd13373;
      46262:data<=16'd14807;
      46263:data<=16'd14322;
      46264:data<=16'd12569;
      46265:data<=16'd8869;
      46266:data<=16'd4948;
      46267:data<=16'd6270;
      46268:data<=16'd7389;
      46269:data<=16'd5594;
      46270:data<=16'd5802;
      46271:data<=16'd6149;
      46272:data<=16'd6093;
      46273:data<=16'd5615;
      46274:data<=16'd5013;
      46275:data<=16'd7870;
      46276:data<=16'd4429;
      46277:data<=-16'd8599;
      46278:data<=-16'd14243;
      46279:data<=-16'd11872;
      46280:data<=-16'd10806;
      46281:data<=-16'd9512;
      46282:data<=-16'd9423;
      46283:data<=-16'd8884;
      46284:data<=-16'd5539;
      46285:data<=-16'd5671;
      46286:data<=-16'd6545;
      46287:data<=-16'd3845;
      46288:data<=-16'd3104;
      46289:data<=-16'd3917;
      46290:data<=-16'd3589;
      46291:data<=-16'd3798;
      46292:data<=-16'd3068;
      46293:data<=-16'd922;
      46294:data<=-16'd182;
      46295:data<=-16'd902;
      46296:data<=-16'd622;
      46297:data<=16'd649;
      46298:data<=16'd294;
      46299:data<=-16'd544;
      46300:data<=16'd967;
      46301:data<=16'd2520;
      46302:data<=16'd2097;
      46303:data<=16'd1764;
      46304:data<=16'd1823;
      46305:data<=16'd1732;
      46306:data<=16'd3243;
      46307:data<=16'd4711;
      46308:data<=16'd3233;
      46309:data<=16'd2124;
      46310:data<=16'd2710;
      46311:data<=16'd2945;
      46312:data<=16'd4422;
      46313:data<=16'd4814;
      46314:data<=16'd5063;
      46315:data<=16'd11876;
      46316:data<=16'd15258;
      46317:data<=16'd10176;
      46318:data<=16'd15279;
      46319:data<=16'd29241;
      46320:data<=16'd32687;
      46321:data<=16'd28415;
      46322:data<=16'd26729;
      46323:data<=16'd27285;
      46324:data<=16'd27287;
      46325:data<=16'd25570;
      46326:data<=16'd24160;
      46327:data<=16'd22885;
      46328:data<=16'd20644;
      46329:data<=16'd20262;
      46330:data<=16'd19619;
      46331:data<=16'd16789;
      46332:data<=16'd15696;
      46333:data<=16'd15217;
      46334:data<=16'd13916;
      46335:data<=16'd13373;
      46336:data<=16'd11412;
      46337:data<=16'd8643;
      46338:data<=16'd7921;
      46339:data<=16'd8149;
      46340:data<=16'd8105;
      46341:data<=16'd6922;
      46342:data<=16'd5194;
      46343:data<=16'd4805;
      46344:data<=16'd4605;
      46345:data<=16'd3894;
      46346:data<=16'd2977;
      46347:data<=16'd1683;
      46348:data<=16'd1350;
      46349:data<=16'd814;
      46350:data<=-16'd575;
      46351:data<=-16'd743;
      46352:data<=-16'd1727;
      46353:data<=-16'd2667;
      46354:data<=-16'd855;
      46355:data<=-16'd1481;
      46356:data<=-16'd4297;
      46357:data<=-16'd4746;
      46358:data<=-16'd5254;
      46359:data<=-16'd4773;
      46360:data<=-16'd7007;
      46361:data<=-16'd19200;
      46362:data<=-16'd27322;
      46363:data<=-16'd23494;
      46364:data<=-16'd24504;
      46365:data<=-16'd31196;
      46366:data<=-16'd31921;
      46367:data<=-16'd30406;
      46368:data<=-16'd30518;
      46369:data<=-16'd30370;
      46370:data<=-16'd30045;
      46371:data<=-16'd28395;
      46372:data<=-16'd26098;
      46373:data<=-16'd25131;
      46374:data<=-16'd25319;
      46375:data<=-16'd25975;
      46376:data<=-16'd25560;
      46377:data<=-16'd25076;
      46378:data<=-16'd25445;
      46379:data<=-16'd23830;
      46380:data<=-16'd22538;
      46381:data<=-16'd24169;
      46382:data<=-16'd23913;
      46383:data<=-16'd21799;
      46384:data<=-16'd21681;
      46385:data<=-16'd21443;
      46386:data<=-16'd20651;
      46387:data<=-16'd21046;
      46388:data<=-16'd20234;
      46389:data<=-16'd18569;
      46390:data<=-16'd18451;
      46391:data<=-16'd17920;
      46392:data<=-16'd17444;
      46393:data<=-16'd18321;
      46394:data<=-16'd17508;
      46395:data<=-16'd16653;
      46396:data<=-16'd17535;
      46397:data<=-16'd16271;
      46398:data<=-16'd14619;
      46399:data<=-16'd14545;
      46400:data<=-16'd14110;
      46401:data<=-16'd14616;
      46402:data<=-16'd11022;
      46403:data<=-16'd567;
      46404:data<=16'd5832;
      46405:data<=16'd6105;
      46406:data<=16'd6029;
      46407:data<=16'd4549;
      46408:data<=16'd3063;
      46409:data<=16'd2786;
      46410:data<=16'd2369;
      46411:data<=16'd2654;
      46412:data<=16'd1158;
      46413:data<=-16'd795;
      46414:data<=16'd2261;
      46415:data<=16'd7473;
      46416:data<=16'd9931;
      46417:data<=16'd8702;
      46418:data<=16'd6417;
      46419:data<=16'd6886;
      46420:data<=16'd7692;
      46421:data<=16'd6942;
      46422:data<=16'd6793;
      46423:data<=16'd6939;
      46424:data<=16'd7512;
      46425:data<=16'd7730;
      46426:data<=16'd7288;
      46427:data<=16'd8307;
      46428:data<=16'd7903;
      46429:data<=16'd6316;
      46430:data<=16'd7389;
      46431:data<=16'd7565;
      46432:data<=16'd6619;
      46433:data<=16'd7385;
      46434:data<=16'd7421;
      46435:data<=16'd7092;
      46436:data<=16'd7517;
      46437:data<=16'd8326;
      46438:data<=16'd9078;
      46439:data<=16'd7788;
      46440:data<=16'd7406;
      46441:data<=16'd8428;
      46442:data<=16'd7708;
      46443:data<=16'd9077;
      46444:data<=16'd7545;
      46445:data<=-16'd2864;
      46446:data<=-16'd9257;
      46447:data<=-16'd8631;
      46448:data<=-16'd9809;
      46449:data<=-16'd9259;
      46450:data<=-16'd6915;
      46451:data<=-16'd6862;
      46452:data<=-16'd5498;
      46453:data<=-16'd4423;
      46454:data<=-16'd5280;
      46455:data<=-16'd3686;
      46456:data<=-16'd1898;
      46457:data<=-16'd2150;
      46458:data<=-16'd1274;
      46459:data<=-16'd588;
      46460:data<=-16'd1048;
      46461:data<=-16'd252;
      46462:data<=16'd670;
      46463:data<=16'd1491;
      46464:data<=16'd1659;
      46465:data<=-16'd2736;
      46466:data<=-16'd6912;
      46467:data<=-16'd5369;
      46468:data<=-16'd4438;
      46469:data<=-16'd4658;
      46470:data<=-16'd1956;
      46471:data<=-16'd1131;
      46472:data<=-16'd2100;
      46473:data<=-16'd1027;
      46474:data<=16'd126;
      46475:data<=16'd1548;
      46476:data<=16'd2297;
      46477:data<=16'd1374;
      46478:data<=16'd2171;
      46479:data<=16'd2598;
      46480:data<=16'd2071;
      46481:data<=16'd3657;
      46482:data<=16'd3348;
      46483:data<=16'd2784;
      46484:data<=16'd5580;
      46485:data<=16'd5190;
      46486:data<=16'd6275;
      46487:data<=16'd17114;
      46488:data<=16'd25438;
      46489:data<=16'd23875;
      46490:data<=16'd21943;
      46491:data<=16'd22086;
      46492:data<=16'd21869;
      46493:data<=16'd22580;
      46494:data<=16'd22230;
      46495:data<=16'd20372;
      46496:data<=16'd20048;
      46497:data<=16'd19788;
      46498:data<=16'd18472;
      46499:data<=16'd18389;
      46500:data<=16'd18930;
      46501:data<=16'd18710;
      46502:data<=16'd18169;
      46503:data<=16'd17423;
      46504:data<=16'd16856;
      46505:data<=16'd16474;
      46506:data<=16'd16198;
      46507:data<=16'd16683;
      46508:data<=16'd16747;
      46509:data<=16'd15259;
      46510:data<=16'd14032;
      46511:data<=16'd14363;
      46512:data<=16'd14741;
      46513:data<=16'd13922;
      46514:data<=16'd13957;
      46515:data<=16'd16788;
      46516:data<=16'd19781;
      46517:data<=16'd19893;
      46518:data<=16'd18806;
      46519:data<=16'd19196;
      46520:data<=16'd19793;
      46521:data<=16'd18833;
      46522:data<=16'd17249;
      46523:data<=16'd15459;
      46524:data<=16'd14465;
      46525:data<=16'd15067;
      46526:data<=16'd14765;
      46527:data<=16'd14196;
      46528:data<=16'd12408;
      46529:data<=16'd3289;
      46530:data<=-16'd6980;
      46531:data<=-16'd9374;
      46532:data<=-16'd9536;
      46533:data<=-16'd10381;
      46534:data<=-16'd10011;
      46535:data<=-16'd10163;
      46536:data<=-16'd9327;
      46537:data<=-16'd9119;
      46538:data<=-16'd10928;
      46539:data<=-16'd9755;
      46540:data<=-16'd8652;
      46541:data<=-16'd10076;
      46542:data<=-16'd9142;
      46543:data<=-16'd9001;
      46544:data<=-16'd11086;
      46545:data<=-16'd10856;
      46546:data<=-16'd10381;
      46547:data<=-16'd10475;
      46548:data<=-16'd9444;
      46549:data<=-16'd9668;
      46550:data<=-16'd11089;
      46551:data<=-16'd11583;
      46552:data<=-16'd11532;
      46553:data<=-16'd11606;
      46554:data<=-16'd11153;
      46555:data<=-16'd10806;
      46556:data<=-16'd12266;
      46557:data<=-16'd12634;
      46558:data<=-16'd10628;
      46559:data<=-16'd10329;
      46560:data<=-16'd10316;
      46561:data<=-16'd9938;
      46562:data<=-16'd12246;
      46563:data<=-16'd12813;
      46564:data<=-16'd11467;
      46565:data<=-16'd14499;
      46566:data<=-16'd18785;
      46567:data<=-16'd19136;
      46568:data<=-16'd17569;
      46569:data<=-16'd18172;
      46570:data<=-16'd18131;
      46571:data<=-16'd10064;
      46572:data<=-16'd346;
      46573:data<=16'd1533;
      46574:data<=16'd560;
      46575:data<=-16'd860;
      46576:data<=-16'd2485;
      46577:data<=-16'd872;
      46578:data<=-16'd735;
      46579:data<=-16'd2024;
      46580:data<=-16'd1187;
      46581:data<=-16'd3510;
      46582:data<=-16'd5796;
      46583:data<=-16'd3395;
      46584:data<=-16'd2732;
      46585:data<=-16'd3545;
      46586:data<=-16'd3256;
      46587:data<=-16'd4673;
      46588:data<=-16'd5864;
      46589:data<=-16'd5109;
      46590:data<=-16'd4734;
      46591:data<=-16'd5127;
      46592:data<=-16'd4573;
      46593:data<=-16'd3724;
      46594:data<=-16'd5077;
      46595:data<=-16'd5600;
      46596:data<=-16'd4246;
      46597:data<=-16'd5454;
      46598:data<=-16'd5759;
      46599:data<=-16'd4622;
      46600:data<=-16'd7175;
      46601:data<=-16'd8005;
      46602:data<=-16'd6240;
      46603:data<=-16'd6722;
      46604:data<=-16'd5670;
      46605:data<=-16'd4716;
      46606:data<=-16'd6630;
      46607:data<=-16'd7028;
      46608:data<=-16'd6608;
      46609:data<=-16'd6622;
      46610:data<=-16'd6898;
      46611:data<=-16'd6307;
      46612:data<=-16'd4749;
      46613:data<=-16'd13038;
      46614:data<=-16'd25858;
      46615:data<=-16'd23062;
      46616:data<=-16'd14883;
      46617:data<=-16'd14612;
      46618:data<=-16'd13641;
      46619:data<=-16'd13415;
      46620:data<=-16'd14686;
      46621:data<=-16'd12333;
      46622:data<=-16'd12091;
      46623:data<=-16'd12314;
      46624:data<=-16'd10096;
      46625:data<=-16'd10883;
      46626:data<=-16'd10681;
      46627:data<=-16'd8276;
      46628:data<=-16'd8307;
      46629:data<=-16'd7708;
      46630:data<=-16'd6904;
      46631:data<=-16'd6484;
      46632:data<=-16'd3697;
      46633:data<=-16'd2830;
      46634:data<=-16'd3767;
      46635:data<=-16'd2563;
      46636:data<=-16'd2638;
      46637:data<=-16'd3045;
      46638:data<=-16'd494;
      46639:data<=16'd647;
      46640:data<=16'd18;
      46641:data<=16'd1427;
      46642:data<=16'd2130;
      46643:data<=16'd1528;
      46644:data<=16'd3142;
      46645:data<=16'd3967;
      46646:data<=16'd3465;
      46647:data<=16'd5048;
      46648:data<=16'd4764;
      46649:data<=16'd4153;
      46650:data<=16'd7025;
      46651:data<=16'd6708;
      46652:data<=16'd5864;
      46653:data<=16'd7538;
      46654:data<=16'd5303;
      46655:data<=16'd9966;
      46656:data<=16'd23516;
      46657:data<=16'd26141;
      46658:data<=16'd22638;
      46659:data<=16'd23925;
      46660:data<=16'd22768;
      46661:data<=16'd21164;
      46662:data<=16'd21046;
      46663:data<=16'd20265;
      46664:data<=16'd22462;
      46665:data<=16'd20760;
      46666:data<=16'd13394;
      46667:data<=16'd11118;
      46668:data<=16'd12158;
      46669:data<=16'd12516;
      46670:data<=16'd13132;
      46671:data<=16'd12141;
      46672:data<=16'd12107;
      46673:data<=16'd12700;
      46674:data<=16'd11207;
      46675:data<=16'd11427;
      46676:data<=16'd12433;
      46677:data<=16'd11775;
      46678:data<=16'd11882;
      46679:data<=16'd11791;
      46680:data<=16'd11162;
      46681:data<=16'd11708;
      46682:data<=16'd11981;
      46683:data<=16'd11365;
      46684:data<=16'd11133;
      46685:data<=16'd11025;
      46686:data<=16'd10237;
      46687:data<=16'd10505;
      46688:data<=16'd11934;
      46689:data<=16'd11808;
      46690:data<=16'd11853;
      46691:data<=16'd11553;
      46692:data<=16'd8875;
      46693:data<=16'd9257;
      46694:data<=16'd10928;
      46695:data<=16'd10763;
      46696:data<=16'd12619;
      46697:data<=16'd6875;
      46698:data<=-16'd6602;
      46699:data<=-16'd9509;
      46700:data<=-16'd6628;
      46701:data<=-16'd7236;
      46702:data<=-16'd5250;
      46703:data<=-16'd4264;
      46704:data<=-16'd5333;
      46705:data<=-16'd4018;
      46706:data<=-16'd3222;
      46707:data<=-16'd1692;
      46708:data<=-16'd754;
      46709:data<=-16'd2118;
      46710:data<=-16'd1715;
      46711:data<=-16'd2999;
      46712:data<=-16'd2887;
      46713:data<=16'd1894;
      46714:data<=16'd839;
      46715:data<=16'd669;
      46716:data<=16'd8624;
      46717:data<=16'd10372;
      46718:data<=16'd7868;
      46719:data<=16'd9959;
      46720:data<=16'd10075;
      46721:data<=16'd8276;
      46722:data<=16'd7597;
      46723:data<=16'd6713;
      46724:data<=16'd6746;
      46725:data<=16'd5877;
      46726:data<=16'd4582;
      46727:data<=16'd5506;
      46728:data<=16'd5275;
      46729:data<=16'd3597;
      46730:data<=16'd3853;
      46731:data<=16'd3821;
      46732:data<=16'd1600;
      46733:data<=16'd1309;
      46734:data<=16'd2264;
      46735:data<=16'd328;
      46736:data<=16'd845;
      46737:data<=16'd2020;
      46738:data<=-16'd2758;
      46739:data<=16'd1254;
      46740:data<=16'd15030;
      46741:data<=16'd16901;
      46742:data<=16'd13444;
      46743:data<=16'd15070;
      46744:data<=16'd11746;
      46745:data<=16'd8370;
      46746:data<=16'd9495;
      46747:data<=16'd8106;
      46748:data<=16'd7928;
      46749:data<=16'd8646;
      46750:data<=16'd5879;
      46751:data<=16'd4278;
      46752:data<=16'd4302;
      46753:data<=16'd3472;
      46754:data<=16'd2399;
      46755:data<=16'd1674;
      46756:data<=16'd1477;
      46757:data<=16'd45;
      46758:data<=-16'd1368;
      46759:data<=-16'd1466;
      46760:data<=-16'd2015;
      46761:data<=-16'd1585;
      46762:data<=-16'd2414;
      46763:data<=-16'd4673;
      46764:data<=-16'd3301;
      46765:data<=-16'd5216;
      46766:data<=-16'd11887;
      46767:data<=-16'd12759;
      46768:data<=-16'd11840;
      46769:data<=-16'd14193;
      46770:data<=-16'd14650;
      46771:data<=-16'd13347;
      46772:data<=-16'd12170;
      46773:data<=-16'd11840;
      46774:data<=-16'd12323;
      46775:data<=-16'd12680;
      46776:data<=-16'd13802;
      46777:data<=-16'd13588;
      46778:data<=-16'd13722;
      46779:data<=-16'd15023;
      46780:data<=-16'd11987;
      46781:data<=-16'd15675;
      46782:data<=-16'd30068;
      46783:data<=-16'd34270;
      46784:data<=-16'd30495;
      46785:data<=-16'd31181;
      46786:data<=-16'd28958;
      46787:data<=-16'd26774;
      46788:data<=-16'd28767;
      46789:data<=-16'd28269;
      46790:data<=-16'd27378;
      46791:data<=-16'd26059;
      46792:data<=-16'd23820;
      46793:data<=-16'd24858;
      46794:data<=-16'd24441;
      46795:data<=-16'd22278;
      46796:data<=-16'd22489;
      46797:data<=-16'd21732;
      46798:data<=-16'd20710;
      46799:data<=-16'd20359;
      46800:data<=-16'd19464;
      46801:data<=-16'd20193;
      46802:data<=-16'd20019;
      46803:data<=-16'd18337;
      46804:data<=-16'd18290;
      46805:data<=-16'd17752;
      46806:data<=-16'd16935;
      46807:data<=-16'd17209;
      46808:data<=-16'd17009;
      46809:data<=-16'd16985;
      46810:data<=-16'd16581;
      46811:data<=-16'd14854;
      46812:data<=-16'd13591;
      46813:data<=-16'd14625;
      46814:data<=-16'd16271;
      46815:data<=-16'd13173;
      46816:data<=-16'd7224;
      46817:data<=-16'd4205;
      46818:data<=-16'd3553;
      46819:data<=-16'd5139;
      46820:data<=-16'd5281;
      46821:data<=-16'd2884;
      46822:data<=-16'd4679;
      46823:data<=-16'd567;
      46824:data<=16'd13526;
      46825:data<=16'd17333;
      46826:data<=16'd13443;
      46827:data<=16'd14965;
      46828:data<=16'd14587;
      46829:data<=16'd12786;
      46830:data<=16'd13245;
      46831:data<=16'd13112;
      46832:data<=16'd14924;
      46833:data<=16'd15409;
      46834:data<=16'd13687;
      46835:data<=16'd14687;
      46836:data<=16'd14234;
      46837:data<=16'd13009;
      46838:data<=16'd14187;
      46839:data<=16'd14305;
      46840:data<=16'd14660;
      46841:data<=16'd14358;
      46842:data<=16'd12530;
      46843:data<=16'd13479;
      46844:data<=16'd14527;
      46845:data<=16'd14078;
      46846:data<=16'd14199;
      46847:data<=16'd14087;
      46848:data<=16'd14759;
      46849:data<=16'd14324;
      46850:data<=16'd13179;
      46851:data<=16'd14821;
      46852:data<=16'd14727;
      46853:data<=16'd13270;
      46854:data<=16'd13697;
      46855:data<=16'd12941;
      46856:data<=16'd13368;
      46857:data<=16'd14636;
      46858:data<=16'd13958;
      46859:data<=16'd14539;
      46860:data<=16'd14045;
      46861:data<=16'd12466;
      46862:data<=16'd12202;
      46863:data<=16'd11617;
      46864:data<=16'd13985;
      46865:data<=16'd9717;
      46866:data<=-16'd7885;
      46867:data<=-16'd16636;
      46868:data<=-16'd13332;
      46869:data<=-16'd13094;
      46870:data<=-16'd11414;
      46871:data<=-16'd9665;
      46872:data<=-16'd11182;
      46873:data<=-16'd9095;
      46874:data<=-16'd8008;
      46875:data<=-16'd7817;
      46876:data<=-16'd4507;
      46877:data<=-16'd5101;
      46878:data<=-16'd6228;
      46879:data<=-16'd4027;
      46880:data<=-16'd4032;
      46881:data<=-16'd3341;
      46882:data<=-16'd1563;
      46883:data<=-16'd1952;
      46884:data<=-16'd1406;
      46885:data<=-16'd884;
      46886:data<=-16'd1363;
      46887:data<=-16'd505;
      46888:data<=16'd229;
      46889:data<=16'd253;
      46890:data<=16'd591;
      46891:data<=16'd1262;
      46892:data<=16'd1433;
      46893:data<=16'd675;
      46894:data<=16'd1589;
      46895:data<=16'd3827;
      46896:data<=16'd4050;
      46897:data<=16'd2807;
      46898:data<=16'd1885;
      46899:data<=16'd2406;
      46900:data<=16'd3516;
      46901:data<=16'd3965;
      46902:data<=16'd4529;
      46903:data<=16'd3993;
      46904:data<=16'd4234;
      46905:data<=16'd5623;
      46906:data<=16'd4165;
      46907:data<=16'd9359;
      46908:data<=16'd22222;
      46909:data<=16'd24890;
      46910:data<=16'd22168;
      46911:data<=16'd23773;
      46912:data<=16'd21775;
      46913:data<=16'd20829;
      46914:data<=16'd22624;
      46915:data<=16'd20638;
      46916:data<=16'd23294;
      46917:data<=16'd27856;
      46918:data<=16'd25751;
      46919:data<=16'd25633;
      46920:data<=16'd27267;
      46921:data<=16'd25253;
      46922:data<=16'd23507;
      46923:data<=16'd22113;
      46924:data<=16'd21341;
      46925:data<=16'd21165;
      46926:data<=16'd19324;
      46927:data<=16'd18390;
      46928:data<=16'd17520;
      46929:data<=16'd15857;
      46930:data<=16'd16272;
      46931:data<=16'd15791;
      46932:data<=16'd13376;
      46933:data<=16'd11964;
      46934:data<=16'd11116;
      46935:data<=16'd10433;
      46936:data<=16'd9442;
      46937:data<=16'd8169;
      46938:data<=16'd7291;
      46939:data<=16'd6673;
      46940:data<=16'd6714;
      46941:data<=16'd5266;
      46942:data<=16'd3428;
      46943:data<=16'd4181;
      46944:data<=16'd3134;
      46945:data<=16'd849;
      46946:data<=-16'd68;
      46947:data<=-16'd1488;
      46948:data<=16'd302;
      46949:data<=-16'd2083;
      46950:data<=-16'd15534;
      46951:data<=-16'd22488;
      46952:data<=-16'd20412;
      46953:data<=-16'd21420;
      46954:data<=-16'd20212;
      46955:data<=-16'd17955;
      46956:data<=-16'd19676;
      46957:data<=-16'd19908;
      46958:data<=-16'd19926;
      46959:data<=-16'd19704;
      46960:data<=-16'd18048;
      46961:data<=-16'd18581;
      46962:data<=-16'd18404;
      46963:data<=-16'd18839;
      46964:data<=-16'd20301;
      46965:data<=-16'd17462;
      46966:data<=-16'd19064;
      46967:data<=-16'd25854;
      46968:data<=-16'd25452;
      46969:data<=-16'd23529;
      46970:data<=-16'd25247;
      46971:data<=-16'd24630;
      46972:data<=-16'd23825;
      46973:data<=-16'd23916;
      46974:data<=-16'd22606;
      46975:data<=-16'd22306;
      46976:data<=-16'd23316;
      46977:data<=-16'd23355;
      46978:data<=-16'd21972;
      46979:data<=-16'd20630;
      46980:data<=-16'd20007;
      46981:data<=-16'd19999;
      46982:data<=-16'd21112;
      46983:data<=-16'd21202;
      46984:data<=-16'd20374;
      46985:data<=-16'd20515;
      46986:data<=-16'd18777;
      46987:data<=-16'd16754;
      46988:data<=-16'd16904;
      46989:data<=-16'd17129;
      46990:data<=-16'd18057;
      46991:data<=-16'd13179;
      46992:data<=-16'd563;
      46993:data<=16'd4475;
      46994:data<=16'd2002;
      46995:data<=16'd2713;
      46996:data<=16'd2689;
      46997:data<=16'd1272;
      46998:data<=16'd1588;
      46999:data<=16'd1553;
      47000:data<=16'd1445;
      47001:data<=16'd317;
      47002:data<=-16'd722;
      47003:data<=16'd332;
      47004:data<=16'd256;
      47005:data<=16'd299;
      47006:data<=16'd651;
      47007:data<=-16'd1301;
      47008:data<=-16'd1727;
      47009:data<=-16'd1198;
      47010:data<=-16'd1900;
      47011:data<=-16'd1251;
      47012:data<=-16'd1036;
      47013:data<=-16'd1337;
      47014:data<=-16'd1438;
      47015:data<=-16'd2504;
      47016:data<=16'd623;
      47017:data<=16'd6579;
      47018:data<=16'd7670;
      47019:data<=16'd6056;
      47020:data<=16'd5177;
      47021:data<=16'd4898;
      47022:data<=16'd5104;
      47023:data<=16'd5134;
      47024:data<=16'd5756;
      47025:data<=16'd5225;
      47026:data<=16'd3792;
      47027:data<=16'd4767;
      47028:data<=16'd4757;
      47029:data<=16'd3548;
      47030:data<=16'd3762;
      47031:data<=16'd3406;
      47032:data<=16'd4995;
      47033:data<=16'd3479;
      47034:data<=-16'd7366;
      47035:data<=-16'd13323;
      47036:data<=-16'd11264;
      47037:data<=-16'd12449;
      47038:data<=-16'd11186;
      47039:data<=-16'd6352;
      47040:data<=-16'd6372;
      47041:data<=-16'd7016;
      47042:data<=-16'd5862;
      47043:data<=-16'd5577;
      47044:data<=-16'd4434;
      47045:data<=-16'd3409;
      47046:data<=-16'd3251;
      47047:data<=-16'd2602;
      47048:data<=-16'd2121;
      47049:data<=-16'd1682;
      47050:data<=-16'd813;
      47051:data<=16'd475;
      47052:data<=16'd1430;
      47053:data<=16'd1751;
      47054:data<=16'd2649;
      47055:data<=16'd2423;
      47056:data<=16'd1422;
      47057:data<=16'd2776;
      47058:data<=16'd3811;
      47059:data<=16'd3576;
      47060:data<=16'd4115;
      47061:data<=16'd4076;
      47062:data<=16'd4253;
      47063:data<=16'd4672;
      47064:data<=16'd4881;
      47065:data<=16'd6202;
      47066:data<=16'd4137;
      47067:data<=-16'd870;
      47068:data<=-16'd2287;
      47069:data<=-16'd1770;
      47070:data<=-16'd503;
      47071:data<=16'd1454;
      47072:data<=16'd2059;
      47073:data<=16'd2943;
      47074:data<=16'd2135;
      47075:data<=16'd4623;
      47076:data<=16'd17399;
      47077:data<=16'd24811;
      47078:data<=16'd21849;
      47079:data<=16'd22686;
      47080:data<=16'd22328;
      47081:data<=16'd18494;
      47082:data<=16'd20494;
      47083:data<=16'd21937;
      47084:data<=16'd20027;
      47085:data<=16'd20228;
      47086:data<=16'd19418;
      47087:data<=16'd18061;
      47088:data<=16'd19186;
      47089:data<=16'd20128;
      47090:data<=16'd19247;
      47091:data<=16'd17835;
      47092:data<=16'd17623;
      47093:data<=16'd16959;
      47094:data<=16'd15622;
      47095:data<=16'd16821;
      47096:data<=16'd17518;
      47097:data<=16'd15772;
      47098:data<=16'd14960;
      47099:data<=16'd14563;
      47100:data<=16'd14765;
      47101:data<=16'd16189;
      47102:data<=16'd16662;
      47103:data<=16'd16224;
      47104:data<=16'd15338;
      47105:data<=16'd14704;
      47106:data<=16'd14099;
      47107:data<=16'd13194;
      47108:data<=16'd14343;
      47109:data<=16'd14562;
      47110:data<=16'd13097;
      47111:data<=16'd13712;
      47112:data<=16'd12122;
      47113:data<=16'd10803;
      47114:data<=16'd13004;
      47115:data<=16'd11306;
      47116:data<=16'd12342;
      47117:data<=16'd15713;
      47118:data<=16'd6343;
      47119:data<=-16'd2558;
      47120:data<=16'd202;
      47121:data<=16'd931;
      47122:data<=16'd140;
      47123:data<=16'd1509;
      47124:data<=16'd911;
      47125:data<=16'd1008;
      47126:data<=16'd858;
      47127:data<=16'd123;
      47128:data<=16'd438;
      47129:data<=-16'd1225;
      47130:data<=-16'd1786;
      47131:data<=-16'd948;
      47132:data<=-16'd2740;
      47133:data<=-16'd3515;
      47134:data<=-16'd3162;
      47135:data<=-16'd3815;
      47136:data<=-16'd3914;
      47137:data<=-16'd4300;
      47138:data<=-16'd4505;
      47139:data<=-16'd5056;
      47140:data<=-16'd6602;
      47141:data<=-16'd6495;
      47142:data<=-16'd6478;
      47143:data<=-16'd6889;
      47144:data<=-16'd6302;
      47145:data<=-16'd7521;
      47146:data<=-16'd8809;
      47147:data<=-16'd8669;
      47148:data<=-16'd8930;
      47149:data<=-16'd8185;
      47150:data<=-16'd7924;
      47151:data<=-16'd9295;
      47152:data<=-16'd10390;
      47153:data<=-16'd10948;
      47154:data<=-16'd9768;
      47155:data<=-16'd8869;
      47156:data<=-16'd9089;
      47157:data<=-16'd8510;
      47158:data<=-16'd10634;
      47159:data<=-16'd9567;
      47160:data<=16'd652;
      47161:data<=16'd7327;
      47162:data<=16'd7309;
      47163:data<=16'd7204;
      47164:data<=16'd5074;
      47165:data<=16'd4112;
      47166:data<=16'd3873;
      47167:data<=-16'd1172;
      47168:data<=-16'd3936;
      47169:data<=-16'd2505;
      47170:data<=-16'd3777;
      47171:data<=-16'd5785;
      47172:data<=-16'd5752;
      47173:data<=-16'd5521;
      47174:data<=-16'd5492;
      47175:data<=-16'd4984;
      47176:data<=-16'd5318;
      47177:data<=-16'd7341;
      47178:data<=-16'd7371;
      47179:data<=-16'd6351;
      47180:data<=-16'd7682;
      47181:data<=-16'd7028;
      47182:data<=-16'd5927;
      47183:data<=-16'd8155;
      47184:data<=-16'd8011;
      47185:data<=-16'd6875;
      47186:data<=-16'd7932;
      47187:data<=-16'd6628;
      47188:data<=-16'd5745;
      47189:data<=-16'd7967;
      47190:data<=-16'd8672;
      47191:data<=-16'd7539;
      47192:data<=-16'd6789;
      47193:data<=-16'd6919;
      47194:data<=-16'd6777;
      47195:data<=-16'd6956;
      47196:data<=-16'd9420;
      47197:data<=-16'd9474;
      47198:data<=-16'd7686;
      47199:data<=-16'd9498;
      47200:data<=-16'd8504;
      47201:data<=-16'd8252;
      47202:data<=-16'd19361;
      47203:data<=-16'd28133;
      47204:data<=-16'd26189;
      47205:data<=-16'd25141;
      47206:data<=-16'd24620;
      47207:data<=-16'd22378;
      47208:data<=-16'd23505;
      47209:data<=-16'd23958;
      47210:data<=-16'd21546;
      47211:data<=-16'd20651;
      47212:data<=-16'd20259;
      47213:data<=-16'd18967;
      47214:data<=-16'd18613;
      47215:data<=-16'd19170;
      47216:data<=-16'd18034;
      47217:data<=-16'd14079;
      47218:data<=-16'd10481;
      47219:data<=-16'd9712;
      47220:data<=-16'd10927;
      47221:data<=-16'd11879;
      47222:data<=-16'd10577;
      47223:data<=-16'd9409;
      47224:data<=-16'd9928;
      47225:data<=-16'd9169;
      47226:data<=-16'd8326;
      47227:data<=-16'd8754;
      47228:data<=-16'd8034;
      47229:data<=-16'd7297;
      47230:data<=-16'd7295;
      47231:data<=-16'd6893;
      47232:data<=-16'd6413;
      47233:data<=-16'd4999;
      47234:data<=-16'd3797;
      47235:data<=-16'd3751;
      47236:data<=-16'd3210;
      47237:data<=-16'd3380;
      47238:data<=-16'd2889;
      47239:data<=-16'd311;
      47240:data<=16'd745;
      47241:data<=16'd1445;
      47242:data<=16'd1858;
      47243:data<=16'd1724;
      47244:data<=16'd9348;
      47245:data<=16'd20274;
      47246:data<=16'd22013;
      47247:data<=16'd20198;
      47248:data<=16'd20914;
      47249:data<=16'd20392;
      47250:data<=16'd19302;
      47251:data<=16'd19382;
      47252:data<=16'd19928;
      47253:data<=16'd19861;
      47254:data<=16'd18722;
      47255:data<=16'd17923;
      47256:data<=16'd17098;
      47257:data<=16'd16827;
      47258:data<=16'd17987;
      47259:data<=16'd17722;
      47260:data<=16'd16728;
      47261:data<=16'd16769;
      47262:data<=16'd16369;
      47263:data<=16'd15825;
      47264:data<=16'd15192;
      47265:data<=16'd15435;
      47266:data<=16'd15808;
      47267:data<=16'd12474;
      47268:data<=16'd9301;
      47269:data<=16'd8940;
      47270:data<=16'd8599;
      47271:data<=16'd10170;
      47272:data<=16'd10618;
      47273:data<=16'd8581;
      47274:data<=16'd9723;
      47275:data<=16'd9846;
      47276:data<=16'd8586;
      47277:data<=16'd10848;
      47278:data<=16'd11063;
      47279:data<=16'd10078;
      47280:data<=16'd10311;
      47281:data<=16'd8194;
      47282:data<=16'd8495;
      47283:data<=16'd10216;
      47284:data<=16'd9867;
      47285:data<=16'd10223;
      47286:data<=16'd3277;
      47287:data<=-16'd8099;
      47288:data<=-16'd8828;
      47289:data<=-16'd5724;
      47290:data<=-16'd6237;
      47291:data<=-16'd5692;
      47292:data<=-16'd5765;
      47293:data<=-16'd6284;
      47294:data<=-16'd5691;
      47295:data<=-16'd5100;
      47296:data<=-16'd3375;
      47297:data<=-16'd2816;
      47298:data<=-16'd3400;
      47299:data<=-16'd2848;
      47300:data<=-16'd3430;
      47301:data<=-16'd3099;
      47302:data<=-16'd716;
      47303:data<=-16'd176;
      47304:data<=-16'd620;
      47305:data<=-16'd557;
      47306:data<=-16'd388;
      47307:data<=-16'd247;
      47308:data<=-16'd121;
      47309:data<=16'd895;
      47310:data<=16'd720;
      47311:data<=-16'd35;
      47312:data<=16'd1089;
      47313:data<=16'd658;
      47314:data<=16'd773;
      47315:data<=16'd2729;
      47316:data<=16'd1563;
      47317:data<=16'd3435;
      47318:data<=16'd8802;
      47319:data<=16'd8269;
      47320:data<=16'd7007;
      47321:data<=16'd8319;
      47322:data<=16'd8090;
      47323:data<=16'd8402;
      47324:data<=16'd8134;
      47325:data<=16'd8066;
      47326:data<=16'd8411;
      47327:data<=16'd5846;
      47328:data<=16'd10760;
      47329:data<=16'd22165;
      47330:data<=16'd23269;
      47331:data<=16'd20601;
      47332:data<=16'd21666;
      47333:data<=16'd18695;
      47334:data<=16'd15978;
      47335:data<=16'd16396;
      47336:data<=16'd14745;
      47337:data<=16'd13750;
      47338:data<=16'd13931;
      47339:data<=16'd12022;
      47340:data<=16'd9306;
      47341:data<=16'd8331;
      47342:data<=16'd9095;
      47343:data<=16'd8425;
      47344:data<=16'd7037;
      47345:data<=16'd6804;
      47346:data<=16'd5024;
      47347:data<=16'd3721;
      47348:data<=16'd4322;
      47349:data<=16'd3532;
      47350:data<=16'd2974;
      47351:data<=16'd2711;
      47352:data<=16'd1278;
      47353:data<=16'd579;
      47354:data<=-16'd362;
      47355:data<=-16'd1086;
      47356:data<=-16'd895;
      47357:data<=-16'd1575;
      47358:data<=-16'd1850;
      47359:data<=-16'd2687;
      47360:data<=-16'd3791;
      47361:data<=-16'd3224;
      47362:data<=-16'd3821;
      47363:data<=-16'd3486;
      47364:data<=-16'd3386;
      47365:data<=-16'd6630;
      47366:data<=-16'd5742;
      47367:data<=-16'd6617;
      47368:data<=-16'd13041;
      47369:data<=-16'd11814;
      47370:data<=-16'd15151;
      47371:data<=-16'd29696;
      47372:data<=-16'd32380;
      47373:data<=-16'd28277;
      47374:data<=-16'd29907;
      47375:data<=-16'd28360;
      47376:data<=-16'd27331;
      47377:data<=-16'd28750;
      47378:data<=-16'd26967;
      47379:data<=-16'd26436;
      47380:data<=-16'd25951;
      47381:data<=-16'd24168;
      47382:data<=-16'd24148;
      47383:data<=-16'd23717;
      47384:data<=-16'd23849;
      47385:data<=-16'd23634;
      47386:data<=-16'd21792;
      47387:data<=-16'd21707;
      47388:data<=-16'd20859;
      47389:data<=-16'd20145;
      47390:data<=-16'd21684;
      47391:data<=-16'd20659;
      47392:data<=-16'd19519;
      47393:data<=-16'd19855;
      47394:data<=-16'd18659;
      47395:data<=-16'd18680;
      47396:data<=-16'd19268;
      47397:data<=-16'd18917;
      47398:data<=-16'd18307;
      47399:data<=-16'd16628;
      47400:data<=-16'd16216;
      47401:data<=-16'd15907;
      47402:data<=-16'd15347;
      47403:data<=-16'd16692;
      47404:data<=-16'd15338;
      47405:data<=-16'd13852;
      47406:data<=-16'd14402;
      47407:data<=-16'd12137;
      47408:data<=-16'd12542;
      47409:data<=-16'd13352;
      47410:data<=-16'd11086;
      47411:data<=-16'd13521;
      47412:data<=-16'd8204;
      47413:data<=16'd6811;
      47414:data<=16'd8831;
      47415:data<=16'd4369;
      47416:data<=16'd5617;
      47417:data<=16'd6786;
      47418:data<=16'd10545;
      47419:data<=16'd13520;
      47420:data<=16'd11050;
      47421:data<=16'd10035;
      47422:data<=16'd9862;
      47423:data<=16'd9467;
      47424:data<=16'd9667;
      47425:data<=16'd8786;
      47426:data<=16'd9618;
      47427:data<=16'd9609;
      47428:data<=16'd7837;
      47429:data<=16'd8525;
      47430:data<=16'd8035;
      47431:data<=16'd7138;
      47432:data<=16'd8122;
      47433:data<=16'd7997;
      47434:data<=16'd9592;
      47435:data<=16'd11295;
      47436:data<=16'd10361;
      47437:data<=16'd10414;
      47438:data<=16'd9749;
      47439:data<=16'd9814;
      47440:data<=16'd12087;
      47441:data<=16'd11371;
      47442:data<=16'd10298;
      47443:data<=16'd10543;
      47444:data<=16'd9967;
      47445:data<=16'd10843;
      47446:data<=16'd11665;
      47447:data<=16'd12145;
      47448:data<=16'd12222;
      47449:data<=16'd10539;
      47450:data<=16'd11239;
      47451:data<=16'd10786;
      47452:data<=16'd9530;
      47453:data<=16'd13670;
      47454:data<=16'd8881;
      47455:data<=-16'd4998;
      47456:data<=-16'd7257;
      47457:data<=-16'd4375;
      47458:data<=-16'd5391;
      47459:data<=-16'd3761;
      47460:data<=-16'd3024;
      47461:data<=-16'd3648;
      47462:data<=-16'd2358;
      47463:data<=-16'd2538;
      47464:data<=-16'd2575;
      47465:data<=-16'd1093;
      47466:data<=16'd208;
      47467:data<=-16'd441;
      47468:data<=-16'd4757;
      47469:data<=-16'd7027;
      47470:data<=-16'd5128;
      47471:data<=-16'd3841;
      47472:data<=-16'd2475;
      47473:data<=-16'd1565;
      47474:data<=-16'd1745;
      47475:data<=-16'd1328;
      47476:data<=-16'd2065;
      47477:data<=-16'd1562;
      47478:data<=16'd566;
      47479:data<=16'd458;
      47480:data<=16'd1192;
      47481:data<=16'd1818;
      47482:data<=16'd33;
      47483:data<=16'd1036;
      47484:data<=16'd3289;
      47485:data<=16'd3488;
      47486:data<=16'd3475;
      47487:data<=16'd2836;
      47488:data<=16'd2508;
      47489:data<=16'd3113;
      47490:data<=16'd4446;
      47491:data<=16'd6311;
      47492:data<=16'd5433;
      47493:data<=16'd5139;
      47494:data<=16'd6141;
      47495:data<=16'd3692;
      47496:data<=16'd9315;
      47497:data<=16'd23179;
      47498:data<=16'd24920;
      47499:data<=16'd20539;
      47500:data<=16'd22636;
      47501:data<=16'd22521;
      47502:data<=16'd21124;
      47503:data<=16'd22516;
      47504:data<=16'd21541;
      47505:data<=16'd20785;
      47506:data<=16'd20650;
      47507:data<=16'd18196;
      47508:data<=16'd17802;
      47509:data<=16'd18968;
      47510:data<=16'd18524;
      47511:data<=16'd18155;
      47512:data<=16'd17000;
      47513:data<=16'd15091;
      47514:data<=16'd15390;
      47515:data<=16'd16372;
      47516:data<=16'd15465;
      47517:data<=16'd15406;
      47518:data<=16'd18401;
      47519:data<=16'd20613;
      47520:data<=16'd20158;
      47521:data<=16'd19829;
      47522:data<=16'd19687;
      47523:data<=16'd19038;
      47524:data<=16'd18381;
      47525:data<=16'd17376;
      47526:data<=16'd16730;
      47527:data<=16'd16070;
      47528:data<=16'd15211;
      47529:data<=16'd14926;
      47530:data<=16'd13380;
      47531:data<=16'd12013;
      47532:data<=16'd12283;
      47533:data<=16'd10830;
      47534:data<=16'd8901;
      47535:data<=16'd7391;
      47536:data<=16'd6153;
      47537:data<=16'd7699;
      47538:data<=16'd3002;
      47539:data<=-16'd10428;
      47540:data<=-16'd15705;
      47541:data<=-16'd13074;
      47542:data<=-16'd14048;
      47543:data<=-16'd14774;
      47544:data<=-16'd14031;
      47545:data<=-16'd14869;
      47546:data<=-16'd15009;
      47547:data<=-16'd14921;
      47548:data<=-16'd14710;
      47549:data<=-16'd13975;
      47550:data<=-16'd13858;
      47551:data<=-16'd13312;
      47552:data<=-16'd13772;
      47553:data<=-16'd15195;
      47554:data<=-16'd14581;
      47555:data<=-16'd13976;
      47556:data<=-16'd13890;
      47557:data<=-16'd12924;
      47558:data<=-16'd13715;
      47559:data<=-16'd15324;
      47560:data<=-16'd14725;
      47561:data<=-16'd13979;
      47562:data<=-16'd14678;
      47563:data<=-16'd14425;
      47564:data<=-16'd13347;
      47565:data<=-16'd14248;
      47566:data<=-16'd14624;
      47567:data<=-16'd13885;
      47568:data<=-16'd17150;
      47569:data<=-16'd20299;
      47570:data<=-16'd18976;
      47571:data<=-16'd18971;
      47572:data<=-16'd19905;
      47573:data<=-16'd19183;
      47574:data<=-16'd19023;
      47575:data<=-16'd18004;
      47576:data<=-16'd16879;
      47577:data<=-16'd17179;
      47578:data<=-16'd17946;
      47579:data<=-16'd19238;
      47580:data<=-16'd13802;
      47581:data<=-16'd1303;
      47582:data<=16'd3350;
      47583:data<=16'd264;
      47584:data<=-16'd265;
      47585:data<=16'd77;
      47586:data<=-16'd152;
      47587:data<=16'd308;
      47588:data<=16'd173;
      47589:data<=-16'd190;
      47590:data<=-16'd1275;
      47591:data<=-16'd2485;
      47592:data<=-16'd2231;
      47593:data<=-16'd2093;
      47594:data<=-16'd1935;
      47595:data<=-16'd1351;
      47596:data<=-16'd2203;
      47597:data<=-16'd3419;
      47598:data<=-16'd3479;
      47599:data<=-16'd3642;
      47600:data<=-16'd3768;
      47601:data<=-16'd2760;
      47602:data<=-16'd2890;
      47603:data<=-16'd4767;
      47604:data<=-16'd4637;
      47605:data<=-16'd3859;
      47606:data<=-16'd4504;
      47607:data<=-16'd3465;
      47608:data<=-16'd3062;
      47609:data<=-16'd4552;
      47610:data<=-16'd4235;
      47611:data<=-16'd4511;
      47612:data<=-16'd4764;
      47613:data<=-16'd3051;
      47614:data<=-16'd3626;
      47615:data<=-16'd4291;
      47616:data<=-16'd4411;
      47617:data<=-16'd5609;
      47618:data<=-16'd2056;
      47619:data<=16'd1347;
      47620:data<=16'd535;
      47621:data<=16'd1911;
      47622:data<=-16'd3106;
      47623:data<=-16'd15120;
      47624:data<=-16'd18161;
      47625:data<=-16'd16460;
      47626:data<=-16'd17068;
      47627:data<=-16'd15461;
      47628:data<=-16'd14537;
      47629:data<=-16'd14543;
      47630:data<=-16'd13022;
      47631:data<=-16'd12624;
      47632:data<=-16'd12152;
      47633:data<=-16'd10895;
      47634:data<=-16'd9257;
      47635:data<=-16'd7275;
      47636:data<=-16'd7720;
      47637:data<=-16'd8287;
      47638:data<=-16'd6957;
      47639:data<=-16'd6302;
      47640:data<=-16'd4945;
      47641:data<=-16'd3286;
      47642:data<=-16'd3294;
      47643:data<=-16'd3275;
      47644:data<=-16'd3016;
      47645:data<=-16'd2479;
      47646:data<=-16'd1627;
      47647:data<=-16'd359;
      47648:data<=16'd1889;
      47649:data<=16'd2231;
      47650:data<=16'd1093;
      47651:data<=16'd1077;
      47652:data<=16'd1478;
      47653:data<=16'd3444;
      47654:data<=16'd4103;
      47655:data<=16'd2352;
      47656:data<=16'd3632;
      47657:data<=16'd3929;
      47658:data<=16'd3004;
      47659:data<=16'd6156;
      47660:data<=16'd6319;
      47661:data<=16'd5527;
      47662:data<=16'd7923;
      47663:data<=16'd5601;
      47664:data<=16'd8426;
      47665:data<=16'd21264;
      47666:data<=16'd26377;
      47667:data<=16'd24542;
      47668:data<=16'd22929;
      47669:data<=16'd18051;
      47670:data<=16'd15538;
      47671:data<=16'd17135;
      47672:data<=16'd17511;
      47673:data<=16'd17168;
      47674:data<=16'd16210;
      47675:data<=16'd15602;
      47676:data<=16'd15233;
      47677:data<=16'd14216;
      47678:data<=16'd15626;
      47679:data<=16'd16404;
      47680:data<=16'd14741;
      47681:data<=16'd14941;
      47682:data<=16'd14361;
      47683:data<=16'd13060;
      47684:data<=16'd14571;
      47685:data<=16'd14985;
      47686:data<=16'd13594;
      47687:data<=16'd13370;
      47688:data<=16'd13505;
      47689:data<=16'd12693;
      47690:data<=16'd11952;
      47691:data<=16'd13085;
      47692:data<=16'd12942;
      47693:data<=16'd11107;
      47694:data<=16'd12043;
      47695:data<=16'd11855;
      47696:data<=16'd10772;
      47697:data<=16'd12895;
      47698:data<=16'd11784;
      47699:data<=16'd9702;
      47700:data<=16'd10695;
      47701:data<=16'd8813;
      47702:data<=16'd8658;
      47703:data<=16'd10345;
      47704:data<=16'd8683;
      47705:data<=16'd10293;
      47706:data<=16'd7736;
      47707:data<=-16'd4502;
      47708:data<=-16'd9618;
      47709:data<=-16'd7168;
      47710:data<=-16'd6731;
      47711:data<=-16'd6396;
      47712:data<=-16'd6605;
      47713:data<=-16'd6921;
      47714:data<=-16'd6737;
      47715:data<=-16'd6243;
      47716:data<=-16'd3648;
      47717:data<=-16'd3688;
      47718:data<=-16'd3409;
      47719:data<=16'd1985;
      47720:data<=16'd2760;
      47721:data<=16'd1045;
      47722:data<=16'd3738;
      47723:data<=16'd4143;
      47724:data<=16'd3328;
      47725:data<=16'd3498;
      47726:data<=16'd2080;
      47727:data<=16'd2273;
      47728:data<=16'd2511;
      47729:data<=16'd1800;
      47730:data<=16'd2149;
      47731:data<=16'd1215;
      47732:data<=16'd1500;
      47733:data<=16'd2218;
      47734:data<=-16'd250;
      47735:data<=-16'd1201;
      47736:data<=-16'd1357;
      47737:data<=-16'd2546;
      47738:data<=-16'd1776;
      47739:data<=-16'd1601;
      47740:data<=-16'd2479;
      47741:data<=-16'd3703;
      47742:data<=-16'd5074;
      47743:data<=-16'd3774;
      47744:data<=-16'd3758;
      47745:data<=-16'd4502;
      47746:data<=-16'd3491;
      47747:data<=-16'd6977;
      47748:data<=-16'd5655;
      47749:data<=16'd6831;
      47750:data<=16'd12753;
      47751:data<=16'd10683;
      47752:data<=16'd10411;
      47753:data<=16'd8564;
      47754:data<=16'd6919;
      47755:data<=16'd7291;
      47756:data<=16'd6046;
      47757:data<=16'd5582;
      47758:data<=16'd5821;
      47759:data<=16'd4131;
      47760:data<=16'd2035;
      47761:data<=16'd1202;
      47762:data<=16'd1292;
      47763:data<=16'd957;
      47764:data<=16'd1102;
      47765:data<=16'd663;
      47766:data<=-16'd1776;
      47767:data<=-16'd1821;
      47768:data<=-16'd2435;
      47769:data<=-16'd7139;
      47770:data<=-16'd8369;
      47771:data<=-16'd7688;
      47772:data<=-16'd9547;
      47773:data<=-16'd9670;
      47774:data<=-16'd9879;
      47775:data<=-16'd10430;
      47776:data<=-16'd8987;
      47777:data<=-16'd9650;
      47778:data<=-16'd11150;
      47779:data<=-16'd11480;
      47780:data<=-16'd11837;
      47781:data<=-16'd10639;
      47782:data<=-16'd10060;
      47783:data<=-16'd9777;
      47784:data<=-16'd8994;
      47785:data<=-16'd11402;
      47786:data<=-16'd11882;
      47787:data<=-16'd10138;
      47788:data<=-16'd11391;
      47789:data<=-16'd9412;
      47790:data<=-16'd10331;
      47791:data<=-16'd22289;
      47792:data<=-16'd29141;
      47793:data<=-16'd26858;
      47794:data<=-16'd26786;
      47795:data<=-16'd26459;
      47796:data<=-16'd24773;
      47797:data<=-16'd25347;
      47798:data<=-16'd25410;
      47799:data<=-16'd24460;
      47800:data<=-16'd23802;
      47801:data<=-16'd22503;
      47802:data<=-16'd20777;
      47803:data<=-16'd20553;
      47804:data<=-16'd21880;
      47805:data<=-16'd20974;
      47806:data<=-16'd18506;
      47807:data<=-16'd18020;
      47808:data<=-16'd17294;
      47809:data<=-16'd16809;
      47810:data<=-16'd18346;
      47811:data<=-16'd17914;
      47812:data<=-16'd15891;
      47813:data<=-16'd15311;
      47814:data<=-16'd14766;
      47815:data<=-16'd14167;
      47816:data<=-16'd14856;
      47817:data<=-16'd15664;
      47818:data<=-16'd13101;
      47819:data<=-16'd7723;
      47820:data<=-16'd5664;
      47821:data<=-16'd6569;
      47822:data<=-16'd6557;
      47823:data<=-16'd6883;
      47824:data<=-16'd6740;
      47825:data<=-16'd5893;
      47826:data<=-16'd5777;
      47827:data<=-16'd4563;
      47828:data<=-16'd4090;
      47829:data<=-16'd4240;
      47830:data<=-16'd2270;
      47831:data<=-16'd2588;
      47832:data<=-16'd1260;
      47833:data<=16'd8405;
      47834:data<=16'd16128;
      47835:data<=16'd17191;
      47836:data<=16'd17553;
      47837:data<=16'd16442;
      47838:data<=16'd15449;
      47839:data<=16'd16298;
      47840:data<=16'd15960;
      47841:data<=16'd16624;
      47842:data<=16'd17581;
      47843:data<=16'd15916;
      47844:data<=16'd15414;
      47845:data<=16'd15873;
      47846:data<=16'd15371;
      47847:data<=16'd16020;
      47848:data<=16'd16186;
      47849:data<=16'd15393;
      47850:data<=16'd15764;
      47851:data<=16'd15565;
      47852:data<=16'd14744;
      47853:data<=16'd15120;
      47854:data<=16'd15502;
      47855:data<=16'd15308;
      47856:data<=16'd15323;
      47857:data<=16'd14789;
      47858:data<=16'd13491;
      47859:data<=16'd13556;
      47860:data<=16'd14766;
      47861:data<=16'd14475;
      47862:data<=16'd13870;
      47863:data<=16'd14351;
      47864:data<=16'd14327;
      47865:data<=16'd14096;
      47866:data<=16'd14466;
      47867:data<=16'd14939;
      47868:data<=16'd13571;
      47869:data<=16'd9385;
      47870:data<=16'd7027;
      47871:data<=16'd7065;
      47872:data<=16'd6493;
      47873:data<=16'd8743;
      47874:data<=16'd8821;
      47875:data<=-16'd187;
      47876:data<=-16'd7489;
      47877:data<=-16'd7718;
      47878:data<=-16'd6663;
      47879:data<=-16'd4353;
      47880:data<=-16'd3474;
      47881:data<=-16'd4808;
      47882:data<=-16'd3899;
      47883:data<=-16'd3577;
      47884:data<=-16'd3527;
      47885:data<=-16'd772;
      47886:data<=16'd168;
      47887:data<=-16'd717;
      47888:data<=-16'd745;
      47889:data<=-16'd826;
      47890:data<=16'd188;
      47891:data<=16'd1701;
      47892:data<=16'd2232;
      47893:data<=16'd2190;
      47894:data<=16'd1451;
      47895:data<=16'd1594;
      47896:data<=16'd2523;
      47897:data<=16'd3160;
      47898:data<=16'd4243;
      47899:data<=16'd3792;
      47900:data<=16'd2737;
      47901:data<=16'd3354;
      47902:data<=16'd3081;
      47903:data<=16'd3375;
      47904:data<=16'd4907;
      47905:data<=16'd4358;
      47906:data<=16'd4238;
      47907:data<=16'd4861;
      47908:data<=16'd4124;
      47909:data<=16'd4625;
      47910:data<=16'd5655;
      47911:data<=16'd6065;
      47912:data<=16'd6314;
      47913:data<=16'd5207;
      47914:data<=16'd5131;
      47915:data<=16'd5705;
      47916:data<=16'd6302;
      47917:data<=16'd13069;
      47918:data<=16'd22300;
      47919:data<=16'd25622;
      47920:data<=16'd26062;
      47921:data<=16'd26048;
      47922:data<=16'd25482;
      47923:data<=16'd25901;
      47924:data<=16'd25379;
      47925:data<=16'd23845;
      47926:data<=16'd22868;
      47927:data<=16'd21670;
      47928:data<=16'd20548;
      47929:data<=16'd19661;
      47930:data<=16'd19267;
      47931:data<=16'd18877;
      47932:data<=16'd16912;
      47933:data<=16'd15529;
      47934:data<=16'd14709;
      47935:data<=16'd12222;
      47936:data<=16'd10960;
      47937:data<=16'd10774;
      47938:data<=16'd9219;
      47939:data<=16'd8649;
      47940:data<=16'd8678;
      47941:data<=16'd7016;
      47942:data<=16'd5268;
      47943:data<=16'd4940;
      47944:data<=16'd5049;
      47945:data<=16'd4510;
      47946:data<=16'd4255;
      47947:data<=16'd3448;
      47948:data<=16'd1187;
      47949:data<=16'd1254;
      47950:data<=16'd2184;
      47951:data<=16'd761;
      47952:data<=16'd879;
      47953:data<=16'd382;
      47954:data<=-16'd2426;
      47955:data<=-16'd2162;
      47956:data<=-16'd2270;
      47957:data<=-16'd3124;
      47958:data<=-16'd1624;
      47959:data<=-16'd7750;
      47960:data<=-16'd18821;
      47961:data<=-16'd20633;
      47962:data<=-16'd18721;
      47963:data<=-16'd19443;
      47964:data<=-16'd18324;
      47965:data<=-16'd17379;
      47966:data<=-16'd18272;
      47967:data<=-16'd18142;
      47968:data<=-16'd18422;
      47969:data<=-16'd21100;
      47970:data<=-16'd23134;
      47971:data<=-16'd22325;
      47972:data<=-16'd22721;
      47973:data<=-16'd24225;
      47974:data<=-16'd22366;
      47975:data<=-16'd20897;
      47976:data<=-16'd21080;
      47977:data<=-16'd19315;
      47978:data<=-16'd19485;
      47979:data<=-16'd21080;
      47980:data<=-16'd19784;
      47981:data<=-16'd19106;
      47982:data<=-16'd19143;
      47983:data<=-16'd17999;
      47984:data<=-16'd18102;
      47985:data<=-16'd18609;
      47986:data<=-16'd18292;
      47987:data<=-16'd17579;
      47988:data<=-16'd16779;
      47989:data<=-16'd16500;
      47990:data<=-16'd15755;
      47991:data<=-16'd16164;
      47992:data<=-16'd17343;
      47993:data<=-16'd15676;
      47994:data<=-16'd15242;
      47995:data<=-16'd15835;
      47996:data<=-16'd13321;
      47997:data<=-16'd13594;
      47998:data<=-16'd14922;
      47999:data<=-16'd13491;
      48000:data<=-16'd14607;
      48001:data<=-16'd10099;
      48002:data<=16'd2029;
      48003:data<=16'd4790;
      48004:data<=16'd919;
      48005:data<=16'd1304;
      48006:data<=16'd1397;
      48007:data<=16'd1304;
      48008:data<=16'd2520;
      48009:data<=16'd1180;
      48010:data<=-16'd396;
      48011:data<=-16'd391;
      48012:data<=-16'd450;
      48013:data<=-16'd26;
      48014:data<=16'd285;
      48015:data<=-16'd426;
      48016:data<=-16'd1539;
      48017:data<=-16'd2511;
      48018:data<=-16'd2294;
      48019:data<=16'd196;
      48020:data<=16'd3656;
      48021:data<=16'd4783;
      48022:data<=16'd3530;
      48023:data<=16'd2541;
      48024:data<=16'd2338;
      48025:data<=16'd2870;
      48026:data<=16'd3168;
      48027:data<=16'd2520;
      48028:data<=16'd2602;
      48029:data<=16'd2734;
      48030:data<=16'd2905;
      48031:data<=16'd4141;
      48032:data<=16'd3927;
      48033:data<=16'd3445;
      48034:data<=16'd4002;
      48035:data<=16'd3723;
      48036:data<=16'd5133;
      48037:data<=16'd6246;
      48038:data<=16'd4670;
      48039:data<=16'd4943;
      48040:data<=16'd4035;
      48041:data<=16'd3313;
      48042:data<=16'd7661;
      48043:data<=16'd3792;
      48044:data<=-16'd8049;
      48045:data<=-16'd10225;
      48046:data<=-16'd7739;
      48047:data<=-16'd7902;
      48048:data<=-16'd5717;
      48049:data<=-16'd4666;
      48050:data<=-16'd5065;
      48051:data<=-16'd3532;
      48052:data<=-16'd3779;
      48053:data<=-16'd4118;
      48054:data<=-16'd2137;
      48055:data<=-16'd1333;
      48056:data<=-16'd1309;
      48057:data<=-16'd757;
      48058:data<=-16'd663;
      48059:data<=-16'd227;
      48060:data<=16'd1290;
      48061:data<=16'd2594;
      48062:data<=16'd2692;
      48063:data<=16'd2924;
      48064:data<=16'd3480;
      48065:data<=16'd3036;
      48066:data<=16'd2943;
      48067:data<=16'd4103;
      48068:data<=16'd5034;
      48069:data<=16'd3519;
      48070:data<=-16'd873;
      48071:data<=-16'd3357;
      48072:data<=-16'd2231;
      48073:data<=-16'd1105;
      48074:data<=-16'd89;
      48075:data<=16'd115;
      48076:data<=-16'd597;
      48077:data<=16'd325;
      48078:data<=16'd776;
      48079:data<=16'd1792;
      48080:data<=16'd4416;
      48081:data<=16'd3786;
      48082:data<=16'd3786;
      48083:data<=16'd4810;
      48084:data<=16'd2090;
      48085:data<=16'd7376;
      48086:data<=16'd19722;
      48087:data<=16'd21343;
      48088:data<=16'd18554;
      48089:data<=16'd19889;
      48090:data<=16'd18478;
      48091:data<=16'd17726;
      48092:data<=16'd19523;
      48093:data<=16'd18424;
      48094:data<=16'd17666;
      48095:data<=16'd17779;
      48096:data<=16'd15881;
      48097:data<=16'd15538;
      48098:data<=16'd17135;
      48099:data<=16'd17109;
      48100:data<=16'd15446;
      48101:data<=16'd13715;
      48102:data<=16'd12683;
      48103:data<=16'd12686;
      48104:data<=16'd13565;
      48105:data<=16'd13779;
      48106:data<=16'd12607;
      48107:data<=16'd11726;
      48108:data<=16'd11593;
      48109:data<=16'd11609;
      48110:data<=16'd11937;
      48111:data<=16'd12051;
      48112:data<=16'd11650;
      48113:data<=16'd11514;
      48114:data<=16'd11602;
      48115:data<=16'd10724;
      48116:data<=16'd10246;
      48117:data<=16'd11530;
      48118:data<=16'd10781;
      48119:data<=16'd10161;
      48120:data<=16'd14663;
      48121:data<=16'd16213;
      48122:data<=16'd13772;
      48123:data<=16'd15622;
      48124:data<=16'd15020;
      48125:data<=16'd12098;
      48126:data<=16'd14546;
      48127:data<=16'd10320;
      48128:data<=-16'd1202;
      48129:data<=-16'd4452;
      48130:data<=-16'd3565;
      48131:data<=-16'd4554;
      48132:data<=-16'd4099;
      48133:data<=-16'd4211;
      48134:data<=-16'd4322;
      48135:data<=-16'd4576;
      48136:data<=-16'd6986;
      48137:data<=-16'd7306;
      48138:data<=-16'd6633;
      48139:data<=-16'd7636;
      48140:data<=-16'd7092;
      48141:data<=-16'd6934;
      48142:data<=-16'd8354;
      48143:data<=-16'd8102;
      48144:data<=-16'd7841;
      48145:data<=-16'd8381;
      48146:data<=-16'd7709;
      48147:data<=-16'd7618;
      48148:data<=-16'd9233;
      48149:data<=-16'd9723;
      48150:data<=-16'd8842;
      48151:data<=-16'd9268;
      48152:data<=-16'd9470;
      48153:data<=-16'd8429;
      48154:data<=-16'd9430;
      48155:data<=-16'd10696;
      48156:data<=-16'd10116;
      48157:data<=-16'd10508;
      48158:data<=-16'd10525;
      48159:data<=-16'd9668;
      48160:data<=-16'd10481;
      48161:data<=-16'd10851;
      48162:data<=-16'd10780;
      48163:data<=-16'd11558;
      48164:data<=-16'd10786;
      48165:data<=-16'd9448;
      48166:data<=-16'd9274;
      48167:data<=-16'd10339;
      48168:data<=-16'd12110;
      48169:data<=-16'd9495;
      48170:data<=-16'd2878;
      48171:data<=-16'd132;
      48172:data<=-16'd1575;
      48173:data<=-16'd3154;
      48174:data<=-16'd3894;
      48175:data<=-16'd3553;
      48176:data<=-16'd3541;
      48177:data<=-16'd3873;
      48178:data<=-16'd3381;
      48179:data<=-16'd4114;
      48180:data<=-16'd5720;
      48181:data<=-16'd5870;
      48182:data<=-16'd5958;
      48183:data<=-16'd6049;
      48184:data<=-16'd5178;
      48185:data<=-16'd5809;
      48186:data<=-16'd7618;
      48187:data<=-16'd7536;
      48188:data<=-16'd6972;
      48189:data<=-16'd7080;
      48190:data<=-16'd6263;
      48191:data<=-16'd6382;
      48192:data<=-16'd8022;
      48193:data<=-16'd7958;
      48194:data<=-16'd7236;
      48195:data<=-16'd7379;
      48196:data<=-16'd6863;
      48197:data<=-16'd7157;
      48198:data<=-16'd8443;
      48199:data<=-16'd8343;
      48200:data<=-16'd7905;
      48201:data<=-16'd7674;
      48202:data<=-16'd7470;
      48203:data<=-16'd8031;
      48204:data<=-16'd7806;
      48205:data<=-16'd7865;
      48206:data<=-16'd9233;
      48207:data<=-16'd8807;
      48208:data<=-16'd8481;
      48209:data<=-16'd8490;
      48210:data<=-16'd6476;
      48211:data<=-16'd11235;
      48212:data<=-16'd22254;
      48213:data<=-16'd24662;
      48214:data<=-16'd21635;
      48215:data<=-16'd22128;
      48216:data<=-16'd21664;
      48217:data<=-16'd21100;
      48218:data<=-16'd21877;
      48219:data<=-16'd18724;
      48220:data<=-16'd14060;
      48221:data<=-16'd11896;
      48222:data<=-16'd11467;
      48223:data<=-16'd12038;
      48224:data<=-16'd11482;
      48225:data<=-16'd10554;
      48226:data<=-16'd10751;
      48227:data<=-16'd9824;
      48228:data<=-16'd9069;
      48229:data<=-16'd9376;
      48230:data<=-16'd8334;
      48231:data<=-16'd7462;
      48232:data<=-16'd7363;
      48233:data<=-16'd6583;
      48234:data<=-16'd6387;
      48235:data<=-16'd6108;
      48236:data<=-16'd4275;
      48237:data<=-16'd2605;
      48238:data<=-16'd1968;
      48239:data<=-16'd1762;
      48240:data<=-16'd2411;
      48241:data<=-16'd2740;
      48242:data<=-16'd664;
      48243:data<=16'd999;
      48244:data<=16'd467;
      48245:data<=16'd905;
      48246:data<=16'd763;
      48247:data<=16'd168;
      48248:data<=16'd3287;
      48249:data<=16'd5142;
      48250:data<=16'd4455;
      48251:data<=16'd5257;
      48252:data<=16'd3671;
      48253:data<=16'd6178;
      48254:data<=16'd17885;
      48255:data<=16'd23071;
      48256:data<=16'd20509;
      48257:data<=16'd20985;
      48258:data<=16'd20199;
      48259:data<=16'd18393;
      48260:data<=16'd19572;
      48261:data<=16'd19889;
      48262:data<=16'd19886;
      48263:data<=16'd19726;
      48264:data<=16'd18434;
      48265:data<=16'd18465;
      48266:data<=16'd18174;
      48267:data<=16'd18014;
      48268:data<=16'd19249;
      48269:data<=16'd17123;
      48270:data<=16'd12392;
      48271:data<=16'd9703;
      48272:data<=16'd9186;
      48273:data<=16'd10125;
      48274:data<=16'd10903;
      48275:data<=16'd10434;
      48276:data<=16'd10107;
      48277:data<=16'd9946;
      48278:data<=16'd8992;
      48279:data<=16'd8846;
      48280:data<=16'd10988;
      48281:data<=16'd11831;
      48282:data<=16'd10307;
      48283:data<=16'd10340;
      48284:data<=16'd10178;
      48285:data<=16'd9609;
      48286:data<=16'd11552;
      48287:data<=16'd11609;
      48288:data<=16'd10475;
      48289:data<=16'd11209;
      48290:data<=16'd9777;
      48291:data<=16'd9219;
      48292:data<=16'd10586;
      48293:data<=16'd9903;
      48294:data<=16'd10784;
      48295:data<=16'd7821;
      48296:data<=-16'd2523;
      48297:data<=-16'd6783;
      48298:data<=-16'd4701;
      48299:data<=-16'd4414;
      48300:data<=-16'd3852;
      48301:data<=-16'd3782;
      48302:data<=-16'd4156;
      48303:data<=-16'd3224;
      48304:data<=-16'd2883;
      48305:data<=-16'd1521;
      48306:data<=-16'd387;
      48307:data<=-16'd1400;
      48308:data<=-16'd1143;
      48309:data<=-16'd500;
      48310:data<=-16'd21;
      48311:data<=16'd1271;
      48312:data<=16'd980;
      48313:data<=16'd863;
      48314:data<=16'd1574;
      48315:data<=16'd905;
      48316:data<=16'd1289;
      48317:data<=16'd2564;
      48318:data<=16'd2273;
      48319:data<=16'd2476;
      48320:data<=16'd5517;
      48321:data<=16'd9065;
      48322:data<=16'd9298;
      48323:data<=16'd9145;
      48324:data<=16'd10625;
      48325:data<=16'd9491;
      48326:data<=16'd8317;
      48327:data<=16'd9054;
      48328:data<=16'd8155;
      48329:data<=16'd7991;
      48330:data<=16'd7714;
      48331:data<=16'd6009;
      48332:data<=16'd6839;
      48333:data<=16'd6830;
      48334:data<=16'd6169;
      48335:data<=16'd6924;
      48336:data<=16'd3664;
      48337:data<=16'd4793;
      48338:data<=16'd15010;
      48339:data<=16'd18832;
      48340:data<=16'd16456;
      48341:data<=16'd16512;
      48342:data<=16'd14549;
      48343:data<=16'd12003;
      48344:data<=16'd12094;
      48345:data<=16'd11232;
      48346:data<=16'd10367;
      48347:data<=16'd10607;
      48348:data<=16'd9670;
      48349:data<=16'd7871;
      48350:data<=16'd7083;
      48351:data<=16'd6986;
      48352:data<=16'd6173;
      48353:data<=16'd5870;
      48354:data<=16'd5526;
      48355:data<=16'd3183;
      48356:data<=16'd1906;
      48357:data<=16'd2052;
      48358:data<=16'd1328;
      48359:data<=16'd1354;
      48360:data<=16'd846;
      48361:data<=-16'd911;
      48362:data<=-16'd1404;
      48363:data<=-16'd2047;
      48364:data<=-16'd2808;
      48365:data<=-16'd2246;
      48366:data<=-16'd2144;
      48367:data<=-16'd2933;
      48368:data<=-16'd3707;
      48369:data<=-16'd3817;
      48370:data<=-16'd5670;
      48371:data<=-16'd10140;
      48372:data<=-16'd10721;
      48373:data<=-16'd9777;
      48374:data<=-16'd12833;
      48375:data<=-16'd12775;
      48376:data<=-16'd11317;
      48377:data<=-16'd12690;
      48378:data<=-16'd10381;
      48379:data<=-16'd12696;
      48380:data<=-16'd24168;
      48381:data<=-16'd28688;
      48382:data<=-16'd26598;
      48383:data<=-16'd26708;
      48384:data<=-16'd25417;
      48385:data<=-16'd24213;
      48386:data<=-16'd24871;
      48387:data<=-16'd24159;
      48388:data<=-16'd23469;
      48389:data<=-16'd22908;
      48390:data<=-16'd21488;
      48391:data<=-16'd20442;
      48392:data<=-16'd20237;
      48393:data<=-16'd20809;
      48394:data<=-16'd20389;
      48395:data<=-16'd19505;
      48396:data<=-16'd19517;
      48397:data<=-16'd18180;
      48398:data<=-16'd17449;
      48399:data<=-16'd18483;
      48400:data<=-16'd17775;
      48401:data<=-16'd16960;
      48402:data<=-16'd16375;
      48403:data<=-16'd14737;
      48404:data<=-16'd14913;
      48405:data<=-16'd15191;
      48406:data<=-16'd14261;
      48407:data<=-16'd14324;
      48408:data<=-16'd13769;
      48409:data<=-16'd12997;
      48410:data<=-16'd12774;
      48411:data<=-16'd12192;
      48412:data<=-16'd12754;
      48413:data<=-16'd12533;
      48414:data<=-16'd11145;
      48415:data<=-16'd11130;
      48416:data<=-16'd10375;
      48417:data<=-16'd10084;
      48418:data<=-16'd11092;
      48419:data<=-16'd10260;
      48420:data<=-16'd8486;
      48421:data<=-16'd1964;
      48422:data<=16'd9045;
      48423:data<=16'd12683;
      48424:data<=16'd10780;
      48425:data<=16'd11162;
      48426:data<=16'd10712;
      48427:data<=16'd10132;
      48428:data<=16'd10725;
      48429:data<=16'd10011;
      48430:data<=16'd9632;
      48431:data<=16'd9404;
      48432:data<=16'd8859;
      48433:data<=16'd9432;
      48434:data<=16'd9611;
      48435:data<=16'd9385;
      48436:data<=16'd9488;
      48437:data<=16'd9617;
      48438:data<=16'd10251;
      48439:data<=16'd10329;
      48440:data<=16'd9699;
      48441:data<=16'd8842;
      48442:data<=16'd8320;
      48443:data<=16'd9706;
      48444:data<=16'd10399;
      48445:data<=16'd9696;
      48446:data<=16'd10073;
      48447:data<=16'd9212;
      48448:data<=16'd8655;
      48449:data<=16'd10533;
      48450:data<=16'd10660;
      48451:data<=16'd10308;
      48452:data<=16'd10561;
      48453:data<=16'd9406;
      48454:data<=16'd9834;
      48455:data<=16'd10887;
      48456:data<=16'd10936;
      48457:data<=16'd11681;
      48458:data<=16'd10836;
      48459:data<=16'd9688;
      48460:data<=16'd9498;
      48461:data<=16'd8960;
      48462:data<=16'd11201;
      48463:data<=16'd9802;
      48464:data<=-16'd33;
      48465:data<=-16'd5418;
      48466:data<=-16'd4184;
      48467:data<=-16'd3973;
      48468:data<=-16'd2397;
      48469:data<=-16'd1007;
      48470:data<=-16'd3806;
      48471:data<=-16'd7542;
      48472:data<=-16'd9109;
      48473:data<=-16'd7412;
      48474:data<=-16'd5228;
      48475:data<=-16'd5268;
      48476:data<=-16'd4927;
      48477:data<=-16'd4366;
      48478:data<=-16'd4540;
      48479:data<=-16'd3421;
      48480:data<=-16'd1817;
      48481:data<=-16'd939;
      48482:data<=-16'd576;
      48483:data<=-16'd538;
      48484:data<=-16'd455;
      48485:data<=-16'd569;
      48486:data<=16'd707;
      48487:data<=16'd2951;
      48488:data<=16'd2826;
      48489:data<=16'd2419;
      48490:data<=16'd3234;
      48491:data<=16'd3206;
      48492:data<=16'd3935;
      48493:data<=16'd5034;
      48494:data<=16'd4551;
      48495:data<=16'd4234;
      48496:data<=16'd4129;
      48497:data<=16'd3891;
      48498:data<=16'd4138;
      48499:data<=16'd4593;
      48500:data<=16'd5582;
      48501:data<=16'd5488;
      48502:data<=16'd5084;
      48503:data<=16'd6391;
      48504:data<=16'd5591;
      48505:data<=16'd6722;
      48506:data<=16'd15609;
      48507:data<=16'd21490;
      48508:data<=16'd20398;
      48509:data<=16'd20280;
      48510:data<=16'd19415;
      48511:data<=16'd18208;
      48512:data<=16'd19795;
      48513:data<=16'd19146;
      48514:data<=16'd17719;
      48515:data<=16'd18036;
      48516:data<=16'd16163;
      48517:data<=16'd15588;
      48518:data<=16'd17152;
      48519:data<=16'd15841;
      48520:data<=16'd16427;
      48521:data<=16'd20489;
      48522:data<=16'd21109;
      48523:data<=16'd19890;
      48524:data<=16'd20527;
      48525:data<=16'd20177;
      48526:data<=16'd18751;
      48527:data<=16'd18148;
      48528:data<=16'd16933;
      48529:data<=16'd15245;
      48530:data<=16'd14686;
      48531:data<=16'd13893;
      48532:data<=16'd12574;
      48533:data<=16'd11972;
      48534:data<=16'd11097;
      48535:data<=16'd10190;
      48536:data<=16'd9307;
      48537:data<=16'd7172;
      48538:data<=16'd6050;
      48539:data<=16'd6088;
      48540:data<=16'd5444;
      48541:data<=16'd5495;
      48542:data<=16'd4235;
      48543:data<=16'd1720;
      48544:data<=16'd1618;
      48545:data<=16'd876;
      48546:data<=-16'd62;
      48547:data<=-16'd591;
      48548:data<=-16'd8328;
      48549:data<=-16'd17212;
      48550:data<=-16'd17441;
      48551:data<=-16'd16264;
      48552:data<=-16'd16625;
      48553:data<=-16'd15561;
      48554:data<=-16'd15622;
      48555:data<=-16'd16035;
      48556:data<=-16'd16296;
      48557:data<=-16'd16782;
      48558:data<=-16'd15706;
      48559:data<=-16'd15299;
      48560:data<=-16'd15553;
      48561:data<=-16'd15346;
      48562:data<=-16'd16349;
      48563:data<=-16'd16035;
      48564:data<=-16'd15180;
      48565:data<=-16'd15793;
      48566:data<=-16'd14266;
      48567:data<=-16'd13543;
      48568:data<=-16'd15130;
      48569:data<=-16'd14286;
      48570:data<=-16'd15232;
      48571:data<=-16'd19332;
      48572:data<=-16'd19928;
      48573:data<=-16'd18735;
      48574:data<=-16'd19314;
      48575:data<=-16'd19623;
      48576:data<=-16'd19005;
      48577:data<=-16'd18507;
      48578:data<=-16'd17743;
      48579:data<=-16'd16419;
      48580:data<=-16'd16860;
      48581:data<=-16'd18503;
      48582:data<=-16'd18266;
      48583:data<=-16'd18002;
      48584:data<=-16'd17221;
      48585:data<=-16'd15124;
      48586:data<=-16'd15863;
      48587:data<=-16'd16315;
      48588:data<=-16'd15123;
      48589:data<=-16'd15026;
      48590:data<=-16'd8237;
      48591:data<=16'd1656;
      48592:data<=16'd1986;
      48593:data<=-16'd367;
      48594:data<=-16'd220;
      48595:data<=-16'd1518;
      48596:data<=-16'd910;
      48597:data<=16'd265;
      48598:data<=-16'd644;
      48599:data<=-16'd1178;
      48600:data<=-16'd2619;
      48601:data<=-16'd3295;
      48602:data<=-16'd2226;
      48603:data<=-16'd2435;
      48604:data<=-16'd2241;
      48605:data<=-16'd2717;
      48606:data<=-16'd4475;
      48607:data<=-16'd3817;
      48608:data<=-16'd3630;
      48609:data<=-16'd4370;
      48610:data<=-16'd3224;
      48611:data<=-16'd3733;
      48612:data<=-16'd5503;
      48613:data<=-16'd5680;
      48614:data<=-16'd5573;
      48615:data<=-16'd5309;
      48616:data<=-16'd5180;
      48617:data<=-16'd5368;
      48618:data<=-16'd6056;
      48619:data<=-16'd7201;
      48620:data<=-16'd5177;
      48621:data<=-16'd1017;
      48622:data<=16'd930;
      48623:data<=16'd1139;
      48624:data<=16'd215;
      48625:data<=-16'd529;
      48626:data<=-16'd796;
      48627:data<=-16'd1532;
      48628:data<=-16'd378;
      48629:data<=-16'd227;
      48630:data<=-16'd1606;
      48631:data<=-16'd494;
      48632:data<=-16'd5470;
      48633:data<=-16'd15250;
      48634:data<=-16'd15908;
      48635:data<=-16'd13714;
      48636:data<=-16'd14116;
      48637:data<=-16'd11276;
      48638:data<=-16'd10184;
      48639:data<=-16'd11007;
      48640:data<=-16'd9263;
      48641:data<=-16'd8975;
      48642:data<=-16'd8513;
      48643:data<=-16'd6188;
      48644:data<=-16'd5465;
      48645:data<=-16'd4749;
      48646:data<=-16'd3627;
      48647:data<=-16'd3532;
      48648:data<=-16'd3659;
      48649:data<=-16'd3086;
      48650:data<=-16'd1098;
      48651:data<=-16'd106;
      48652:data<=-16'd268;
      48653:data<=16'd651;
      48654:data<=16'd528;
      48655:data<=16'd1087;
      48656:data<=16'd3673;
      48657:data<=16'd3903;
      48658:data<=16'd3418;
      48659:data<=16'd3738;
      48660:data<=16'd3096;
      48661:data<=16'd3817;
      48662:data<=16'd5406;
      48663:data<=16'd6185;
      48664:data<=16'd6454;
      48665:data<=16'd5818;
      48666:data<=16'd5956;
      48667:data<=16'd6097;
      48668:data<=16'd6525;
      48669:data<=16'd8671;
      48670:data<=16'd6969;
      48671:data<=16'd3395;
      48672:data<=16'd2309;
      48673:data<=16'd343;
      48674:data<=16'd5600;
      48675:data<=16'd17673;
      48676:data<=16'd19973;
      48677:data<=16'd17500;
      48678:data<=16'd18101;
      48679:data<=16'd16175;
      48680:data<=16'd16571;
      48681:data<=16'd19306;
      48682:data<=16'd18283;
      48683:data<=16'd17898;
      48684:data<=16'd17246;
      48685:data<=16'd14945;
      48686:data<=16'd15814;
      48687:data<=16'd16976;
      48688:data<=16'd16242;
      48689:data<=16'd15896;
      48690:data<=16'd15608;
      48691:data<=16'd15288;
      48692:data<=16'd14590;
      48693:data<=16'd14692;
      48694:data<=16'd15717;
      48695:data<=16'd14681;
      48696:data<=16'd13661;
      48697:data<=16'd13376;
      48698:data<=16'd11568;
      48699:data<=16'd11568;
      48700:data<=16'd13138;
      48701:data<=16'd12743;
      48702:data<=16'd11712;
      48703:data<=16'd10866;
      48704:data<=16'd10448;
      48705:data<=16'd10615;
      48706:data<=16'd10763;
      48707:data<=16'd11383;
      48708:data<=16'd11197;
      48709:data<=16'd10361;
      48710:data<=16'd9859;
      48711:data<=16'd9212;
      48712:data<=16'd10443;
      48713:data<=16'd10564;
      48714:data<=16'd8395;
      48715:data<=16'd9545;
      48716:data<=16'd5541;
      48717:data<=-16'd5823;
      48718:data<=-16'd7447;
      48719:data<=-16'd3679;
      48720:data<=-16'd4965;
      48721:data<=-16'd1809;
      48722:data<=16'd2689;
      48723:data<=16'd1180;
      48724:data<=16'd1407;
      48725:data<=16'd3240;
      48726:data<=16'd3007;
      48727:data<=16'd3316;
      48728:data<=16'd3027;
      48729:data<=16'd2049;
      48730:data<=16'd2052;
      48731:data<=16'd2193;
      48732:data<=16'd2115;
      48733:data<=16'd1444;
      48734:data<=16'd1180;
      48735:data<=16'd1533;
      48736:data<=16'd473;
      48737:data<=-16'd760;
      48738:data<=-16'd920;
      48739:data<=-16'd926;
      48740:data<=-16'd939;
      48741:data<=-16'd1107;
      48742:data<=-16'd925;
      48743:data<=-16'd1457;
      48744:data<=-16'd3021;
      48745:data<=-16'd2911;
      48746:data<=-16'd2773;
      48747:data<=-16'd3413;
      48748:data<=-16'd2660;
      48749:data<=-16'd3315;
      48750:data<=-16'd4974;
      48751:data<=-16'd4892;
      48752:data<=-16'd4784;
      48753:data<=-16'd4534;
      48754:data<=-16'd4757;
      48755:data<=-16'd5136;
      48756:data<=-16'd5033;
      48757:data<=-16'd7413;
      48758:data<=-16'd4241;
      48759:data<=16'd6933;
      48760:data<=16'd10232;
      48761:data<=16'd7344;
      48762:data<=16'd7266;
      48763:data<=16'd5285;
      48764:data<=16'd4895;
      48765:data<=16'd6379;
      48766:data<=16'd4772;
      48767:data<=16'd5377;
      48768:data<=16'd4490;
      48769:data<=16'd1061;
      48770:data<=16'd2707;
      48771:data<=16'd734;
      48772:data<=-16'd5500;
      48773:data<=-16'd5363;
      48774:data<=-16'd4977;
      48775:data<=-16'd6916;
      48776:data<=-16'd6678;
      48777:data<=-16'd7260;
      48778:data<=-16'd7530;
      48779:data<=-16'd6387;
      48780:data<=-16'd6893;
      48781:data<=-16'd8310;
      48782:data<=-16'd9356;
      48783:data<=-16'd9424;
      48784:data<=-16'd9034;
      48785:data<=-16'd8663;
      48786:data<=-16'd8073;
      48787:data<=-16'd9230;
      48788:data<=-16'd10263;
      48789:data<=-16'd9652;
      48790:data<=-16'd10249;
      48791:data<=-16'd9985;
      48792:data<=-16'd8693;
      48793:data<=-16'd9247;
      48794:data<=-16'd9969;
      48795:data<=-16'd10436;
      48796:data<=-16'd9999;
      48797:data<=-16'd9198;
      48798:data<=-16'd9250;
      48799:data<=-16'd8067;
      48800:data<=-16'd12871;
      48801:data<=-16'd24184;
      48802:data<=-16'd26697;
      48803:data<=-16'd23220;
      48804:data<=-16'd22782;
      48805:data<=-16'd21720;
      48806:data<=-16'd22391;
      48807:data<=-16'd23376;
      48808:data<=-16'd20999;
      48809:data<=-16'd20609;
      48810:data<=-16'd19867;
      48811:data<=-16'd18167;
      48812:data<=-16'd19839;
      48813:data<=-16'd19886;
      48814:data<=-16'd18254;
      48815:data<=-16'd17755;
      48816:data<=-16'd16589;
      48817:data<=-16'd16672;
      48818:data<=-16'd16627;
      48819:data<=-16'd15823;
      48820:data<=-16'd16160;
      48821:data<=-16'd13000;
      48822:data<=-16'd7793;
      48823:data<=-16'd6091;
      48824:data<=-16'd6540;
      48825:data<=-16'd7392;
      48826:data<=-16'd6893;
      48827:data<=-16'd5977;
      48828:data<=-16'd6167;
      48829:data<=-16'd5080;
      48830:data<=-16'd4878;
      48831:data<=-16'd5260;
      48832:data<=-16'd3280;
      48833:data<=-16'd2620;
      48834:data<=-16'd2649;
      48835:data<=-16'd2332;
      48836:data<=-16'd2927;
      48837:data<=-16'd980;
      48838:data<=16'd490;
      48839:data<=16'd537;
      48840:data<=16'd2179;
      48841:data<=16'd749;
      48842:data<=16'd3648;
      48843:data<=16'd15370;
      48844:data<=16'd19760;
      48845:data<=16'd17482;
      48846:data<=16'd18245;
      48847:data<=16'd17522;
      48848:data<=16'd16466;
      48849:data<=16'd17290;
      48850:data<=16'd17685;
      48851:data<=16'd18674;
      48852:data<=16'd18172;
      48853:data<=16'd17070;
      48854:data<=16'd17252;
      48855:data<=16'd16130;
      48856:data<=16'd16308;
      48857:data<=16'd17236;
      48858:data<=16'd15881;
      48859:data<=16'd15810;
      48860:data<=16'd15826;
      48861:data<=16'd14504;
      48862:data<=16'd14965;
      48863:data<=16'd15637;
      48864:data<=16'd15578;
      48865:data<=16'd15264;
      48866:data<=16'd14443;
      48867:data<=16'd14220;
      48868:data<=16'd13585;
      48869:data<=16'd13744;
      48870:data<=16'd14812;
      48871:data<=16'd11931;
      48872:data<=16'd7324;
      48873:data<=16'd5277;
      48874:data<=16'd4960;
      48875:data<=16'd6018;
      48876:data<=16'd6634;
      48877:data<=16'd6610;
      48878:data<=16'd6498;
      48879:data<=16'd5066;
      48880:data<=16'd5556;
      48881:data<=16'd6953;
      48882:data<=16'd6771;
      48883:data<=16'd8381;
      48884:data<=16'd5159;
      48885:data<=-16'd5210;
      48886:data<=-16'd9333;
      48887:data<=-16'd7004;
      48888:data<=-16'd5927;
      48889:data<=-16'd5166;
      48890:data<=-16'd5133;
      48891:data<=-16'd5538;
      48892:data<=-16'd5541;
      48893:data<=-16'd5359;
      48894:data<=-16'd2846;
      48895:data<=-16'd1283;
      48896:data<=-16'd2196;
      48897:data<=-16'd1729;
      48898:data<=-16'd1779;
      48899:data<=-16'd1559;
      48900:data<=16'd673;
      48901:data<=16'd543;
      48902:data<=-16'd206;
      48903:data<=16'd720;
      48904:data<=16'd688;
      48905:data<=16'd926;
      48906:data<=16'd1991;
      48907:data<=16'd2875;
      48908:data<=16'd3415;
      48909:data<=16'd3309;
      48910:data<=16'd3779;
      48911:data<=16'd3368;
      48912:data<=16'd2817;
      48913:data<=16'd4840;
      48914:data<=16'd4937;
      48915:data<=16'd4059;
      48916:data<=16'd5394;
      48917:data<=16'd4358;
      48918:data<=16'd4235;
      48919:data<=16'd6334;
      48920:data<=16'd5456;
      48921:data<=16'd7189;
      48922:data<=16'd11520;
      48923:data<=16'd12545;
      48924:data<=16'd12598;
      48925:data<=16'd11552;
      48926:data<=16'd14926;
      48927:data<=16'd25332;
      48928:data<=16'd28433;
      48929:data<=16'd24943;
      48930:data<=16'd24859;
      48931:data<=16'd23711;
      48932:data<=16'd22063;
      48933:data<=16'd22075;
      48934:data<=16'd20359;
      48935:data<=16'd19444;
      48936:data<=16'd18965;
      48937:data<=16'd16994;
      48938:data<=16'd15444;
      48939:data<=16'd13687;
      48940:data<=16'd12331;
      48941:data<=16'd11621;
      48942:data<=16'd11062;
      48943:data<=16'd10957;
      48944:data<=16'd8605;
      48945:data<=16'd6419;
      48946:data<=16'd6661;
      48947:data<=16'd5618;
      48948:data<=16'd5451;
      48949:data<=16'd5535;
      48950:data<=16'd2787;
      48951:data<=16'd1844;
      48952:data<=16'd1704;
      48953:data<=16'd482;
      48954:data<=16'd854;
      48955:data<=16'd255;
      48956:data<=-16'd984;
      48957:data<=-16'd1735;
      48958:data<=-16'd3331;
      48959:data<=-16'd3626;
      48960:data<=-16'd3973;
      48961:data<=-16'd4000;
      48962:data<=-16'd3278;
      48963:data<=-16'd5838;
      48964:data<=-16'd6567;
      48965:data<=-16'd5718;
      48966:data<=-16'd7464;
      48967:data<=-16'd4819;
      48968:data<=-16'd7156;
      48969:data<=-16'd20181;
      48970:data<=-16'd24184;
      48971:data<=-16'd22333;
      48972:data<=-16'd26814;
      48973:data<=-16'd27940;
      48974:data<=-16'd26295;
      48975:data<=-16'd27640;
      48976:data<=-16'd27869;
      48977:data<=-16'd26982;
      48978:data<=-16'd25819;
      48979:data<=-16'd24927;
      48980:data<=-16'd24400;
      48981:data<=-16'd23346;
      48982:data<=-16'd23883;
      48983:data<=-16'd23682;
      48984:data<=-16'd22380;
      48985:data<=-16'd22606;
      48986:data<=-16'd20647;
      48987:data<=-16'd19405;
      48988:data<=-16'd21276;
      48989:data<=-16'd20313;
      48990:data<=-16'd19115;
      48991:data<=-16'd18856;
      48992:data<=-16'd16832;
      48993:data<=-16'd16941;
      48994:data<=-16'd17622;
      48995:data<=-16'd16813;
      48996:data<=-16'd16550;
      48997:data<=-16'd15376;
      48998:data<=-16'd14545;
      48999:data<=-16'd14129;
      49000:data<=-16'd13711;
      49001:data<=-16'd15215;
      49002:data<=-16'd14636;
      49003:data<=-16'd13138;
      49004:data<=-16'd13537;
      49005:data<=-16'd11768;
      49006:data<=-16'd11696;
      49007:data<=-16'd13076;
      49008:data<=-16'd11620;
      49009:data<=-16'd12797;
      49010:data<=-16'd9580;
      49011:data<=16'd1953;
      49012:data<=16'd5655;
      49013:data<=16'd2781;
      49014:data<=16'd3203;
      49015:data<=16'd2732;
      49016:data<=16'd2021;
      49017:data<=16'd2860;
      49018:data<=16'd2605;
      49019:data<=16'd1800;
      49020:data<=16'd338;
      49021:data<=16'd825;
      49022:data<=16'd4637;
      49023:data<=16'd6905;
      49024:data<=16'd6646;
      49025:data<=16'd5360;
      49026:data<=16'd4141;
      49027:data<=16'd4410;
      49028:data<=16'd4353;
      49029:data<=16'd3918;
      49030:data<=16'd3971;
      49031:data<=16'd3294;
      49032:data<=16'd3278;
      49033:data<=16'd3877;
      49034:data<=16'd3600;
      49035:data<=16'd3169;
      49036:data<=16'd2300;
      49037:data<=16'd2396;
      49038:data<=16'd4161;
      49039:data<=16'd4437;
      49040:data<=16'd3609;
      49041:data<=16'd3404;
      49042:data<=16'd3093;
      49043:data<=16'd3245;
      49044:data<=16'd4387;
      49045:data<=16'd5513;
      49046:data<=16'd5078;
      49047:data<=16'd4258;
      49048:data<=16'd4952;
      49049:data<=16'd4027;
      49050:data<=16'd3598;
      49051:data<=16'd7464;
      49052:data<=16'd5115;
      49053:data<=-16'd5426;
      49054:data<=-16'd10003;
      49055:data<=-16'd8943;
      49056:data<=-16'd8558;
      49057:data<=-16'd6064;
      49058:data<=-16'd4325;
      49059:data<=-16'd5418;
      49060:data<=-16'd5225;
      49061:data<=-16'd4554;
      49062:data<=-16'd3718;
      49063:data<=-16'd1779;
      49064:data<=-16'd999;
      49065:data<=-16'd1051;
      49066:data<=-16'd1039;
      49067:data<=-16'd889;
      49068:data<=16'd165;
      49069:data<=16'd1022;
      49070:data<=16'd1744;
      49071:data<=16'd1533;
      49072:data<=-16'd1469;
      49073:data<=-16'd4047;
      49074:data<=-16'd4608;
      49075:data<=-16'd4003;
      49076:data<=-16'd1826;
      49077:data<=-16'd1257;
      49078:data<=-16'd1742;
      49079:data<=-16'd497;
      49080:data<=-16'd701;
      49081:data<=-16'd259;
      49082:data<=16'd2836;
      49083:data<=16'd3338;
      49084:data<=16'd2802;
      49085:data<=16'd3574;
      49086:data<=16'd3263;
      49087:data<=16'd3755;
      49088:data<=16'd5341;
      49089:data<=16'd5733;
      49090:data<=16'd5454;
      49091:data<=16'd5841;
      49092:data<=16'd6112;
      49093:data<=16'd4074;
      49094:data<=16'd6680;
      49095:data<=16'd17832;
      49096:data<=16'd23156;
      49097:data<=16'd20447;
      49098:data<=16'd20292;
      49099:data<=16'd19434;
      49100:data<=16'd18463;
      49101:data<=16'd20662;
      49102:data<=16'd19725;
      49103:data<=16'd18043;
      49104:data<=16'd18093;
      49105:data<=16'd16377;
      49106:data<=16'd16189;
      49107:data<=16'd17230;
      49108:data<=16'd16913;
      49109:data<=16'd16384;
      49110:data<=16'd14936;
      49111:data<=16'd14460;
      49112:data<=16'd14859;
      49113:data<=16'd14483;
      49114:data<=16'd14866;
      49115:data<=16'd13418;
      49116:data<=16'd12196;
      49117:data<=16'd13740;
      49118:data<=16'd12128;
      49119:data<=16'd11268;
      49120:data<=16'd13524;
      49121:data<=16'd11999;
      49122:data<=16'd12478;
      49123:data<=16'd16839;
      49124:data<=16'd16829;
      49125:data<=16'd15615;
      49126:data<=16'd16254;
      49127:data<=16'd15861;
      49128:data<=16'd14922;
      49129:data<=16'd14004;
      49130:data<=16'd13537;
      49131:data<=16'd12834;
      49132:data<=16'd11400;
      49133:data<=16'd10319;
      49134:data<=16'd9632;
      49135:data<=16'd10753;
      49136:data<=16'd8668;
      49137:data<=-16'd1804;
      49138:data<=-16'd9746;
      49139:data<=-16'd9759;
      49140:data<=-16'd9310;
      49141:data<=-16'd9078;
      49142:data<=-16'd8636;
      49143:data<=-16'd8969;
      49144:data<=-16'd9273;
      49145:data<=-16'd10542;
      49146:data<=-16'd10645;
      49147:data<=-16'd9764;
      49148:data<=-16'd10053;
      49149:data<=-16'd9266;
      49150:data<=-16'd10020;
      49151:data<=-16'd12223;
      49152:data<=-16'd10971;
      49153:data<=-16'd10173;
      49154:data<=-16'd10798;
      49155:data<=-16'd10031;
      49156:data<=-16'd10574;
      49157:data<=-16'd11165;
      49158:data<=-16'd10903;
      49159:data<=-16'd11097;
      49160:data<=-16'd10029;
      49161:data<=-16'd9746;
      49162:data<=-16'd10337;
      49163:data<=-16'd9966;
      49164:data<=-16'd10713;
      49165:data<=-16'd10457;
      49166:data<=-16'd9360;
      49167:data<=-16'd9659;
      49168:data<=-16'd8319;
      49169:data<=-16'd8715;
      49170:data<=-16'd11168;
      49171:data<=-16'd9541;
      49172:data<=-16'd10216;
      49173:data<=-16'd15158;
      49174:data<=-16'd15790;
      49175:data<=-16'd14653;
      49176:data<=-16'd15782;
      49177:data<=-16'd16742;
      49178:data<=-16'd14333;
      49179:data<=-16'd5588;
      49180:data<=16'd1980;
      49181:data<=16'd1040;
      49182:data<=-16'd1172;
      49183:data<=-16'd1025;
      49184:data<=-16'd1345;
      49185:data<=-16'd1204;
      49186:data<=-16'd1169;
      49187:data<=-16'd1741;
      49188:data<=-16'd2302;
      49189:data<=-16'd3368;
      49190:data<=-16'd3463;
      49191:data<=-16'd2972;
      49192:data<=-16'd2975;
      49193:data<=-16'd2355;
      49194:data<=-16'd3004;
      49195:data<=-16'd4898;
      49196:data<=-16'd5081;
      49197:data<=-16'd4673;
      49198:data<=-16'd4285;
      49199:data<=-16'd3618;
      49200:data<=-16'd4285;
      49201:data<=-16'd5509;
      49202:data<=-16'd6111;
      49203:data<=-16'd6226;
      49204:data<=-16'd5799;
      49205:data<=-16'd5547;
      49206:data<=-16'd5568;
      49207:data<=-16'd6205;
      49208:data<=-16'd7315;
      49209:data<=-16'd7221;
      49210:data<=-16'd7066;
      49211:data<=-16'd7285;
      49212:data<=-16'd6648;
      49213:data<=-16'd7280;
      49214:data<=-16'd8611;
      49215:data<=-16'd8069;
      49216:data<=-16'd7154;
      49217:data<=-16'd7174;
      49218:data<=-16'd7517;
      49219:data<=-16'd6539;
      49220:data<=-16'd7507;
      49221:data<=-16'd15920;
      49222:data<=-16'd21864;
      49223:data<=-16'd17077;
      49224:data<=-16'd13170;
      49225:data<=-16'd13964;
      49226:data<=-16'd13602;
      49227:data<=-16'd13996;
      49228:data<=-16'd13926;
      49229:data<=-16'd11934;
      49230:data<=-16'd11347;
      49231:data<=-16'd10853;
      49232:data<=-16'd9923;
      49233:data<=-16'd9583;
      49234:data<=-16'd8822;
      49235:data<=-16'd8298;
      49236:data<=-16'd7641;
      49237:data<=-16'd6875;
      49238:data<=-16'd6108;
      49239:data<=-16'd4156;
      49240:data<=-16'd3526;
      49241:data<=-16'd3541;
      49242:data<=-16'd2385;
      49243:data<=-16'd3124;
      49244:data<=-16'd2458;
      49245:data<=16'd958;
      49246:data<=16'd1298;
      49247:data<=16'd943;
      49248:data<=16'd1673;
      49249:data<=16'd1072;
      49250:data<=16'd2322;
      49251:data<=16'd4798;
      49252:data<=16'd5233;
      49253:data<=16'd4980;
      49254:data<=16'd5194;
      49255:data<=16'd5782;
      49256:data<=16'd5621;
      49257:data<=16'd6032;
      49258:data<=16'd7723;
      49259:data<=16'd7345;
      49260:data<=16'd7382;
      49261:data<=16'd7764;
      49262:data<=16'd6761;
      49263:data<=16'd14166;
      49264:data<=16'd24903;
      49265:data<=16'd24588;
      49266:data<=16'd22031;
      49267:data<=16'd22730;
      49268:data<=16'd21308;
      49269:data<=16'd21582;
      49270:data<=16'd22479;
      49271:data<=16'd21426;
      49272:data<=16'd20225;
      49273:data<=16'd16374;
      49274:data<=16'd13594;
      49275:data<=16'd14625;
      49276:data<=16'd15030;
      49277:data<=16'd15609;
      49278:data<=16'd15265;
      49279:data<=16'd13596;
      49280:data<=16'd13929;
      49281:data<=16'd13347;
      49282:data<=16'd13154;
      49283:data<=16'd14836;
      49284:data<=16'd13559;
      49285:data<=16'd12824;
      49286:data<=16'd13618;
      49287:data<=16'd11814;
      49288:data<=16'd11635;
      49289:data<=16'd12844;
      49290:data<=16'd12143;
      49291:data<=16'd11944;
      49292:data<=16'd11429;
      49293:data<=16'd10410;
      49294:data<=16'd10718;
      49295:data<=16'd11439;
      49296:data<=16'd11720;
      49297:data<=16'd10887;
      49298:data<=16'd10657;
      49299:data<=16'd10865;
      49300:data<=16'd9515;
      49301:data<=16'd10176;
      49302:data<=16'd10954;
      49303:data<=16'd9696;
      49304:data<=16'd10686;
      49305:data<=16'd5879;
      49306:data<=-16'd5283;
      49307:data<=-16'd6702;
      49308:data<=-16'd2861;
      49309:data<=-16'd3788;
      49310:data<=-16'd3345;
      49311:data<=-16'd2497;
      49312:data<=-16'd3938;
      49313:data<=-16'd3206;
      49314:data<=-16'd1624;
      49315:data<=-16'd1494;
      49316:data<=-16'd1292;
      49317:data<=-16'd558;
      49318:data<=-16'd807;
      49319:data<=-16'd1604;
      49320:data<=-16'd91;
      49321:data<=16'd1115;
      49322:data<=16'd1121;
      49323:data<=16'd4128;
      49324:data<=16'd5877;
      49325:data<=16'd4767;
      49326:data<=16'd5830;
      49327:data<=16'd6263;
      49328:data<=16'd5836;
      49329:data<=16'd6702;
      49330:data<=16'd6072;
      49331:data<=16'd5932;
      49332:data<=16'd6140;
      49333:data<=16'd4817;
      49334:data<=16'd5301;
      49335:data<=16'd5494;
      49336:data<=16'd4502;
      49337:data<=16'd4816;
      49338:data<=16'd3471;
      49339:data<=16'd1689;
      49340:data<=16'd1489;
      49341:data<=16'd1221;
      49342:data<=16'd1618;
      49343:data<=16'd1177;
      49344:data<=16'd558;
      49345:data<=-16'd538;
      49346:data<=-16'd3935;
      49347:data<=16'd804;
      49348:data<=16'd11734;
      49349:data<=16'd12891;
      49350:data<=16'd10137;
      49351:data<=16'd9865;
      49352:data<=16'd7345;
      49353:data<=16'd7072;
      49354:data<=16'd7457;
      49355:data<=16'd5383;
      49356:data<=16'd5780;
      49357:data<=16'd4902;
      49358:data<=16'd2287;
      49359:data<=16'd2505;
      49360:data<=16'd2014;
      49361:data<=16'd1236;
      49362:data<=16'd1509;
      49363:data<=16'd268;
      49364:data<=-16'd908;
      49365:data<=-16'd1512;
      49366:data<=-16'd1823;
      49367:data<=-16'd1841;
      49368:data<=-16'd2561;
      49369:data<=-16'd2588;
      49370:data<=-16'd3374;
      49371:data<=-16'd4955;
      49372:data<=-16'd5060;
      49373:data<=-16'd7407;
      49374:data<=-16'd10187;
      49375:data<=-16'd9597;
      49376:data<=-16'd10237;
      49377:data<=-16'd11414;
      49378:data<=-16'd10988;
      49379:data<=-16'd11194;
      49380:data<=-16'd10763;
      49381:data<=-16'd10296;
      49382:data<=-16'd11003;
      49383:data<=-16'd12046;
      49384:data<=-16'd12765;
      49385:data<=-16'd11400;
      49386:data<=-16'd11576;
      49387:data<=-16'd12511;
      49388:data<=-16'd9605;
      49389:data<=-16'd14128;
      49390:data<=-16'd25855;
      49391:data<=-16'd27558;
      49392:data<=-16'd24438;
      49393:data<=-16'd24859;
      49394:data<=-16'd23441;
      49395:data<=-16'd23194;
      49396:data<=-16'd24310;
      49397:data<=-16'd22566;
      49398:data<=-16'd21711;
      49399:data<=-16'd21047;
      49400:data<=-16'd18915;
      49401:data<=-16'd18688;
      49402:data<=-16'd19488;
      49403:data<=-16'd19347;
      49404:data<=-16'd18484;
      49405:data<=-16'd17370;
      49406:data<=-16'd16392;
      49407:data<=-16'd15749;
      49408:data<=-16'd16498;
      49409:data<=-16'd16964;
      49410:data<=-16'd15753;
      49411:data<=-16'd14989;
      49412:data<=-16'd13973;
      49413:data<=-16'd13438;
      49414:data<=-16'd14748;
      49415:data<=-16'd14319;
      49416:data<=-16'd12947;
      49417:data<=-16'd12377;
      49418:data<=-16'd11009;
      49419:data<=-16'd10981;
      49420:data<=-16'd11815;
      49421:data<=-16'd11969;
      49422:data<=-16'd12032;
      49423:data<=-16'd9054;
      49424:data<=-16'd5419;
      49425:data<=-16'd4589;
      49426:data<=-16'd4313;
      49427:data<=-16'd5709;
      49428:data<=-16'd5574;
      49429:data<=-16'd3557;
      49430:data<=-16'd6187;
      49431:data<=-16'd2587;
      49432:data<=16'd10116;
      49433:data<=16'd13068;
      49434:data<=16'd9617;
      49435:data<=16'd10589;
      49436:data<=16'd9862;
      49437:data<=16'd9051;
      49438:data<=16'd10674;
      49439:data<=16'd11069;
      49440:data<=16'd11846;
      49441:data<=16'd11640;
      49442:data<=16'd10390;
      49443:data<=16'd10662;
      49444:data<=16'd10229;
      49445:data<=16'd10781;
      49446:data<=16'd12239;
      49447:data<=16'd11291;
      49448:data<=16'd11004;
      49449:data<=16'd10898;
      49450:data<=16'd9655;
      49451:data<=16'd10604;
      49452:data<=16'd11535;
      49453:data<=16'd10790;
      49454:data<=16'd10516;
      49455:data<=16'd10358;
      49456:data<=16'd10120;
      49457:data<=16'd9919;
      49458:data<=16'd10525;
      49459:data<=16'd11348;
      49460:data<=16'd10457;
      49461:data<=16'd10114;
      49462:data<=16'd10072;
      49463:data<=16'd9415;
      49464:data<=16'd10848;
      49465:data<=16'd11333;
      49466:data<=16'd10063;
      49467:data<=16'd9850;
      49468:data<=16'd8921;
      49469:data<=16'd9245;
      49470:data<=16'd9818;
      49471:data<=16'd9153;
      49472:data<=16'd11832;
      49473:data<=16'd7521;
      49474:data<=-16'd6986;
      49475:data<=-16'd11776;
      49476:data<=-16'd7551;
      49477:data<=-16'd6736;
      49478:data<=-16'd6068;
      49479:data<=-16'd5470;
      49480:data<=-16'd5777;
      49481:data<=-16'd4969;
      49482:data<=-16'd4657;
      49483:data<=-16'd3034;
      49484:data<=-16'd1512;
      49485:data<=-16'd1938;
      49486:data<=-16'd969;
      49487:data<=-16'd875;
      49488:data<=-16'd1597;
      49489:data<=16'd2;
      49490:data<=16'd998;
      49491:data<=16'd1160;
      49492:data<=16'd1136;
      49493:data<=16'd428;
      49494:data<=16'd910;
      49495:data<=16'd1832;
      49496:data<=16'd2955;
      49497:data<=16'd3503;
      49498:data<=16'd2552;
      49499:data<=16'd3422;
      49500:data<=16'd4076;
      49501:data<=16'd3344;
      49502:data<=16'd4880;
      49503:data<=16'd5462;
      49504:data<=16'd4924;
      49505:data<=16'd5265;
      49506:data<=16'd4096;
      49507:data<=16'd4569;
      49508:data<=16'd6335;
      49509:data<=16'd6531;
      49510:data<=16'd6912;
      49511:data<=16'd5278;
      49512:data<=16'd4752;
      49513:data<=16'd6120;
      49514:data<=16'd3909;
      49515:data<=16'd8555;
      49516:data<=16'd19784;
      49517:data<=16'd21246;
      49518:data<=16'd18541;
      49519:data<=16'd18387;
      49520:data<=16'd17418;
      49521:data<=16'd18648;
      49522:data<=16'd18663;
      49523:data<=16'd17646;
      49524:data<=16'd20389;
      49525:data<=16'd20242;
      49526:data<=16'd18483;
      49527:data<=16'd19835;
      49528:data<=16'd19347;
      49529:data<=16'd17963;
      49530:data<=16'd17067;
      49531:data<=16'd15497;
      49532:data<=16'd15296;
      49533:data<=16'd14866;
      49534:data<=16'd14041;
      49535:data<=16'd13376;
      49536:data<=16'd11455;
      49537:data<=16'd10839;
      49538:data<=16'd10613;
      49539:data<=16'd8842;
      49540:data<=16'd7635;
      49541:data<=16'd6287;
      49542:data<=16'd5310;
      49543:data<=16'd5031;
      49544:data<=16'd3923;
      49545:data<=16'd3151;
      49546:data<=16'd1533;
      49547:data<=16'd138;
      49548:data<=16'd843;
      49549:data<=-16'd12;
      49550:data<=-16'd710;
      49551:data<=-16'd867;
      49552:data<=-16'd3265;
      49553:data<=-16'd3242;
      49554:data<=-16'd3148;
      49555:data<=-16'd4619;
      49556:data<=-16'd1968;
      49557:data<=-16'd5166;
      49558:data<=-16'd17165;
      49559:data<=-16'd21594;
      49560:data<=-16'd19076;
      49561:data<=-16'd18682;
      49562:data<=-16'd18054;
      49563:data<=-16'd17139;
      49564:data<=-16'd17916;
      49565:data<=-16'd18619;
      49566:data<=-16'd18028;
      49567:data<=-16'd17484;
      49568:data<=-16'd17537;
      49569:data<=-16'd16220;
      49570:data<=-16'd15952;
      49571:data<=-16'd17602;
      49572:data<=-16'd16871;
      49573:data<=-16'd17376;
      49574:data<=-16'd20224;
      49575:data<=-16'd19443;
      49576:data<=-16'd18762;
      49577:data<=-16'd20378;
      49578:data<=-16'd20007;
      49579:data<=-16'd19244;
      49580:data<=-16'd18189;
      49581:data<=-16'd16513;
      49582:data<=-16'd17073;
      49583:data<=-16'd17993;
      49584:data<=-16'd17854;
      49585:data<=-16'd17253;
      49586:data<=-16'd16114;
      49587:data<=-16'd15703;
      49588:data<=-16'd15151;
      49589:data<=-16'd15241;
      49590:data<=-16'd16653;
      49591:data<=-16'd15599;
      49592:data<=-16'd14339;
      49593:data<=-16'd14458;
      49594:data<=-16'd12660;
      49595:data<=-16'd12657;
      49596:data<=-16'd13840;
      49597:data<=-16'd13135;
      49598:data<=-16'd14516;
      49599:data<=-16'd10865;
      49600:data<=16'd802;
      49601:data<=16'd4760;
      49602:data<=16'd804;
      49603:data<=16'd249;
      49604:data<=16'd807;
      49605:data<=16'd710;
      49606:data<=16'd1572;
      49607:data<=16'd1140;
      49608:data<=-16'd135;
      49609:data<=-16'd848;
      49610:data<=-16'd876;
      49611:data<=-16'd550;
      49612:data<=-16'd737;
      49613:data<=-16'd672;
      49614:data<=-16'd1257;
      49615:data<=-16'd3148;
      49616:data<=-16'd3469;
      49617:data<=-16'd2573;
      49618:data<=-16'd2276;
      49619:data<=-16'd1982;
      49620:data<=-16'd2267;
      49621:data<=-16'd3535;
      49622:data<=-16'd4537;
      49623:data<=-16'd3066;
      49624:data<=16'd755;
      49625:data<=16'd2375;
      49626:data<=16'd1014;
      49627:data<=-16'd149;
      49628:data<=-16'd576;
      49629:data<=-16'd190;
      49630:data<=16'd173;
      49631:data<=-16'd20;
      49632:data<=16'd368;
      49633:data<=16'd276;
      49634:data<=16'd265;
      49635:data<=16'd961;
      49636:data<=16'd737;
      49637:data<=16'd1010;
      49638:data<=16'd746;
      49639:data<=16'd858;
      49640:data<=16'd4918;
      49641:data<=16'd2887;
      49642:data<=-16'd7755;
      49643:data<=-16'd11658;
      49644:data<=-16'd9450;
      49645:data<=-16'd8863;
      49646:data<=-16'd6724;
      49647:data<=-16'd5388;
      49648:data<=-16'd6299;
      49649:data<=-16'd5768;
      49650:data<=-16'd5486;
      49651:data<=-16'd4760;
      49652:data<=-16'd2463;
      49653:data<=-16'd1466;
      49654:data<=-16'd1061;
      49655:data<=-16'd359;
      49656:data<=-16'd182;
      49657:data<=16'd164;
      49658:data<=16'd1300;
      49659:data<=16'd2640;
      49660:data<=16'd2664;
      49661:data<=16'd2479;
      49662:data<=16'd3030;
      49663:data<=16'd2681;
      49664:data<=16'd3638;
      49665:data<=16'd5809;
      49666:data<=16'd5833;
      49667:data<=16'd6084;
      49668:data<=16'd6626;
      49669:data<=16'd5718;
      49670:data<=16'd6056;
      49671:data<=16'd7486;
      49672:data<=16'd8619;
      49673:data<=16'd7617;
      49674:data<=16'd3912;
      49675:data<=16'd2886;
      49676:data<=16'd4126;
      49677:data<=16'd4793;
      49678:data<=16'd6425;
      49679:data<=16'd5944;
      49680:data<=16'd5383;
      49681:data<=16'd6487;
      49682:data<=16'd3686;
      49683:data<=16'd7048;
      49684:data<=16'd19926;
      49685:data<=16'd23588;
      49686:data<=16'd19917;
      49687:data<=16'd20301;
      49688:data<=16'd19437;
      49689:data<=16'd18692;
      49690:data<=16'd20945;
      49691:data<=16'd20615;
      49692:data<=16'd18994;
      49693:data<=16'd18154;
      49694:data<=16'd16869;
      49695:data<=16'd17027;
      49696:data<=16'd18319;
      49697:data<=16'd18040;
      49698:data<=16'd16327;
      49699:data<=16'd15603;
      49700:data<=16'd15937;
      49701:data<=16'd15529;
      49702:data<=16'd15535;
      49703:data<=16'd15794;
      49704:data<=16'd14795;
      49705:data<=16'd14063;
      49706:data<=16'd13074;
      49707:data<=16'd11831;
      49708:data<=16'd12730;
      49709:data<=16'd13856;
      49710:data<=16'd13461;
      49711:data<=16'd12624;
      49712:data<=16'd11640;
      49713:data<=16'd11012;
      49714:data<=16'd11074;
      49715:data<=16'd12196;
      49716:data<=16'd12768;
      49717:data<=16'd11089;
      49718:data<=16'd10383;
      49719:data<=16'd10275;
      49720:data<=16'd9398;
      49721:data<=16'd10915;
      49722:data<=16'd10856;
      49723:data<=16'd9624;
      49724:data<=16'd13697;
      49725:data<=16'd12563;
      49726:data<=16'd2241;
      49727:data<=-16'd1797;
      49728:data<=16'd399;
      49729:data<=-16'd30;
      49730:data<=-16'd731;
      49731:data<=-16'd808;
      49732:data<=-16'd1080;
      49733:data<=-16'd963;
      49734:data<=-16'd1465;
      49735:data<=-16'd1380;
      49736:data<=-16'd987;
      49737:data<=-16'd1544;
      49738:data<=-16'd1394;
      49739:data<=-16'd1457;
      49740:data<=-16'd2807;
      49741:data<=-16'd3744;
      49742:data<=-16'd4061;
      49743:data<=-16'd3715;
      49744:data<=-16'd3030;
      49745:data<=-16'd3559;
      49746:data<=-16'd4966;
      49747:data<=-16'd5788;
      49748:data<=-16'd5574;
      49749:data<=-16'd5421;
      49750:data<=-16'd5809;
      49751:data<=-16'd5506;
      49752:data<=-16'd5641;
      49753:data<=-16'd7239;
      49754:data<=-16'd7956;
      49755:data<=-16'd7535;
      49756:data<=-16'd7042;
      49757:data<=-16'd6466;
      49758:data<=-16'd7119;
      49759:data<=-16'd8630;
      49760:data<=-16'd8971;
      49761:data<=-16'd8367;
      49762:data<=-16'd7887;
      49763:data<=-16'd7773;
      49764:data<=-16'd7485;
      49765:data<=-16'd8542;
      49766:data<=-16'd11403;
      49767:data<=-16'd8563;
      49768:data<=16'd1115;
      49769:data<=16'd6106;
      49770:data<=16'd4479;
      49771:data<=16'd3084;
      49772:data<=16'd2488;
      49773:data<=16'd1965;
      49774:data<=16'd414;
      49775:data<=-16'd2302;
      49776:data<=-16'd2634;
      49777:data<=-16'd2945;
      49778:data<=-16'd5456;
      49779:data<=-16'd5733;
      49780:data<=-16'd4589;
      49781:data<=-16'd4407;
      49782:data<=-16'd4167;
      49783:data<=-16'd5510;
      49784:data<=-16'd7442;
      49785:data<=-16'd7222;
      49786:data<=-16'd6693;
      49787:data<=-16'd6761;
      49788:data<=-16'd6813;
      49789:data<=-16'd7645;
      49790:data<=-16'd8927;
      49791:data<=-16'd8904;
      49792:data<=-16'd7567;
      49793:data<=-16'd7585;
      49794:data<=-16'd8514;
      49795:data<=-16'd7988;
      49796:data<=-16'd8229;
      49797:data<=-16'd9365;
      49798:data<=-16'd9031;
      49799:data<=-16'd8799;
      49800:data<=-16'd8279;
      49801:data<=-16'd7100;
      49802:data<=-16'd8193;
      49803:data<=-16'd9990;
      49804:data<=-16'd9815;
      49805:data<=-16'd8924;
      49806:data<=-16'd8557;
      49807:data<=-16'd8044;
      49808:data<=-16'd7013;
      49809:data<=-16'd10298;
      49810:data<=-16'd19173;
      49811:data<=-16'd24083;
      49812:data<=-16'd22551;
      49813:data<=-16'd21275;
      49814:data<=-16'd21200;
      49815:data<=-16'd21343;
      49816:data<=-16'd21326;
      49817:data<=-16'd20030;
      49818:data<=-16'd18851;
      49819:data<=-16'd18046;
      49820:data<=-16'd17132;
      49821:data<=-16'd16876;
      49822:data<=-16'd17048;
      49823:data<=-16'd17009;
      49824:data<=-16'd14466;
      49825:data<=-16'd10258;
      49826:data<=-16'd9256;
      49827:data<=-16'd9972;
      49828:data<=-16'd9905;
      49829:data<=-16'd10340;
      49830:data<=-16'd9784;
      49831:data<=-16'd8724;
      49832:data<=-16'd8651;
      49833:data<=-16'd7835;
      49834:data<=-16'd6949;
      49835:data<=-16'd6454;
      49836:data<=-16'd5839;
      49837:data<=-16'd5924;
      49838:data<=-16'd5547;
      49839:data<=-16'd4535;
      49840:data<=-16'd3027;
      49841:data<=-16'd1142;
      49842:data<=-16'd1704;
      49843:data<=-16'd2478;
      49844:data<=-16'd928;
      49845:data<=-16'd361;
      49846:data<=16'd312;
      49847:data<=16'd1809;
      49848:data<=16'd2117;
      49849:data<=16'd2734;
      49850:data<=16'd1656;
      49851:data<=16'd1883;
      49852:data<=16'd11188;
      49853:data<=16'd19901;
      49854:data<=16'd18961;
      49855:data<=16'd17582;
      49856:data<=16'd18398;
      49857:data<=16'd16807;
      49858:data<=16'd16402;
      49859:data<=16'd18201;
      49860:data<=16'd17981;
      49861:data<=16'd16636;
      49862:data<=16'd16284;
      49863:data<=16'd15573;
      49864:data<=16'd15135;
      49865:data<=16'd16134;
      49866:data<=16'd15934;
      49867:data<=16'd14536;
      49868:data<=16'd14509;
      49869:data<=16'd14237;
      49870:data<=16'd13007;
      49871:data<=16'd13021;
      49872:data<=16'd14079;
      49873:data<=16'd14512;
      49874:data<=16'd12557;
      49875:data<=16'd8889;
      49876:data<=16'd7374;
      49877:data<=16'd8432;
      49878:data<=16'd9415;
      49879:data<=16'd9406;
      49880:data<=16'd8849;
      49881:data<=16'd8825;
      49882:data<=16'd8878;
      49883:data<=16'd8661;
      49884:data<=16'd9815;
      49885:data<=16'd10496;
      49886:data<=16'd9128;
      49887:data<=16'd8664;
      49888:data<=16'd8683;
      49889:data<=16'd8254;
      49890:data<=16'd9201;
      49891:data<=16'd9734;
      49892:data<=16'd9774;
      49893:data<=16'd9177;
      49894:data<=16'd2053;
      49895:data<=-16'd6593;
      49896:data<=-16'd5985;
      49897:data<=-16'd2575;
      49898:data<=-16'd3559;
      49899:data<=-16'd3880;
      49900:data<=-16'd3334;
      49901:data<=-16'd3803;
      49902:data<=-16'd2413;
      49903:data<=-16'd599;
      49904:data<=-16'd579;
      49905:data<=-16'd738;
      49906:data<=-16'd734;
      49907:data<=-16'd597;
      49908:data<=16'd205;
      49909:data<=16'd1054;
      49910:data<=16'd1313;
      49911:data<=16'd1236;
      49912:data<=16'd1330;
      49913:data<=16'd1013;
      49914:data<=16'd528;
      49915:data<=16'd1676;
      49916:data<=16'd3186;
      49917:data<=16'd2977;
      49918:data<=16'd2619;
      49919:data<=16'd2651;
      49920:data<=16'd2252;
      49921:data<=16'd3102;
      49922:data<=16'd4451;
      49923:data<=16'd3654;
      49924:data<=16'd4452;
      49925:data<=16'd8254;
      49926:data<=16'd8387;
      49927:data<=16'd6837;
      49928:data<=16'd9074;
      49929:data<=16'd9549;
      49930:data<=16'd8005;
      49931:data<=16'd8545;
      49932:data<=16'd7629;
      49933:data<=16'd6904;
      49934:data<=16'd6896;
      49935:data<=16'd5442;
      49936:data<=16'd11262;
      49937:data<=16'd20381;
      49938:data<=16'd19782;
      49939:data<=16'd17106;
      49940:data<=16'd16985;
      49941:data<=16'd14220;
      49942:data<=16'd13138;
      49943:data<=16'd13176;
      49944:data<=16'd11450;
      49945:data<=16'd11203;
      49946:data<=16'd9488;
      49947:data<=16'd6300;
      49948:data<=16'd6128;
      49949:data<=16'd6325;
      49950:data<=16'd5538;
      49951:data<=16'd5030;
      49952:data<=16'd3847;
      49953:data<=16'd2232;
      49954:data<=16'd1186;
      49955:data<=16'd1365;
      49956:data<=16'd1475;
      49957:data<=16'd696;
      49958:data<=16'd582;
      49959:data<=-16'd355;
      49960:data<=-16'd2126;
      49961:data<=-16'd2272;
      49962:data<=-16'd2540;
      49963:data<=-16'd2874;
      49964:data<=-16'd2144;
      49965:data<=-16'd2945;
      49966:data<=-16'd5046;
      49967:data<=-16'd5905;
      49968:data<=-16'd5139;
      49969:data<=-16'd4578;
      49970:data<=-16'd5256;
      49971:data<=-16'd5774;
      49972:data<=-16'd6805;
      49973:data<=-16'd7483;
      49974:data<=-16'd7297;
      49975:data<=-16'd10624;
      49976:data<=-16'd12295;
      49977:data<=-16'd10097;
      49978:data<=-16'd16848;
      49979:data<=-16'd27047;
      49980:data<=-16'd26959;
      49981:data<=-16'd24686;
      49982:data<=-16'd24636;
      49983:data<=-16'd23332;
      49984:data<=-16'd24280;
      49985:data<=-16'd25118;
      49986:data<=-16'd23253;
      49987:data<=-16'd22374;
      49988:data<=-16'd21491;
      49989:data<=-16'd19967;
      49990:data<=-16'd20351;
      49991:data<=-16'd21663;
      49992:data<=-16'd21127;
      49993:data<=-16'd19306;
      49994:data<=-16'd18763;
      49995:data<=-16'd18298;
      49996:data<=-16'd17609;
      49997:data<=-16'd18627;
      49998:data<=-16'd18240;
      49999:data<=-16'd16584;
      50000:data<=-16'd16851;
      50001:data<=-16'd16193;
      50002:data<=-16'd15233;
      50003:data<=-16'd16010;
      50004:data<=-16'd15512;
      50005:data<=-16'd14694;
      50006:data<=-16'd14938;
      50007:data<=-16'd14477;
      50008:data<=-16'd13421;
      50009:data<=-16'd12888;
      50010:data<=-16'd14013;
      50011:data<=-16'd14084;
      50012:data<=-16'd11834;
      50013:data<=-16'd11775;
      50014:data<=-16'd11723;
      50015:data<=-16'd10604;
      50016:data<=-16'd12283;
      50017:data<=-16'd11517;
      50018:data<=-16'd10079;
      50019:data<=-16'd12477;
      50020:data<=-16'd6385;
      50021:data<=16'd5151;
      50022:data<=16'd5538;
      50023:data<=16'd2297;
      50024:data<=16'd4742;
      50025:data<=16'd7065;
      50026:data<=16'd8043;
      50027:data<=16'd8308;
      50028:data<=16'd6872;
      50029:data<=16'd5612;
      50030:data<=16'd4939;
      50031:data<=16'd4699;
      50032:data<=16'd4945;
      50033:data<=16'd5084;
      50034:data<=16'd5233;
      50035:data<=16'd4892;
      50036:data<=16'd4432;
      50037:data<=16'd4432;
      50038:data<=16'd4073;
      50039:data<=16'd4215;
      50040:data<=16'd5509;
      50041:data<=16'd7028;
      50042:data<=16'd7788;
      50043:data<=16'd6734;
      50044:data<=16'd5724;
      50045:data<=16'd6408;
      50046:data<=16'd7119;
      50047:data<=16'd7987;
      50048:data<=16'd8877;
      50049:data<=16'd8663;
      50050:data<=16'd8299;
      50051:data<=16'd7561;
      50052:data<=16'd7556;
      50053:data<=16'd9292;
      50054:data<=16'd9511;
      50055:data<=16'd8875;
      50056:data<=16'd9024;
      50057:data<=16'd8217;
      50058:data<=16'd8331;
      50059:data<=16'd9135;
      50060:data<=16'd9765;
      50061:data<=16'd11526;
      50062:data<=16'd6677;
      50063:data<=-16'd4531;
      50064:data<=-16'd7256;
      50065:data<=-16'd3128;
      50066:data<=-16'd2382;
      50067:data<=-16'd2417;
      50068:data<=-16'd1867;
      50069:data<=-16'd2168;
      50070:data<=-16'd1586;
      50071:data<=-16'd751;
      50072:data<=16'd446;
      50073:data<=16'd2071;
      50074:data<=16'd1453;
      50075:data<=-16'd1022;
      50076:data<=-16'd2670;
      50077:data<=-16'd2417;
      50078:data<=-16'd923;
      50079:data<=16'd332;
      50080:data<=16'd696;
      50081:data<=16'd522;
      50082:data<=16'd434;
      50083:data<=16'd318;
      50084:data<=16'd1008;
      50085:data<=16'd3210;
      50086:data<=16'd3707;
      50087:data<=16'd2867;
      50088:data<=16'd3891;
      50089:data<=16'd3902;
      50090:data<=16'd3207;
      50091:data<=16'd4323;
      50092:data<=16'd4610;
      50093:data<=16'd5291;
      50094:data<=16'd6264;
      50095:data<=16'd4971;
      50096:data<=16'd5192;
      50097:data<=16'd6475;
      50098:data<=16'd6854;
      50099:data<=16'd7799;
      50100:data<=16'd6975;
      50101:data<=16'd6808;
      50102:data<=16'd6887;
      50103:data<=16'd4079;
      50104:data<=16'd10111;
      50105:data<=16'd22307;
      50106:data<=16'd23200;
      50107:data<=16'd19749;
      50108:data<=16'd19930;
      50109:data<=16'd19197;
      50110:data<=16'd20071;
      50111:data<=16'd20155;
      50112:data<=16'd18060;
      50113:data<=16'd18607;
      50114:data<=16'd17438;
      50115:data<=16'd15603;
      50116:data<=16'd17781;
      50117:data<=16'd18177;
      50118:data<=16'd16750;
      50119:data<=16'd16615;
      50120:data<=16'd15327;
      50121:data<=16'd14462;
      50122:data<=16'd15408;
      50123:data<=16'd15807;
      50124:data<=16'd15512;
      50125:data<=16'd16659;
      50126:data<=16'd18641;
      50127:data<=16'd17801;
      50128:data<=16'd16545;
      50129:data<=16'd17811;
      50130:data<=16'd17358;
      50131:data<=16'd16004;
      50132:data<=16'd16295;
      50133:data<=16'd15546;
      50134:data<=16'd14307;
      50135:data<=16'd13244;
      50136:data<=16'd12281;
      50137:data<=16'd12061;
      50138:data<=16'd10900;
      50139:data<=16'd10372;
      50140:data<=16'd9894;
      50141:data<=16'd7591;
      50142:data<=16'd7649;
      50143:data<=16'd7019;
      50144:data<=16'd4978;
      50145:data<=16'd7450;
      50146:data<=16'd3407;
      50147:data<=-16'd9724;
      50148:data<=-16'd13823;
      50149:data<=-16'd10554;
      50150:data<=-16'd10890;
      50151:data<=-16'd11339;
      50152:data<=-16'd10777;
      50153:data<=-16'd11503;
      50154:data<=-16'd12527;
      50155:data<=-16'd12769;
      50156:data<=-16'd11891;
      50157:data<=-16'd11289;
      50158:data<=-16'd10969;
      50159:data<=-16'd11329;
      50160:data<=-16'd13082;
      50161:data<=-16'd13029;
      50162:data<=-16'd12119;
      50163:data<=-16'd12336;
      50164:data<=-16'd11265;
      50165:data<=-16'd11174;
      50166:data<=-16'd12740;
      50167:data<=-16'd12745;
      50168:data<=-16'd12616;
      50169:data<=-16'd12308;
      50170:data<=-16'd11241;
      50171:data<=-16'd11168;
      50172:data<=-16'd11377;
      50173:data<=-16'd11708;
      50174:data<=-16'd12076;
      50175:data<=-16'd13189;
      50176:data<=-16'd15437;
      50177:data<=-16'd15018;
      50178:data<=-16'd14542;
      50179:data<=-16'd16383;
      50180:data<=-16'd15235;
      50181:data<=-16'd14302;
      50182:data<=-16'd14813;
      50183:data<=-16'd12830;
      50184:data<=-16'd13958;
      50185:data<=-16'd15420;
      50186:data<=-16'd13723;
      50187:data<=-16'd15679;
      50188:data<=-16'd11505;
      50189:data<=16'd1333;
      50190:data<=16'd3909;
      50191:data<=-16'd698;
      50192:data<=-16'd778;
      50193:data<=-16'd532;
      50194:data<=-16'd462;
      50195:data<=-16'd205;
      50196:data<=-16'd1105;
      50197:data<=-16'd1051;
      50198:data<=-16'd2097;
      50199:data<=-16'd3297;
      50200:data<=-16'd2419;
      50201:data<=-16'd2569;
      50202:data<=-16'd2385;
      50203:data<=-16'd1855;
      50204:data<=-16'd3685;
      50205:data<=-16'd4326;
      50206:data<=-16'd3568;
      50207:data<=-16'd3748;
      50208:data<=-16'd3034;
      50209:data<=-16'd2693;
      50210:data<=-16'd4038;
      50211:data<=-16'd4755;
      50212:data<=-16'd4523;
      50213:data<=-16'd4231;
      50214:data<=-16'd4076;
      50215:data<=-16'd4328;
      50216:data<=-16'd5156;
      50217:data<=-16'd5700;
      50218:data<=-16'd5233;
      50219:data<=-16'd5174;
      50220:data<=-16'd5436;
      50221:data<=-16'd4966;
      50222:data<=-16'd5151;
      50223:data<=-16'd6031;
      50224:data<=-16'd6733;
      50225:data<=-16'd5554;
      50226:data<=-16'd1768;
      50227:data<=-16'd1028;
      50228:data<=-16'd2425;
      50229:data<=-16'd883;
      50230:data<=-16'd5262;
      50231:data<=-16'd16058;
      50232:data<=-16'd18950;
      50233:data<=-16'd16086;
      50234:data<=-16'd15767;
      50235:data<=-16'd15191;
      50236:data<=-16'd14120;
      50237:data<=-16'd13611;
      50238:data<=-16'd12604;
      50239:data<=-16'd12319;
      50240:data<=-16'd11621;
      50241:data<=-16'd9407;
      50242:data<=-16'd7746;
      50243:data<=-16'd7448;
      50244:data<=-16'd7642;
      50245:data<=-16'd7206;
      50246:data<=-16'd6159;
      50247:data<=-16'd4672;
      50248:data<=-16'd2913;
      50249:data<=-16'd2629;
      50250:data<=-16'd3011;
      50251:data<=-16'd2764;
      50252:data<=-16'd2966;
      50253:data<=-16'd1800;
      50254:data<=16'd517;
      50255:data<=16'd905;
      50256:data<=16'd1174;
      50257:data<=16'd1902;
      50258:data<=16'd1406;
      50259:data<=16'd1413;
      50260:data<=16'd2547;
      50261:data<=16'd3726;
      50262:data<=16'd4085;
      50263:data<=16'd3589;
      50264:data<=16'd3629;
      50265:data<=16'd3800;
      50266:data<=16'd4704;
      50267:data<=16'd6220;
      50268:data<=16'd5289;
      50269:data<=16'd5119;
      50270:data<=16'd5959;
      50271:data<=16'd3610;
      50272:data<=16'd7744;
      50273:data<=16'd19948;
      50274:data<=16'd23604;
      50275:data<=16'd19076;
      50276:data<=16'd16595;
      50277:data<=16'd14995;
      50278:data<=16'd14630;
      50279:data<=16'd15618;
      50280:data<=16'd15051;
      50281:data<=16'd14844;
      50282:data<=16'd14700;
      50283:data<=16'd13332;
      50284:data<=16'd13505;
      50285:data<=16'd15074;
      50286:data<=16'd15500;
      50287:data<=16'd14395;
      50288:data<=16'd13523;
      50289:data<=16'd13456;
      50290:data<=16'd12568;
      50291:data<=16'd12557;
      50292:data<=16'd13991;
      50293:data<=16'd13524;
      50294:data<=16'd12837;
      50295:data<=16'd13021;
      50296:data<=16'd11489;
      50297:data<=16'd10924;
      50298:data<=16'd12299;
      50299:data<=16'd12119;
      50300:data<=16'd11315;
      50301:data<=16'd11330;
      50302:data<=16'd10845;
      50303:data<=16'd10179;
      50304:data<=16'd10613;
      50305:data<=16'd11085;
      50306:data<=16'd10169;
      50307:data<=16'd9643;
      50308:data<=16'd9474;
      50309:data<=16'd8583;
      50310:data<=16'd9799;
      50311:data<=16'd10733;
      50312:data<=16'd9391;
      50313:data<=16'd10492;
      50314:data<=16'd7078;
      50315:data<=-16'd4334;
      50316:data<=-16'd8072;
      50317:data<=-16'd4070;
      50318:data<=-16'd4299;
      50319:data<=-16'd4546;
      50320:data<=-16'd3149;
      50321:data<=-16'd4088;
      50322:data<=-16'd3412;
      50323:data<=-16'd1823;
      50324:data<=-16'd2132;
      50325:data<=-16'd732;
      50326:data<=16'd1738;
      50327:data<=16'd1973;
      50328:data<=16'd2053;
      50329:data<=16'd3648;
      50330:data<=16'd4309;
      50331:data<=16'd3679;
      50332:data<=16'd3683;
      50333:data<=16'd3277;
      50334:data<=16'd2485;
      50335:data<=16'd2602;
      50336:data<=16'd1917;
      50337:data<=16'd1269;
      50338:data<=16'd1751;
      50339:data<=16'd1318;
      50340:data<=16'd825;
      50341:data<=16'd321;
      50342:data<=-16'd740;
      50343:data<=-16'd764;
      50344:data<=-16'd1400;
      50345:data<=-16'd1811;
      50346:data<=-16'd638;
      50347:data<=-16'd1707;
      50348:data<=-16'd3231;
      50349:data<=-16'd3121;
      50350:data<=-16'd3735;
      50351:data<=-16'd3504;
      50352:data<=-16'd3432;
      50353:data<=-16'd3982;
      50354:data<=-16'd4088;
      50355:data<=-16'd6980;
      50356:data<=-16'd4563;
      50357:data<=16'd6811;
      50358:data<=16'd10928;
      50359:data<=16'd7671;
      50360:data<=16'd7074;
      50361:data<=16'd5336;
      50362:data<=16'd3944;
      50363:data<=16'd4496;
      50364:data<=16'd2990;
      50365:data<=16'd2880;
      50366:data<=16'd2867;
      50367:data<=16'd658;
      50368:data<=16'd787;
      50369:data<=16'd670;
      50370:data<=-16'd696;
      50371:data<=-16'd6;
      50372:data<=-16'd602;
      50373:data<=-16'd2182;
      50374:data<=-16'd2152;
      50375:data<=-16'd3523;
      50376:data<=-16'd6065;
      50377:data<=-16'd6877;
      50378:data<=-16'd6678;
      50379:data<=-16'd7617;
      50380:data<=-16'd9085;
      50381:data<=-16'd8837;
      50382:data<=-16'd8196;
      50383:data<=-16'd8431;
      50384:data<=-16'd8334;
      50385:data<=-16'd8772;
      50386:data<=-16'd9712;
      50387:data<=-16'd9906;
      50388:data<=-16'd9964;
      50389:data<=-16'd9808;
      50390:data<=-16'd9400;
      50391:data<=-16'd9715;
      50392:data<=-16'd11248;
      50393:data<=-16'd12151;
      50394:data<=-16'd10487;
      50395:data<=-16'd9882;
      50396:data<=-16'd10504;
      50397:data<=-16'd8839;
      50398:data<=-16'd12537;
      50399:data<=-16'd22968;
      50400:data<=-16'd26706;
      50401:data<=-16'd23925;
      50402:data<=-16'd23077;
      50403:data<=-16'd22820;
      50404:data<=-16'd22674;
      50405:data<=-16'd22659;
      50406:data<=-16'd20956;
      50407:data<=-16'd20099;
      50408:data<=-16'd20010;
      50409:data<=-16'd18569;
      50410:data<=-16'd18128;
      50411:data<=-16'd19038;
      50412:data<=-16'd18645;
      50413:data<=-16'd17262;
      50414:data<=-16'd16527;
      50415:data<=-16'd16131;
      50416:data<=-16'd15987;
      50417:data<=-16'd16806;
      50418:data<=-16'd16944;
      50419:data<=-16'd15547;
      50420:data<=-16'd14624;
      50421:data<=-16'd13866;
      50422:data<=-16'd12913;
      50423:data<=-16'd13518;
      50424:data<=-16'd14119;
      50425:data<=-16'd12226;
      50426:data<=-16'd9039;
      50427:data<=-16'd7136;
      50428:data<=-16'd7298;
      50429:data<=-16'd7691;
      50430:data<=-16'd7474;
      50431:data<=-16'd7471;
      50432:data<=-16'd7013;
      50433:data<=-16'd6062;
      50434:data<=-16'd5192;
      50435:data<=-16'd4789;
      50436:data<=-16'd5729;
      50437:data<=-16'd5207;
      50438:data<=-16'd3213;
      50439:data<=-16'd4622;
      50440:data<=-16'd2661;
      50441:data<=16'd8393;
      50442:data<=16'd15380;
      50443:data<=16'd13844;
      50444:data<=16'd13705;
      50445:data<=16'd13902;
      50446:data<=16'd12005;
      50447:data<=16'd12226;
      50448:data<=16'd13159;
      50449:data<=16'd13570;
      50450:data<=16'd14249;
      50451:data<=16'd13277;
      50452:data<=16'd12176;
      50453:data<=16'd12633;
      50454:data<=16'd13180;
      50455:data<=16'd13614;
      50456:data<=16'd13552;
      50457:data<=16'd13206;
      50458:data<=16'd12935;
      50459:data<=16'd12072;
      50460:data<=16'd12405;
      50461:data<=16'd13500;
      50462:data<=16'd13007;
      50463:data<=16'd12740;
      50464:data<=16'd12601;
      50465:data<=16'd11473;
      50466:data<=16'd11720;
      50467:data<=16'd12751;
      50468:data<=16'd12739;
      50469:data<=16'd12372;
      50470:data<=16'd11770;
      50471:data<=16'd11221;
      50472:data<=16'd11095;
      50473:data<=16'd11420;
      50474:data<=16'd11996;
      50475:data<=16'd11082;
      50476:data<=16'd8545;
      50477:data<=16'd6539;
      50478:data<=16'd6143;
      50479:data<=16'd6643;
      50480:data<=16'd7268;
      50481:data<=16'd8651;
      50482:data<=16'd7089;
      50483:data<=-16'd1588;
      50484:data<=-16'd8789;
      50485:data<=-16'd7259;
      50486:data<=-16'd4165;
      50487:data<=-16'd3905;
      50488:data<=-16'd3976;
      50489:data<=-16'd3892;
      50490:data<=-16'd3676;
      50491:data<=-16'd3313;
      50492:data<=-16'd2300;
      50493:data<=-16'd861;
      50494:data<=-16'd855;
      50495:data<=-16'd1266;
      50496:data<=-16'd1246;
      50497:data<=-16'd1183;
      50498:data<=16'd238;
      50499:data<=16'd1336;
      50500:data<=16'd614;
      50501:data<=16'd288;
      50502:data<=16'd250;
      50503:data<=16'd77;
      50504:data<=16'd1102;
      50505:data<=16'd2720;
      50506:data<=16'd3468;
      50507:data<=16'd3250;
      50508:data<=16'd3133;
      50509:data<=16'd3104;
      50510:data<=16'd3380;
      50511:data<=16'd4995;
      50512:data<=16'd5536;
      50513:data<=16'd4758;
      50514:data<=16'd5342;
      50515:data<=16'd5201;
      50516:data<=16'd5063;
      50517:data<=16'd7081;
      50518:data<=16'd7383;
      50519:data<=16'd6449;
      50520:data<=16'd6501;
      50521:data<=16'd6162;
      50522:data<=16'd6572;
      50523:data<=16'd6308;
      50524:data<=16'd7040;
      50525:data<=16'd15264;
      50526:data<=16'd24040;
      50527:data<=16'd24896;
      50528:data<=16'd23417;
      50529:data<=16'd23669;
      50530:data<=16'd24040;
      50531:data<=16'd23400;
      50532:data<=16'd21796;
      50533:data<=16'd21090;
      50534:data<=16'd20603;
      50535:data<=16'd19215;
      50536:data<=16'd18363;
      50537:data<=16'd17646;
      50538:data<=16'd16983;
      50539:data<=16'd16648;
      50540:data<=16'd15760;
      50541:data<=16'd14816;
      50542:data<=16'd13194;
      50543:data<=16'd11370;
      50544:data<=16'd11210;
      50545:data<=16'd10684;
      50546:data<=16'd9755;
      50547:data<=16'd9753;
      50548:data<=16'd8310;
      50549:data<=16'd6372;
      50550:data<=16'd5697;
      50551:data<=16'd4783;
      50552:data<=16'd4488;
      50553:data<=16'd4743;
      50554:data<=16'd3592;
      50555:data<=16'd2030;
      50556:data<=16'd998;
      50557:data<=16'd20;
      50558:data<=-16'd773;
      50559:data<=-16'd893;
      50560:data<=-16'd1005;
      50561:data<=-16'd2443;
      50562:data<=-16'd3381;
      50563:data<=-16'd2981;
      50564:data<=-16'd3554;
      50565:data<=-16'd3090;
      50566:data<=-16'd3350;
      50567:data<=-16'd11439;
      50568:data<=-16'd20280;
      50569:data<=-16'd20219;
      50570:data<=-16'd18531;
      50571:data<=-16'd19513;
      50572:data<=-16'd18628;
      50573:data<=-16'd18249;
      50574:data<=-16'd19262;
      50575:data<=-16'd18463;
      50576:data<=-16'd19129;
      50577:data<=-16'd21475;
      50578:data<=-16'd21023;
      50579:data<=-16'd20562;
      50580:data<=-16'd21904;
      50581:data<=-16'd21379;
      50582:data<=-16'd20095;
      50583:data<=-16'd19675;
      50584:data<=-16'd18580;
      50585:data<=-16'd18507;
      50586:data<=-16'd19769;
      50587:data<=-16'd19549;
      50588:data<=-16'd18662;
      50589:data<=-16'd18248;
      50590:data<=-16'd17444;
      50591:data<=-16'd17004;
      50592:data<=-16'd17185;
      50593:data<=-16'd17182;
      50594:data<=-16'd16753;
      50595:data<=-16'd15758;
      50596:data<=-16'd15045;
      50597:data<=-16'd14598;
      50598:data<=-16'd14084;
      50599:data<=-16'd14784;
      50600:data<=-16'd14924;
      50601:data<=-16'd13540;
      50602:data<=-16'd13273;
      50603:data<=-16'd12320;
      50604:data<=-16'd11267;
      50605:data<=-16'd13277;
      50606:data<=-16'd13132;
      50607:data<=-16'd11518;
      50608:data<=-16'd11744;
      50609:data<=-16'd4798;
      50610:data<=16'd4892;
      50611:data<=16'd4372;
      50612:data<=16'd2193;
      50613:data<=16'd4165;
      50614:data<=16'd3882;
      50615:data<=16'd3550;
      50616:data<=16'd3739;
      50617:data<=16'd2005;
      50618:data<=16'd1240;
      50619:data<=16'd1391;
      50620:data<=16'd1968;
      50621:data<=16'd2802;
      50622:data<=16'd2196;
      50623:data<=16'd1656;
      50624:data<=16'd402;
      50625:data<=-16'd1122;
      50626:data<=16'd1071;
      50627:data<=16'd3703;
      50628:data<=16'd4179;
      50629:data<=16'd4375;
      50630:data<=16'd3250;
      50631:data<=16'd2628;
      50632:data<=16'd3304;
      50633:data<=16'd2520;
      50634:data<=16'd2140;
      50635:data<=16'd2719;
      50636:data<=16'd2500;
      50637:data<=16'd2288;
      50638:data<=16'd2203;
      50639:data<=16'd2614;
      50640:data<=16'd2887;
      50641:data<=16'd2405;
      50642:data<=16'd3363;
      50643:data<=16'd4444;
      50644:data<=16'd3956;
      50645:data<=16'd3703;
      50646:data<=16'd4064;
      50647:data<=16'd5010;
      50648:data<=16'd5473;
      50649:data<=16'd6129;
      50650:data<=16'd7785;
      50651:data<=16'd3181;
      50652:data<=-16'd5956;
      50653:data<=-16'd7671;
      50654:data<=-16'd5215;
      50655:data<=-16'd5136;
      50656:data<=-16'd4309;
      50657:data<=-16'd3254;
      50658:data<=-16'd3127;
      50659:data<=-16'd2752;
      50660:data<=-16'd2206;
      50661:data<=-16'd1133;
      50662:data<=-16'd955;
      50663:data<=-16'd1004;
      50664:data<=-16'd27;
      50665:data<=-16'd553;
      50666:data<=-16'd476;
      50667:data<=16'd1782;
      50668:data<=16'd2631;
      50669:data<=16'd2830;
      50670:data<=16'd3007;
      50671:data<=16'd1905;
      50672:data<=16'd1318;
      50673:data<=16'd2123;
      50674:data<=16'd4159;
      50675:data<=16'd5366;
      50676:data<=16'd3445;
      50677:data<=16'd917;
      50678:data<=-16'd261;
      50679:data<=16'd476;
      50680:data<=16'd2526;
      50681:data<=16'd2646;
      50682:data<=16'd2306;
      50683:data<=16'd2961;
      50684:data<=16'd2575;
      50685:data<=16'd2999;
      50686:data<=16'd4384;
      50687:data<=16'd5325;
      50688:data<=16'd5821;
      50689:data<=16'd4494;
      50690:data<=16'd4455;
      50691:data<=16'd4927;
      50692:data<=16'd3045;
      50693:data<=16'd8492;
      50694:data<=16'd18851;
      50695:data<=16'd19785;
      50696:data<=16'd17135;
      50697:data<=16'd17552;
      50698:data<=16'd16835;
      50699:data<=16'd17094;
      50700:data<=16'd17473;
      50701:data<=16'd15863;
      50702:data<=16'd15565;
      50703:data<=16'd15205;
      50704:data<=16'd14557;
      50705:data<=16'd15353;
      50706:data<=16'd15570;
      50707:data<=16'd15464;
      50708:data<=16'd14885;
      50709:data<=16'd13344;
      50710:data<=16'd13045;
      50711:data<=16'd13676;
      50712:data<=16'd14448;
      50713:data<=16'd14612;
      50714:data<=16'd13608;
      50715:data<=16'd13283;
      50716:data<=16'd12652;
      50717:data<=16'd12090;
      50718:data<=16'd13386;
      50719:data<=16'd12924;
      50720:data<=16'd11453;
      50721:data<=16'd11526;
      50722:data<=16'd10718;
      50723:data<=16'd10854;
      50724:data<=16'd11489;
      50725:data<=16'd9900;
      50726:data<=16'd10692;
      50727:data<=16'd13365;
      50728:data<=16'd13227;
      50729:data<=16'd12122;
      50730:data<=16'd12307;
      50731:data<=16'd13493;
      50732:data<=16'd12888;
      50733:data<=16'd11541;
      50734:data<=16'd12851;
      50735:data<=16'd8552;
      50736:data<=-16'd1982;
      50737:data<=-16'd5006;
      50738:data<=-16'd3169;
      50739:data<=-16'd4228;
      50740:data<=-16'd4074;
      50741:data<=-16'd3667;
      50742:data<=-16'd4951;
      50743:data<=-16'd5570;
      50744:data<=-16'd5955;
      50745:data<=-16'd6037;
      50746:data<=-16'd6138;
      50747:data<=-16'd6190;
      50748:data<=-16'd6390;
      50749:data<=-16'd8616;
      50750:data<=-16'd8925;
      50751:data<=-16'd7125;
      50752:data<=-16'd8343;
      50753:data<=-16'd8687;
      50754:data<=-16'd7632;
      50755:data<=-16'd9377;
      50756:data<=-16'd10205;
      50757:data<=-16'd9758;
      50758:data<=-16'd10108;
      50759:data<=-16'd9394;
      50760:data<=-16'd9153;
      50761:data<=-16'd10279;
      50762:data<=-16'd11292;
      50763:data<=-16'd11483;
      50764:data<=-16'd10875;
      50765:data<=-16'd10927;
      50766:data<=-16'd10430;
      50767:data<=-16'd10240;
      50768:data<=-16'd12102;
      50769:data<=-16'd11515;
      50770:data<=-16'd10569;
      50771:data<=-16'd11735;
      50772:data<=-16'd10290;
      50773:data<=-16'd10411;
      50774:data<=-16'd11941;
      50775:data<=-16'd10651;
      50776:data<=-16'd13277;
      50777:data<=-16'd12912;
      50778:data<=-16'd3374;
      50779:data<=-16'd402;
      50780:data<=-16'd3967;
      50781:data<=-16'd3897;
      50782:data<=-16'd4222;
      50783:data<=-16'd4868;
      50784:data<=-16'd3971;
      50785:data<=-16'd4055;
      50786:data<=-16'd4911;
      50787:data<=-16'd6313;
      50788:data<=-16'd6147;
      50789:data<=-16'd5262;
      50790:data<=-16'd5797;
      50791:data<=-16'd4746;
      50792:data<=-16'd5278;
      50793:data<=-16'd8078;
      50794:data<=-16'd7144;
      50795:data<=-16'd6232;
      50796:data<=-16'd6852;
      50797:data<=-16'd5744;
      50798:data<=-16'd6122;
      50799:data<=-16'd7335;
      50800:data<=-16'd7743;
      50801:data<=-16'd8144;
      50802:data<=-16'd7259;
      50803:data<=-16'd7107;
      50804:data<=-16'd7365;
      50805:data<=-16'd7215;
      50806:data<=-16'd8748;
      50807:data<=-16'd8299;
      50808:data<=-16'd6872;
      50809:data<=-16'd7720;
      50810:data<=-16'd7250;
      50811:data<=-16'd7835;
      50812:data<=-16'd9315;
      50813:data<=-16'd7949;
      50814:data<=-16'd7968;
      50815:data<=-16'd7700;
      50816:data<=-16'd6328;
      50817:data<=-16'd7506;
      50818:data<=-16'd7016;
      50819:data<=-16'd10114;
      50820:data<=-16'd19655;
      50821:data<=-16'd21781;
      50822:data<=-16'd18395;
      50823:data<=-16'd18542;
      50824:data<=-16'd18786;
      50825:data<=-16'd19238;
      50826:data<=-16'd18733;
      50827:data<=-16'd14985;
      50828:data<=-16'd12313;
      50829:data<=-16'd11376;
      50830:data<=-16'd11834;
      50831:data<=-16'd12698;
      50832:data<=-16'd11627;
      50833:data<=-16'd11652;
      50834:data<=-16'd11667;
      50835:data<=-16'd9599;
      50836:data<=-16'd9130;
      50837:data<=-16'd9094;
      50838:data<=-16'd8627;
      50839:data<=-16'd8839;
      50840:data<=-16'd7896;
      50841:data<=-16'd7376;
      50842:data<=-16'd6451;
      50843:data<=-16'd3797;
      50844:data<=-16'd3529;
      50845:data<=-16'd3905;
      50846:data<=-16'd2839;
      50847:data<=-16'd2713;
      50848:data<=-16'd1724;
      50849:data<=16'd99;
      50850:data<=16'd702;
      50851:data<=16'd829;
      50852:data<=16'd1158;
      50853:data<=16'd2026;
      50854:data<=16'd1624;
      50855:data<=16'd1518;
      50856:data<=16'd4030;
      50857:data<=16'd3849;
      50858:data<=16'd3049;
      50859:data<=16'd4460;
      50860:data<=16'd2502;
      50861:data<=16'd6143;
      50862:data<=16'd17843;
      50863:data<=16'd20280;
      50864:data<=16'd16998;
      50865:data<=16'd18093;
      50866:data<=16'd17256;
      50867:data<=16'd16551;
      50868:data<=16'd18219;
      50869:data<=16'd17155;
      50870:data<=16'd16336;
      50871:data<=16'd16707;
      50872:data<=16'd15898;
      50873:data<=16'd15606;
      50874:data<=16'd15970;
      50875:data<=16'd16827;
      50876:data<=16'd16495;
      50877:data<=16'd13515;
      50878:data<=16'd10997;
      50879:data<=16'd9853;
      50880:data<=16'd10392;
      50881:data<=16'd12152;
      50882:data<=16'd11709;
      50883:data<=16'd11130;
      50884:data<=16'd11361;
      50885:data<=16'd9891;
      50886:data<=16'd10202;
      50887:data<=16'd12073;
      50888:data<=16'd11703;
      50889:data<=16'd11250;
      50890:data<=16'd11141;
      50891:data<=16'd10220;
      50892:data<=16'd10044;
      50893:data<=16'd11080;
      50894:data<=16'd11872;
      50895:data<=16'd10766;
      50896:data<=16'd9984;
      50897:data<=16'd10390;
      50898:data<=16'd9276;
      50899:data<=16'd9771;
      50900:data<=16'd11239;
      50901:data<=16'd9959;
      50902:data<=16'd10680;
      50903:data<=16'd8172;
      50904:data<=-16'd2026;
      50905:data<=-16'd4995;
      50906:data<=-16'd802;
      50907:data<=-16'd1372;
      50908:data<=-16'd1988;
      50909:data<=-16'd1225;
      50910:data<=-16'd2453;
      50911:data<=-16'd1563;
      50912:data<=16'd394;
      50913:data<=16'd884;
      50914:data<=16'd939;
      50915:data<=16'd340;
      50916:data<=16'd173;
      50917:data<=16'd271;
      50918:data<=16'd878;
      50919:data<=16'd2611;
      50920:data<=16'd2414;
      50921:data<=16'd1768;
      50922:data<=16'd2235;
      50923:data<=16'd1158;
      50924:data<=16'd1577;
      50925:data<=16'd3413;
      50926:data<=16'd2983;
      50927:data<=16'd4413;
      50928:data<=16'd7420;
      50929:data<=16'd7145;
      50930:data<=16'd6467;
      50931:data<=16'd7553;
      50932:data<=16'd8202;
      50933:data<=16'd7981;
      50934:data<=16'd7432;
      50935:data<=16'd6802;
      50936:data<=16'd6361;
      50937:data<=16'd6167;
      50938:data<=16'd5588;
      50939:data<=16'd5018;
      50940:data<=16'd5018;
      50941:data<=16'd4306;
      50942:data<=16'd4117;
      50943:data<=16'd3603;
      50944:data<=16'd485;
      50945:data<=16'd3087;
      50946:data<=16'd12427;
      50947:data<=16'd15350;
      50948:data<=16'd13001;
      50949:data<=16'd12267;
      50950:data<=16'd10392;
      50951:data<=16'd9171;
      50952:data<=16'd9174;
      50953:data<=16'd7724;
      50954:data<=16'd7329;
      50955:data<=16'd6408;
      50956:data<=16'd4337;
      50957:data<=16'd4393;
      50958:data<=16'd3871;
      50959:data<=16'd3019;
      50960:data<=16'd3814;
      50961:data<=16'd2892;
      50962:data<=16'd1201;
      50963:data<=16'd569;
      50964:data<=-16'd253;
      50965:data<=-16'd230;
      50966:data<=16'd162;
      50967:data<=-16'd503;
      50968:data<=-16'd2130;
      50969:data<=-16'd3604;
      50970:data<=-16'd3128;
      50971:data<=-16'd3007;
      50972:data<=-16'd4002;
      50973:data<=-16'd3453;
      50974:data<=-16'd4264;
      50975:data<=-16'd6114;
      50976:data<=-16'd5515;
      50977:data<=-16'd6918;
      50978:data<=-16'd10260;
      50979:data<=-16'd10307;
      50980:data<=-16'd9815;
      50981:data<=-16'd11118;
      50982:data<=-16'd11318;
      50983:data<=-16'd10290;
      50984:data<=-16'd10460;
      50985:data<=-16'd10413;
      50986:data<=-16'd8577;
      50987:data<=-16'd12245;
      50988:data<=-16'd22266;
      50989:data<=-16'd25710;
      50990:data<=-16'd22651;
      50991:data<=-16'd22013;
      50992:data<=-16'd21516;
      50993:data<=-16'd21082;
      50994:data<=-16'd22152;
      50995:data<=-16'd21067;
      50996:data<=-16'd20119;
      50997:data<=-16'd20061;
      50998:data<=-16'd18175;
      50999:data<=-16'd17907;
      51000:data<=-16'd19180;
      51001:data<=-16'd18632;
      51002:data<=-16'd17851;
      51003:data<=-16'd17412;
      51004:data<=-16'd16472;
      51005:data<=-16'd15632;
      51006:data<=-16'd15546;
      51007:data<=-16'd16028;
      51008:data<=-16'd15547;
      51009:data<=-16'd14345;
      51010:data<=-16'd13265;
      51011:data<=-16'd12358;
      51012:data<=-16'd13164;
      51013:data<=-16'd14054;
      51014:data<=-16'd13029;
      51015:data<=-16'd12377;
      51016:data<=-16'd11671;
      51017:data<=-16'd10496;
      51018:data<=-16'd10847;
      51019:data<=-16'd11377;
      51020:data<=-16'd11182;
      51021:data<=-16'd10645;
      51022:data<=-16'd9550;
      51023:data<=-16'd8551;
      51024:data<=-16'd7958;
      51025:data<=-16'd9238;
      51026:data<=-16'd10373;
      51027:data<=-16'd7753;
      51028:data<=-16'd5400;
      51029:data<=-16'd1610;
      51030:data<=16'd7133;
      51031:data<=16'd10290;
      51032:data<=16'd7219;
      51033:data<=16'd7812;
      51034:data<=16'd8690;
      51035:data<=16'd7627;
      51036:data<=16'd7803;
      51037:data<=16'd7676;
      51038:data<=16'd7699;
      51039:data<=16'd7600;
      51040:data<=16'd7072;
      51041:data<=16'd7761;
      51042:data<=16'd7327;
      51043:data<=16'd7280;
      51044:data<=16'd9094;
      51045:data<=16'd8757;
      51046:data<=16'd8561;
      51047:data<=16'd9182;
      51048:data<=16'd7794;
      51049:data<=16'd8642;
      51050:data<=16'd10857;
      51051:data<=16'd10260;
      51052:data<=16'd9796;
      51053:data<=16'd9676;
      51054:data<=16'd8940;
      51055:data<=16'd9629;
      51056:data<=16'd10654;
      51057:data<=16'd10672;
      51058:data<=16'd10510;
      51059:data<=16'd10419;
      51060:data<=16'd9506;
      51061:data<=16'd8763;
      51062:data<=16'd10440;
      51063:data<=16'd11424;
      51064:data<=16'd10187;
      51065:data<=16'd10393;
      51066:data<=16'd10232;
      51067:data<=16'd9063;
      51068:data<=16'd9847;
      51069:data<=16'd10699;
      51070:data<=16'd11398;
      51071:data<=16'd9274;
      51072:data<=16'd735;
      51073:data<=-16'd4628;
      51074:data<=-16'd2328;
      51075:data<=-16'd326;
      51076:data<=16'd159;
      51077:data<=-16'd758;
      51078:data<=-16'd3993;
      51079:data<=-16'd5087;
      51080:data<=-16'd3748;
      51081:data<=-16'd2417;
      51082:data<=-16'd1268;
      51083:data<=-16'd1199;
      51084:data<=-16'd1254;
      51085:data<=-16'd1040;
      51086:data<=-16'd1366;
      51087:data<=-16'd543;
      51088:data<=16'd839;
      51089:data<=16'd1178;
      51090:data<=16'd1677;
      51091:data<=16'd1879;
      51092:data<=16'd934;
      51093:data<=16'd969;
      51094:data<=16'd2921;
      51095:data<=16'd4161;
      51096:data<=16'd3610;
      51097:data<=16'd3221;
      51098:data<=16'd3005;
      51099:data<=16'd3037;
      51100:data<=16'd4443;
      51101:data<=16'd5025;
      51102:data<=16'd4499;
      51103:data<=16'd4699;
      51104:data<=16'd4109;
      51105:data<=16'd3741;
      51106:data<=16'd5379;
      51107:data<=16'd6502;
      51108:data<=16'd6402;
      51109:data<=16'd5879;
      51110:data<=16'd5473;
      51111:data<=16'd5410;
      51112:data<=16'd4622;
      51113:data<=16'd7553;
      51114:data<=16'd16079;
      51115:data<=16'd20292;
      51116:data<=16'd18148;
      51117:data<=16'd17361;
      51118:data<=16'd17940;
      51119:data<=16'd18146;
      51120:data<=16'd18315;
      51121:data<=16'd17206;
      51122:data<=16'd16224;
      51123:data<=16'd15817;
      51124:data<=16'd15335;
      51125:data<=16'd15834;
      51126:data<=16'd15552;
      51127:data<=16'd15305;
      51128:data<=16'd17406;
      51129:data<=16'd17846;
      51130:data<=16'd16569;
      51131:data<=16'd17126;
      51132:data<=16'd17074;
      51133:data<=16'd16136;
      51134:data<=16'd15896;
      51135:data<=16'd14574;
      51136:data<=16'd13250;
      51137:data<=16'd12878;
      51138:data<=16'd12114;
      51139:data<=16'd11771;
      51140:data<=16'd11192;
      51141:data<=16'd9711;
      51142:data<=16'd9259;
      51143:data<=16'd8634;
      51144:data<=16'd6438;
      51145:data<=16'd5207;
      51146:data<=16'd5192;
      51147:data<=16'd4311;
      51148:data<=16'd3629;
      51149:data<=16'd3500;
      51150:data<=16'd1817;
      51151:data<=16'd337;
      51152:data<=16'd320;
      51153:data<=-16'd205;
      51154:data<=16'd575;
      51155:data<=-16'd731;
      51156:data<=-16'd10167;
      51157:data<=-16'd17438;
      51158:data<=-16'd15725;
      51159:data<=-16'd15059;
      51160:data<=-16'd16049;
      51161:data<=-16'd14337;
      51162:data<=-16'd14554;
      51163:data<=-16'd16078;
      51164:data<=-16'd15803;
      51165:data<=-16'd15672;
      51166:data<=-16'd15412;
      51167:data<=-16'd14634;
      51168:data<=-16'd14756;
      51169:data<=-16'd15520;
      51170:data<=-16'd15684;
      51171:data<=-16'd15098;
      51172:data<=-16'd15023;
      51173:data<=-16'd14877;
      51174:data<=-16'd14496;
      51175:data<=-16'd15452;
      51176:data<=-16'd15752;
      51177:data<=-16'd15655;
      51178:data<=-16'd17643;
      51179:data<=-16'd18189;
      51180:data<=-16'd16945;
      51181:data<=-16'd17822;
      51182:data<=-16'd18901;
      51183:data<=-16'd18249;
      51184:data<=-16'd17512;
      51185:data<=-16'd16948;
      51186:data<=-16'd15687;
      51187:data<=-16'd15112;
      51188:data<=-16'd16886;
      51189:data<=-16'd17444;
      51190:data<=-16'd15706;
      51191:data<=-16'd15362;
      51192:data<=-16'd14433;
      51193:data<=-16'd13529;
      51194:data<=-16'd15376;
      51195:data<=-16'd15292;
      51196:data<=-16'd14516;
      51197:data<=-16'd13253;
      51198:data<=-16'd5145;
      51199:data<=16'd1193;
      51200:data<=-16'd828;
      51201:data<=-16'd1905;
      51202:data<=-16'd1319;
      51203:data<=-16'd2056;
      51204:data<=-16'd1463;
      51205:data<=-16'd805;
      51206:data<=-16'd1157;
      51207:data<=-16'd2220;
      51208:data<=-16'd3240;
      51209:data<=-16'd2629;
      51210:data<=-16'd2399;
      51211:data<=-16'd2649;
      51212:data<=-16'd2843;
      51213:data<=-16'd4508;
      51214:data<=-16'd4652;
      51215:data<=-16'd3392;
      51216:data<=-16'd3444;
      51217:data<=-16'd2631;
      51218:data<=-16'd2561;
      51219:data<=-16'd4300;
      51220:data<=-16'd4432;
      51221:data<=-16'd4106;
      51222:data<=-16'd3920;
      51223:data<=-16'd2983;
      51224:data<=-16'd3116;
      51225:data<=-16'd4084;
      51226:data<=-16'd4977;
      51227:data<=-16'd4695;
      51228:data<=-16'd2419;
      51229:data<=-16'd387;
      51230:data<=16'd500;
      51231:data<=-16'd229;
      51232:data<=-16'd2074;
      51233:data<=-16'd1938;
      51234:data<=-16'd1263;
      51235:data<=-16'd1333;
      51236:data<=-16'd864;
      51237:data<=-16'd1345;
      51238:data<=-16'd775;
      51239:data<=-16'd505;
      51240:data<=-16'd6855;
      51241:data<=-16'd13362;
      51242:data<=-16'd13221;
      51243:data<=-16'd11764;
      51244:data<=-16'd10510;
      51245:data<=-16'd8792;
      51246:data<=-16'd8619;
      51247:data<=-16'd8392;
      51248:data<=-16'd7750;
      51249:data<=-16'd7183;
      51250:data<=-16'd5274;
      51251:data<=-16'd3862;
      51252:data<=-16'd3741;
      51253:data<=-16'd2635;
      51254:data<=-16'd1724;
      51255:data<=-16'd2490;
      51256:data<=-16'd2413;
      51257:data<=-16'd525;
      51258:data<=16'd576;
      51259:data<=16'd472;
      51260:data<=16'd514;
      51261:data<=16'd165;
      51262:data<=16'd549;
      51263:data<=16'd2549;
      51264:data<=16'd3131;
      51265:data<=16'd2443;
      51266:data<=16'd2681;
      51267:data<=16'd2601;
      51268:data<=16'd3040;
      51269:data<=16'd4893;
      51270:data<=16'd5448;
      51271:data<=16'd4855;
      51272:data<=16'd4634;
      51273:data<=16'd4592;
      51274:data<=16'd5009;
      51275:data<=16'd5577;
      51276:data<=16'd6626;
      51277:data<=16'd7238;
      51278:data<=16'd4933;
      51279:data<=16'd2375;
      51280:data<=16'd1351;
      51281:data<=16'd1996;
      51282:data<=16'd8928;
      51283:data<=16'd17050;
      51284:data<=16'd17279;
      51285:data<=16'd15455;
      51286:data<=16'd15524;
      51287:data<=16'd15009;
      51288:data<=16'd16375;
      51289:data<=16'd17224;
      51290:data<=16'd15552;
      51291:data<=16'd15277;
      51292:data<=16'd14680;
      51293:data<=16'd13717;
      51294:data<=16'd14929;
      51295:data<=16'd15054;
      51296:data<=16'd13878;
      51297:data<=16'd13505;
      51298:data<=16'd13003;
      51299:data<=16'd12446;
      51300:data<=16'd12900;
      51301:data<=16'd14853;
      51302:data<=16'd15323;
      51303:data<=16'd13267;
      51304:data<=16'd13097;
      51305:data<=16'd13241;
      51306:data<=16'd12513;
      51307:data<=16'd14225;
      51308:data<=16'd14381;
      51309:data<=16'd12504;
      51310:data<=16'd12310;
      51311:data<=16'd11256;
      51312:data<=16'd11107;
      51313:data<=16'd12677;
      51314:data<=16'd12032;
      51315:data<=16'd11294;
      51316:data<=16'd10856;
      51317:data<=16'd9870;
      51318:data<=16'd9853;
      51319:data<=16'd9523;
      51320:data<=16'd10140;
      51321:data<=16'd10621;
      51322:data<=16'd9474;
      51323:data<=16'd9433;
      51324:data<=16'd4413;
      51325:data<=-16'd3729;
      51326:data<=-16'd3621;
      51327:data<=-16'd2444;
      51328:data<=-16'd3874;
      51329:data<=-16'd1451;
      51330:data<=-16'd899;
      51331:data<=-16'd1539;
      51332:data<=16'd896;
      51333:data<=16'd902;
      51334:data<=16'd253;
      51335:data<=16'd802;
      51336:data<=16'd23;
      51337:data<=16'd247;
      51338:data<=16'd262;
      51339:data<=-16'd564;
      51340:data<=-16'd229;
      51341:data<=-16'd638;
      51342:data<=-16'd1101;
      51343:data<=-16'd1054;
      51344:data<=-16'd2017;
      51345:data<=-16'd3018;
      51346:data<=-16'd3650;
      51347:data<=-16'd3324;
      51348:data<=-16'd2946;
      51349:data<=-16'd3664;
      51350:data<=-16'd3933;
      51351:data<=-16'd5159;
      51352:data<=-16'd6287;
      51353:data<=-16'd5375;
      51354:data<=-16'd5639;
      51355:data<=-16'd5441;
      51356:data<=-16'd4975;
      51357:data<=-16'd7218;
      51358:data<=-16'd7606;
      51359:data<=-16'd7051;
      51360:data<=-16'd7133;
      51361:data<=-16'd5107;
      51362:data<=-16'd6178;
      51363:data<=-16'd8523;
      51364:data<=-16'd8132;
      51365:data<=-16'd9500;
      51366:data<=-16'd5495;
      51367:data<=16'd4253;
      51368:data<=16'd5934;
      51369:data<=16'd3072;
      51370:data<=16'd2434;
      51371:data<=16'd1638;
      51372:data<=16'd2056;
      51373:data<=16'd2378;
      51374:data<=16'd1744;
      51375:data<=16'd975;
      51376:data<=-16'd1312;
      51377:data<=-16'd1569;
      51378:data<=-16'd1063;
      51379:data<=-16'd3389;
      51380:data<=-16'd3814;
      51381:data<=-16'd3530;
      51382:data<=-16'd5274;
      51383:data<=-16'd5360;
      51384:data<=-16'd4869;
      51385:data<=-16'd4927;
      51386:data<=-16'd4573;
      51387:data<=-16'd4977;
      51388:data<=-16'd5685;
      51389:data<=-16'd6760;
      51390:data<=-16'd7174;
      51391:data<=-16'd6096;
      51392:data<=-16'd6040;
      51393:data<=-16'd5977;
      51394:data<=-16'd6059;
      51395:data<=-16'd7689;
      51396:data<=-16'd7400;
      51397:data<=-16'd6634;
      51398:data<=-16'd7062;
      51399:data<=-16'd6038;
      51400:data<=-16'd6366;
      51401:data<=-16'd7835;
      51402:data<=-16'd7720;
      51403:data<=-16'd8015;
      51404:data<=-16'd7368;
      51405:data<=-16'd6657;
      51406:data<=-16'd7228;
      51407:data<=-16'd6065;
      51408:data<=-16'd9533;
      51409:data<=-16'd18550;
      51410:data<=-16'd20879;
      51411:data<=-16'd18302;
      51412:data<=-16'd18130;
      51413:data<=-16'd17996;
      51414:data<=-16'd18186;
      51415:data<=-16'd18516;
      51416:data<=-16'd17108;
      51417:data<=-16'd15878;
      51418:data<=-16'd14948;
      51419:data<=-16'd15115;
      51420:data<=-16'd16536;
      51421:data<=-16'd15537;
      51422:data<=-16'd13530;
      51423:data<=-16'd13309;
      51424:data<=-16'd13132;
      51425:data<=-16'd12759;
      51426:data<=-16'd12760;
      51427:data<=-16'd12402;
      51428:data<=-16'd11025;
      51429:data<=-16'd9022;
      51430:data<=-16'd8062;
      51431:data<=-16'd7844;
      51432:data<=-16'd7874;
      51433:data<=-16'd8748;
      51434:data<=-16'd8810;
      51435:data<=-16'd7756;
      51436:data<=-16'd6884;
      51437:data<=-16'd6385;
      51438:data<=-16'd6551;
      51439:data<=-16'd6046;
      51440:data<=-16'd5069;
      51441:data<=-16'd5018;
      51442:data<=-16'd4487;
      51443:data<=-16'd4278;
      51444:data<=-16'd3315;
      51445:data<=-16'd399;
      51446:data<=-16'd590;
      51447:data<=-16'd934;
      51448:data<=16'd576;
      51449:data<=-16'd1657;
      51450:data<=16'd2470;
      51451:data<=16'd14657;
      51452:data<=16'd17159;
      51453:data<=16'd14455;
      51454:data<=16'd15749;
      51455:data<=16'd14334;
      51456:data<=16'd13799;
      51457:data<=16'd16131;
      51458:data<=16'd15458;
      51459:data<=16'd14865;
      51460:data<=16'd14936;
      51461:data<=16'd13894;
      51462:data<=16'd13746;
      51463:data<=16'd13691;
      51464:data<=16'd14125;
      51465:data<=16'd14653;
      51466:data<=16'd14163;
      51467:data<=16'd14201;
      51468:data<=16'd13436;
      51469:data<=16'd13071;
      51470:data<=16'd14466;
      51471:data<=16'd14170;
      51472:data<=16'd13687;
      51473:data<=16'd13494;
      51474:data<=16'd11976;
      51475:data<=16'd12612;
      51476:data<=16'd14167;
      51477:data<=16'd14017;
      51478:data<=16'd12944;
      51479:data<=16'd10505;
      51480:data<=16'd9541;
      51481:data<=16'd10348;
      51482:data<=16'd10364;
      51483:data<=16'd10903;
      51484:data<=16'd10757;
      51485:data<=16'd10386;
      51486:data<=16'd10414;
      51487:data<=16'd8793;
      51488:data<=16'd10034;
      51489:data<=16'd11934;
      51490:data<=16'd10534;
      51491:data<=16'd12107;
      51492:data<=16'd8922;
      51493:data<=-16'd2174;
      51494:data<=-16'd4018;
      51495:data<=-16'd45;
      51496:data<=-16'd1121;
      51497:data<=-16'd814;
      51498:data<=16'd106;
      51499:data<=-16'd1199;
      51500:data<=-16'd749;
      51501:data<=16'd719;
      51502:data<=16'd1777;
      51503:data<=16'd1545;
      51504:data<=16'd790;
      51505:data<=16'd1438;
      51506:data<=16'd1500;
      51507:data<=16'd2070;
      51508:data<=16'd3479;
      51509:data<=16'd2817;
      51510:data<=16'd2560;
      51511:data<=16'd2980;
      51512:data<=16'd2707;
      51513:data<=16'd3711;
      51514:data<=16'd4266;
      51515:data<=16'd4024;
      51516:data<=16'd4444;
      51517:data<=16'd3987;
      51518:data<=16'd3406;
      51519:data<=16'd3811;
      51520:data<=16'd5039;
      51521:data<=16'd5661;
      51522:data<=16'd4428;
      51523:data<=16'd4458;
      51524:data<=16'd4664;
      51525:data<=16'd3835;
      51526:data<=16'd5688;
      51527:data<=16'd6037;
      51528:data<=16'd4999;
      51529:data<=16'd7438;
      51530:data<=16'd6992;
      51531:data<=16'd5836;
      51532:data<=16'd7959;
      51533:data<=16'd6363;
      51534:data<=16'd8824;
      51535:data<=16'd18302;
      51536:data<=16'd20171;
      51537:data<=16'd17606;
      51538:data<=16'd17719;
      51539:data<=16'd15904;
      51540:data<=16'd14657;
      51541:data<=16'd14968;
      51542:data<=16'd13952;
      51543:data<=16'd13291;
      51544:data<=16'd11847;
      51545:data<=16'd9556;
      51546:data<=16'd8680;
      51547:data<=16'd7984;
      51548:data<=16'd7151;
      51549:data<=16'd6996;
      51550:data<=16'd6865;
      51551:data<=16'd5468;
      51552:data<=16'd3704;
      51553:data<=16'd3674;
      51554:data<=16'd3089;
      51555:data<=16'd2008;
      51556:data<=16'd2931;
      51557:data<=16'd1732;
      51558:data<=-16'd1313;
      51559:data<=-16'd1544;
      51560:data<=-16'd1312;
      51561:data<=-16'd1296;
      51562:data<=-16'd960;
      51563:data<=-16'd2350;
      51564:data<=-16'd3309;
      51565:data<=-16'd3243;
      51566:data<=-16'd3720;
      51567:data<=-16'd3718;
      51568:data<=-16'd3802;
      51569:data<=-16'd4308;
      51570:data<=-16'd5457;
      51571:data<=-16'd6663;
      51572:data<=-16'd5718;
      51573:data<=-16'd6075;
      51574:data<=-16'd7138;
      51575:data<=-16'd5028;
      51576:data<=-16'd8957;
      51577:data<=-16'd19089;
      51578:data<=-16'd21722;
      51579:data<=-16'd20390;
      51580:data<=-16'd21567;
      51581:data<=-16'd20324;
      51582:data<=-16'd19757;
      51583:data<=-16'd21925;
      51584:data<=-16'd21174;
      51585:data<=-16'd19506;
      51586:data<=-16'd19331;
      51587:data<=-16'd18225;
      51588:data<=-16'd17911;
      51589:data<=-16'd18970;
      51590:data<=-16'd18671;
      51591:data<=-16'd18202;
      51592:data<=-16'd18460;
      51593:data<=-16'd17202;
      51594:data<=-16'd16187;
      51595:data<=-16'd17387;
      51596:data<=-16'd17211;
      51597:data<=-16'd15790;
      51598:data<=-16'd16005;
      51599:data<=-16'd15150;
      51600:data<=-16'd13564;
      51601:data<=-16'd14489;
      51602:data<=-16'd15085;
      51603:data<=-16'd14123;
      51604:data<=-16'd13741;
      51605:data<=-16'd13250;
      51606:data<=-16'd12607;
      51607:data<=-16'd12589;
      51608:data<=-16'd12807;
      51609:data<=-16'd12605;
      51610:data<=-16'd11843;
      51611:data<=-16'd11778;
      51612:data<=-16'd11241;
      51613:data<=-16'd10173;
      51614:data<=-16'd11582;
      51615:data<=-16'd11547;
      51616:data<=-16'd9618;
      51617:data<=-16'd11147;
      51618:data<=-16'd7808;
      51619:data<=16'd2147;
      51620:data<=16'd4317;
      51621:data<=16'd1436;
      51622:data<=16'd2419;
      51623:data<=16'd2476;
      51624:data<=16'd1915;
      51625:data<=16'd2860;
      51626:data<=16'd1874;
      51627:data<=16'd673;
      51628:data<=16'd1212;
      51629:data<=16'd2387;
      51630:data<=16'd3571;
      51631:data<=16'd3418;
      51632:data<=16'd2679;
      51633:data<=16'd2341;
      51634:data<=16'd1812;
      51635:data<=16'd1701;
      51636:data<=16'd1807;
      51637:data<=16'd1706;
      51638:data<=16'd1404;
      51639:data<=16'd1115;
      51640:data<=16'd1917;
      51641:data<=16'd2288;
      51642:data<=16'd1642;
      51643:data<=16'd1952;
      51644:data<=16'd2428;
      51645:data<=16'd3357;
      51646:data<=16'd4632;
      51647:data<=16'd4296;
      51648:data<=16'd4446;
      51649:data<=16'd4634;
      51650:data<=16'd3721;
      51651:data<=16'd5057;
      51652:data<=16'd6398;
      51653:data<=16'd6044;
      51654:data<=16'd6566;
      51655:data<=16'd5965;
      51656:data<=16'd5133;
      51657:data<=16'd5661;
      51658:data<=16'd5991;
      51659:data<=16'd7520;
      51660:data<=16'd4999;
      51661:data<=-16'd3826;
      51662:data<=-16'd7426;
      51663:data<=-16'd5175;
      51664:data<=-16'd4452;
      51665:data<=-16'd3551;
      51666:data<=-16'd2822;
      51667:data<=-16'd3304;
      51668:data<=-16'd2990;
      51669:data<=-16'd2675;
      51670:data<=-16'd1525;
      51671:data<=16'd61;
      51672:data<=-16'd199;
      51673:data<=-16'd241;
      51674:data<=16'd293;
      51675:data<=16'd77;
      51676:data<=16'd755;
      51677:data<=16'd2309;
      51678:data<=16'd2598;
      51679:data<=16'd1219;
      51680:data<=16'd229;
      51681:data<=16'd273;
      51682:data<=16'd364;
      51683:data<=16'd1677;
      51684:data<=16'd3078;
      51685:data<=16'd2745;
      51686:data<=16'd2852;
      51687:data<=16'd2837;
      51688:data<=16'd2743;
      51689:data<=16'd4717;
      51690:data<=16'd5536;
      51691:data<=16'd4731;
      51692:data<=16'd4810;
      51693:data<=16'd4376;
      51694:data<=16'd4435;
      51695:data<=16'd5495;
      51696:data<=16'd5923;
      51697:data<=16'd6234;
      51698:data<=16'd5773;
      51699:data<=16'd5961;
      51700:data<=16'd6567;
      51701:data<=16'd5049;
      51702:data<=16'd8526;
      51703:data<=16'd17277;
      51704:data<=16'd19835;
      51705:data<=16'd18211;
      51706:data<=16'd18090;
      51707:data<=16'd17394;
      51708:data<=16'd17637;
      51709:data<=16'd18117;
      51710:data<=16'd16998;
      51711:data<=16'd16592;
      51712:data<=16'd15854;
      51713:data<=16'd15060;
      51714:data<=16'd15879;
      51715:data<=16'd15803;
      51716:data<=16'd14828;
      51717:data<=16'd14236;
      51718:data<=16'd13435;
      51719:data<=16'd12844;
      51720:data<=16'd12892;
      51721:data<=16'd13443;
      51722:data<=16'd12974;
      51723:data<=16'd11765;
      51724:data<=16'd11846;
      51725:data<=16'd10969;
      51726:data<=16'd9828;
      51727:data<=16'd10956;
      51728:data<=16'd10827;
      51729:data<=16'd10560;
      51730:data<=16'd12044;
      51731:data<=16'd11204;
      51732:data<=16'd10454;
      51733:data<=16'd11866;
      51734:data<=16'd11756;
      51735:data<=16'd10796;
      51736:data<=16'd9674;
      51737:data<=16'd8724;
      51738:data<=16'd8786;
      51739:data<=16'd7812;
      51740:data<=16'd7148;
      51741:data<=16'd6463;
      51742:data<=16'd4573;
      51743:data<=16'd5805;
      51744:data<=16'd4225;
      51745:data<=-16'd5568;
      51746:data<=-16'd11464;
      51747:data<=-16'd10527;
      51748:data<=-16'd10742;
      51749:data<=-16'd10540;
      51750:data<=-16'd9445;
      51751:data<=-16'd10516;
      51752:data<=-16'd11753;
      51753:data<=-16'd11640;
      51754:data<=-16'd11189;
      51755:data<=-16'd11141;
      51756:data<=-16'd10988;
      51757:data<=-16'd10742;
      51758:data<=-16'd11550;
      51759:data<=-16'd12172;
      51760:data<=-16'd12157;
      51761:data<=-16'd12304;
      51762:data<=-16'd11330;
      51763:data<=-16'd10754;
      51764:data<=-16'd11937;
      51765:data<=-16'd12396;
      51766:data<=-16'd11984;
      51767:data<=-16'd11312;
      51768:data<=-16'd10345;
      51769:data<=-16'd10213;
      51770:data<=-16'd10762;
      51771:data<=-16'd11570;
      51772:data<=-16'd11726;
      51773:data<=-16'd10988;
      51774:data<=-16'd10877;
      51775:data<=-16'd10510;
      51776:data<=-16'd10646;
      51777:data<=-16'd12022;
      51778:data<=-16'd11291;
      51779:data<=-16'd11107;
      51780:data<=-16'd12944;
      51781:data<=-16'd12093;
      51782:data<=-16'd11779;
      51783:data<=-16'd13074;
      51784:data<=-16'd12231;
      51785:data<=-16'd12794;
      51786:data<=-16'd10931;
      51787:data<=-16'd2041;
      51788:data<=16'd2770;
      51789:data<=16'd379;
      51790:data<=-16'd799;
      51791:data<=-16'd600;
      51792:data<=-16'd1078;
      51793:data<=-16'd1049;
      51794:data<=-16'd937;
      51795:data<=-16'd1726;
      51796:data<=-16'd2761;
      51797:data<=-16'd2761;
      51798:data<=-16'd2905;
      51799:data<=-16'd3195;
      51800:data<=-16'd2253;
      51801:data<=-16'd2801;
      51802:data<=-16'd4358;
      51803:data<=-16'd4074;
      51804:data<=-16'd4402;
      51805:data<=-16'd4698;
      51806:data<=-16'd3507;
      51807:data<=-16'd4030;
      51808:data<=-16'd5274;
      51809:data<=-16'd5658;
      51810:data<=-16'd5982;
      51811:data<=-16'd5027;
      51812:data<=-16'd4452;
      51813:data<=-16'd5357;
      51814:data<=-16'd5554;
      51815:data<=-16'd5868;
      51816:data<=-16'd6391;
      51817:data<=-16'd6049;
      51818:data<=-16'd5585;
      51819:data<=-16'd5037;
      51820:data<=-16'd5582;
      51821:data<=-16'd6778;
      51822:data<=-16'd6522;
      51823:data<=-16'd6448;
      51824:data<=-16'd6216;
      51825:data<=-16'd5379;
      51826:data<=-16'd6278;
      51827:data<=-16'd6570;
      51828:data<=-16'd7861;
      51829:data<=-16'd14092;
      51830:data<=-16'd17393;
      51831:data<=-16'd15095;
      51832:data<=-16'd15062;
      51833:data<=-16'd16079;
      51834:data<=-16'd15153;
      51835:data<=-16'd14774;
      51836:data<=-16'd14070;
      51837:data<=-16'd13118;
      51838:data<=-16'd13165;
      51839:data<=-16'd12207;
      51840:data<=-16'd11007;
      51841:data<=-16'd10985;
      51842:data<=-16'd10103;
      51843:data<=-16'd8922;
      51844:data<=-16'd9119;
      51845:data<=-16'd8293;
      51846:data<=-16'd5976;
      51847:data<=-16'd5256;
      51848:data<=-16'd4966;
      51849:data<=-16'd3483;
      51850:data<=-16'd3412;
      51851:data<=-16'd3248;
      51852:data<=-16'd984;
      51853:data<=-16'd314;
      51854:data<=-16'd561;
      51855:data<=16'd757;
      51856:data<=16'd781;
      51857:data<=16'd337;
      51858:data<=16'd2105;
      51859:data<=16'd3418;
      51860:data<=16'd2936;
      51861:data<=16'd2845;
      51862:data<=16'd3510;
      51863:data<=16'd3348;
      51864:data<=16'd3459;
      51865:data<=16'd5268;
      51866:data<=16'd5691;
      51867:data<=16'd5307;
      51868:data<=16'd6399;
      51869:data<=16'd5121;
      51870:data<=16'd6052;
      51871:data<=16'd14998;
      51872:data<=16'd20850;
      51873:data<=16'd19497;
      51874:data<=16'd19112;
      51875:data<=16'd18679;
      51876:data<=16'd17703;
      51877:data<=16'd19059;
      51878:data<=16'd19358;
      51879:data<=16'd17940;
      51880:data<=16'd16437;
      51881:data<=16'd14610;
      51882:data<=16'd14220;
      51883:data<=16'd15148;
      51884:data<=16'd15388;
      51885:data<=16'd14719;
      51886:data<=16'd14187;
      51887:data<=16'd14264;
      51888:data<=16'd13502;
      51889:data<=16'd13364;
      51890:data<=16'd14838;
      51891:data<=16'd14313;
      51892:data<=16'd13432;
      51893:data<=16'd13635;
      51894:data<=16'd11934;
      51895:data<=16'd11896;
      51896:data<=16'd13957;
      51897:data<=16'd13362;
      51898:data<=16'd12612;
      51899:data<=16'd12326;
      51900:data<=16'd10803;
      51901:data<=16'd10941;
      51902:data<=16'd12270;
      51903:data<=16'd12668;
      51904:data<=16'd12061;
      51905:data<=16'd11106;
      51906:data<=16'd11159;
      51907:data<=16'd10753;
      51908:data<=16'd10595;
      51909:data<=16'd11796;
      51910:data<=16'd10818;
      51911:data<=16'd10507;
      51912:data<=16'd10619;
      51913:data<=16'd3432;
      51914:data<=-16'd3119;
      51915:data<=-16'd1321;
      51916:data<=-16'd296;
      51917:data<=-16'd1397;
      51918:data<=-16'd881;
      51919:data<=-16'd1524;
      51920:data<=-16'd1284;
      51921:data<=16'd878;
      51922:data<=16'd1092;
      51923:data<=16'd446;
      51924:data<=16'd522;
      51925:data<=16'd200;
      51926:data<=16'd579;
      51927:data<=16'd1965;
      51928:data<=16'd2076;
      51929:data<=16'd1707;
      51930:data<=16'd3060;
      51931:data<=16'd3624;
      51932:data<=16'd2807;
      51933:data<=16'd4131;
      51934:data<=16'd5738;
      51935:data<=16'd5321;
      51936:data<=16'd5083;
      51937:data<=16'd4666;
      51938:data<=16'd4068;
      51939:data<=16'd4513;
      51940:data<=16'd4272;
      51941:data<=16'd3618;
      51942:data<=16'd3542;
      51943:data<=16'd3137;
      51944:data<=16'd3075;
      51945:data<=16'd2726;
      51946:data<=16'd1086;
      51947:data<=-16'd282;
      51948:data<=-16'd764;
      51949:data<=-16'd456;
      51950:data<=-16'd300;
      51951:data<=-16'd1007;
      51952:data<=-16'd1193;
      51953:data<=-16'd2435;
      51954:data<=-16'd3318;
      51955:data<=16'd2519;
      51956:data<=16'd9935;
      51957:data<=16'd10396;
      51958:data<=16'd8156;
      51959:data<=16'd7130;
      51960:data<=16'd6008;
      51961:data<=16'd5466;
      51962:data<=16'd5301;
      51963:data<=16'd5165;
      51964:data<=16'd4493;
      51965:data<=16'd2475;
      51966:data<=16'd1726;
      51967:data<=16'd2111;
      51968:data<=16'd1465;
      51969:data<=16'd1515;
      51970:data<=16'd1339;
      51971:data<=-16'd506;
      51972:data<=-16'd1339;
      51973:data<=-16'd1113;
      51974:data<=-16'd1328;
      51975:data<=-16'd1760;
      51976:data<=-16'd2396;
      51977:data<=-16'd3301;
      51978:data<=-16'd4370;
      51979:data<=-16'd4611;
      51980:data<=-16'd4943;
      51981:data<=-16'd6508;
      51982:data<=-16'd6294;
      51983:data<=-16'd6049;
      51984:data<=-16'd8463;
      51985:data<=-16'd8621;
      51986:data<=-16'd7298;
      51987:data<=-16'd7454;
      51988:data<=-16'd6539;
      51989:data<=-16'd7050;
      51990:data<=-16'd9103;
      51991:data<=-16'd9050;
      51992:data<=-16'd8865;
      51993:data<=-16'd8461;
      51994:data<=-16'd8573;
      51995:data<=-16'd9774;
      51996:data<=-16'd8998;
      51997:data<=-16'd12913;
      51998:data<=-16'd21511;
      51999:data<=-16'd22419;
      52000:data<=-16'd19654;
      52001:data<=-16'd19919;
      52002:data<=-16'd19371;
      52003:data<=-16'd19658;
      52004:data<=-16'd20080;
      52005:data<=-16'd18457;
      52006:data<=-16'd17744;
      52007:data<=-16'd16806;
      52008:data<=-16'd16634;
      52009:data<=-16'd18187;
      52010:data<=-16'd17340;
      52011:data<=-16'd16095;
      52012:data<=-16'd15908;
      52013:data<=-16'd14707;
      52014:data<=-16'd14774;
      52015:data<=-16'd15675;
      52016:data<=-16'd15179;
      52017:data<=-16'd14087;
      52018:data<=-16'd13073;
      52019:data<=-16'd12546;
      52020:data<=-16'd12087;
      52021:data<=-16'd12508;
      52022:data<=-16'd13456;
      52023:data<=-16'd12448;
      52024:data<=-16'd11847;
      52025:data<=-16'd11489;
      52026:data<=-16'd9577;
      52027:data<=-16'd10439;
      52028:data<=-16'd12157;
      52029:data<=-16'd11163;
      52030:data<=-16'd9890;
      52031:data<=-16'd7674;
      52032:data<=-16'd6643;
      52033:data<=-16'd7876;
      52034:data<=-16'd7683;
      52035:data<=-16'd8044;
      52036:data<=-16'd7212;
      52037:data<=-16'd5457;
      52038:data<=-16'd7973;
      52039:data<=-16'd4387;
      52040:data<=16'd6263;
      52041:data<=16'd8258;
      52042:data<=16'd6249;
      52043:data<=16'd7615;
      52044:data<=16'd6789;
      52045:data<=16'd6443;
      52046:data<=16'd8281;
      52047:data<=16'd8422;
      52048:data<=16'd7900;
      52049:data<=16'd7932;
      52050:data<=16'd8284;
      52051:data<=16'd7943;
      52052:data<=16'd7677;
      52053:data<=16'd9039;
      52054:data<=16'd9198;
      52055:data<=16'd8833;
      52056:data<=16'd9294;
      52057:data<=16'd8035;
      52058:data<=16'd8122;
      52059:data<=16'd9790;
      52060:data<=16'd9179;
      52061:data<=16'd8895;
      52062:data<=16'd8831;
      52063:data<=16'd7814;
      52064:data<=16'd8542;
      52065:data<=16'd9468;
      52066:data<=16'd9477;
      52067:data<=16'd9268;
      52068:data<=16'd8504;
      52069:data<=16'd8478;
      52070:data<=16'd8642;
      52071:data<=16'd9145;
      52072:data<=16'd10105;
      52073:data<=16'd9279;
      52074:data<=16'd9279;
      52075:data<=16'd9641;
      52076:data<=16'd7899;
      52077:data<=16'd8849;
      52078:data<=16'd10146;
      52079:data<=16'd9162;
      52080:data<=16'd10020;
      52081:data<=16'd5033;
      52082:data<=-16'd5638;
      52083:data<=-16'd6939;
      52084:data<=-16'd2969;
      52085:data<=-16'd3541;
      52086:data<=-16'd3879;
      52087:data<=-16'd3078;
      52088:data<=-16'd3342;
      52089:data<=-16'd2417;
      52090:data<=-16'd644;
      52091:data<=16'd2;
      52092:data<=-16'd544;
      52093:data<=-16'd600;
      52094:data<=-16'd133;
      52095:data<=-16'd625;
      52096:data<=16'd70;
      52097:data<=16'd2014;
      52098:data<=16'd1968;
      52099:data<=16'd1242;
      52100:data<=16'd961;
      52101:data<=16'd743;
      52102:data<=16'd2455;
      52103:data<=16'd4358;
      52104:data<=16'd4002;
      52105:data<=16'd3466;
      52106:data<=16'd3385;
      52107:data<=16'd3171;
      52108:data<=16'd3867;
      52109:data<=16'd4992;
      52110:data<=16'd5154;
      52111:data<=16'd4643;
      52112:data<=16'd4303;
      52113:data<=16'd3949;
      52114:data<=16'd3991;
      52115:data<=16'd5154;
      52116:data<=16'd5585;
      52117:data<=16'd5060;
      52118:data<=16'd5262;
      52119:data<=16'd4678;
      52120:data<=16'd4457;
      52121:data<=16'd5767;
      52122:data<=16'd5238;
      52123:data<=16'd8029;
      52124:data<=16'd16780;
      52125:data<=16'd19135;
      52126:data<=16'd15606;
      52127:data<=16'd17024;
      52128:data<=16'd18287;
      52129:data<=16'd16007;
      52130:data<=16'd16290;
      52131:data<=16'd17232;
      52132:data<=16'd16224;
      52133:data<=16'd16073;
      52134:data<=16'd16806;
      52135:data<=16'd16660;
      52136:data<=16'd15479;
      52137:data<=16'd14451;
      52138:data<=16'd13946;
      52139:data<=16'd13332;
      52140:data<=16'd12789;
      52141:data<=16'd12101;
      52142:data<=16'd11474;
      52143:data<=16'd10740;
      52144:data<=16'd9289;
      52145:data<=16'd9054;
      52146:data<=16'd8587;
      52147:data<=16'd5800;
      52148:data<=16'd4819;
      52149:data<=16'd5145;
      52150:data<=16'd4241;
      52151:data<=16'd4655;
      52152:data<=16'd4082;
      52153:data<=16'd1550;
      52154:data<=16'd1436;
      52155:data<=16'd1962;
      52156:data<=16'd1081;
      52157:data<=16'd635;
      52158:data<=16'd52;
      52159:data<=-16'd1366;
      52160:data<=-16'd2372;
      52161:data<=-16'd2055;
      52162:data<=-16'd2569;
      52163:data<=-16'd3284;
      52164:data<=-16'd1254;
      52165:data<=-16'd4886;
      52166:data<=-16'd15717;
      52167:data<=-16'd18556;
      52168:data<=-16'd15441;
      52169:data<=-16'd16230;
      52170:data<=-16'd15594;
      52171:data<=-16'd14912;
      52172:data<=-16'd17208;
      52173:data<=-16'd16528;
      52174:data<=-16'd15082;
      52175:data<=-16'd15259;
      52176:data<=-16'd14580;
      52177:data<=-16'd15189;
      52178:data<=-16'd16110;
      52179:data<=-16'd15183;
      52180:data<=-16'd15038;
      52181:data<=-16'd16173;
      52182:data<=-16'd16542;
      52183:data<=-16'd15767;
      52184:data<=-16'd16057;
      52185:data<=-16'd16892;
      52186:data<=-16'd15534;
      52187:data<=-16'd14700;
      52188:data<=-16'd14739;
      52189:data<=-16'd13145;
      52190:data<=-16'd13702;
      52191:data<=-16'd15612;
      52192:data<=-16'd14654;
      52193:data<=-16'd13870;
      52194:data<=-16'd13870;
      52195:data<=-16'd13051;
      52196:data<=-16'd13715;
      52197:data<=-16'd15026;
      52198:data<=-16'd14378;
      52199:data<=-16'd13039;
      52200:data<=-16'd12624;
      52201:data<=-16'd11911;
      52202:data<=-16'd11483;
      52203:data<=-16'd13024;
      52204:data<=-16'd12533;
      52205:data<=-16'd11025;
      52206:data<=-16'd13177;
      52207:data<=-16'd9718;
      52208:data<=16'd469;
      52209:data<=16'd2461;
      52210:data<=-16'd638;
      52211:data<=16'd553;
      52212:data<=16'd913;
      52213:data<=16'd191;
      52214:data<=16'd990;
      52215:data<=16'd114;
      52216:data<=-16'd1394;
      52217:data<=-16'd1528;
      52218:data<=-16'd1169;
      52219:data<=-16'd637;
      52220:data<=-16'd605;
      52221:data<=-16'd1518;
      52222:data<=-16'd2743;
      52223:data<=-16'd2795;
      52224:data<=-16'd2044;
      52225:data<=-16'd2238;
      52226:data<=-16'd1939;
      52227:data<=-16'd1575;
      52228:data<=-16'd3095;
      52229:data<=-16'd3826;
      52230:data<=-16'd3046;
      52231:data<=-16'd2000;
      52232:data<=-16'd402;
      52233:data<=-16'd370;
      52234:data<=-16'd1730;
      52235:data<=-16'd2093;
      52236:data<=-16'd2038;
      52237:data<=-16'd1641;
      52238:data<=-16'd1286;
      52239:data<=-16'd1498;
      52240:data<=-16'd1284;
      52241:data<=-16'd1242;
      52242:data<=-16'd1031;
      52243:data<=-16'd540;
      52244:data<=-16'd839;
      52245:data<=-16'd453;
      52246:data<=-16'd9;
      52247:data<=16'd980;
      52248:data<=16'd3847;
      52249:data<=16'd772;
      52250:data<=-16'd8420;
      52251:data<=-16'd11458;
      52252:data<=-16'd8830;
      52253:data<=-16'd7659;
      52254:data<=-16'd7100;
      52255:data<=-16'd6610;
      52256:data<=-16'd6302;
      52257:data<=-16'd5946;
      52258:data<=-16'd5871;
      52259:data<=-16'd4246;
      52260:data<=-16'd2370;
      52261:data<=-16'd2356;
      52262:data<=-16'd2008;
      52263:data<=-16'd1451;
      52264:data<=-16'd1645;
      52265:data<=-16'd710;
      52266:data<=16'd917;
      52267:data<=16'd1488;
      52268:data<=16'd1387;
      52269:data<=16'd1416;
      52270:data<=16'd1553;
      52271:data<=16'd2243;
      52272:data<=16'd3944;
      52273:data<=16'd4642;
      52274:data<=16'd3811;
      52275:data<=16'd4064;
      52276:data<=16'd4487;
      52277:data<=16'd3932;
      52278:data<=16'd4796;
      52279:data<=16'd6031;
      52280:data<=16'd5300;
      52281:data<=16'd3999;
      52282:data<=16'd3304;
      52283:data<=16'd3172;
      52284:data<=16'd3912;
      52285:data<=16'd5348;
      52286:data<=16'd5683;
      52287:data<=16'd4640;
      52288:data<=16'd5222;
      52289:data<=16'd5665;
      52290:data<=16'd4309;
      52291:data<=16'd8921;
      52292:data<=16'd18240;
      52293:data<=16'd20630;
      52294:data<=16'd18427;
      52295:data<=16'd18460;
      52296:data<=16'd18551;
      52297:data<=16'd18621;
      52298:data<=16'd18915;
      52299:data<=16'd17922;
      52300:data<=16'd17364;
      52301:data<=16'd16697;
      52302:data<=16'd15479;
      52303:data<=16'd16163;
      52304:data<=16'd16818;
      52305:data<=16'd15473;
      52306:data<=16'd14657;
      52307:data<=16'd14728;
      52308:data<=16'd14202;
      52309:data<=16'd14205;
      52310:data<=16'd15095;
      52311:data<=16'd14730;
      52312:data<=16'd13706;
      52313:data<=16'd13571;
      52314:data<=16'd12809;
      52315:data<=16'd12377;
      52316:data<=16'd13335;
      52317:data<=16'd13035;
      52318:data<=16'd12519;
      52319:data<=16'd12627;
      52320:data<=16'd11348;
      52321:data<=16'd11192;
      52322:data<=16'd12560;
      52323:data<=16'd12542;
      52324:data<=16'd11950;
      52325:data<=16'd10980;
      52326:data<=16'd9941;
      52327:data<=16'd9984;
      52328:data<=16'd10454;
      52329:data<=16'd11320;
      52330:data<=16'd10540;
      52331:data<=16'd9724;
      52332:data<=16'd12419;
      52333:data<=16'd9659;
      52334:data<=16'd315;
      52335:data<=-16'd2124;
      52336:data<=-16'd277;
      52337:data<=-16'd1478;
      52338:data<=-16'd1366;
      52339:data<=-16'd919;
      52340:data<=-16'd1812;
      52341:data<=-16'd1676;
      52342:data<=-16'd1803;
      52343:data<=-16'd1765;
      52344:data<=-16'd1503;
      52345:data<=-16'd1958;
      52346:data<=-16'd1657;
      52347:data<=-16'd2311;
      52348:data<=-16'd3585;
      52349:data<=-16'd3119;
      52350:data<=-16'd3444;
      52351:data<=-16'd3845;
      52352:data<=-16'd2946;
      52353:data<=-16'd3876;
      52354:data<=-16'd5166;
      52355:data<=-16'd4494;
      52356:data<=-16'd3974;
      52357:data<=-16'd3962;
      52358:data<=-16'd3761;
      52359:data<=-16'd4394;
      52360:data<=-16'd6031;
      52361:data<=-16'd6754;
      52362:data<=-16'd6176;
      52363:data<=-16'd6056;
      52364:data<=-16'd6129;
      52365:data<=-16'd6481;
      52366:data<=-16'd7532;
      52367:data<=-16'd7295;
      52368:data<=-16'd6769;
      52369:data<=-16'd6937;
      52370:data<=-16'd6446;
      52371:data<=-16'd7136;
      52372:data<=-16'd7950;
      52373:data<=-16'd7639;
      52374:data<=-16'd8812;
      52375:data<=-16'd5950;
      52376:data<=16'd3036;
      52377:data<=16'd6986;
      52378:data<=16'd4226;
      52379:data<=16'd2867;
      52380:data<=16'd3341;
      52381:data<=16'd2534;
      52382:data<=16'd1175;
      52383:data<=16'd1131;
      52384:data<=16'd625;
      52385:data<=-16'd1441;
      52386:data<=-16'd1642;
      52387:data<=-16'd904;
      52388:data<=-16'd1656;
      52389:data<=-16'd1721;
      52390:data<=-16'd2158;
      52391:data<=-16'd3770;
      52392:data<=-16'd4076;
      52393:data<=-16'd4173;
      52394:data<=-16'd4385;
      52395:data<=-16'd3779;
      52396:data<=-16'd3918;
      52397:data<=-16'd5001;
      52398:data<=-16'd6181;
      52399:data<=-16'd6278;
      52400:data<=-16'd5285;
      52401:data<=-16'd5089;
      52402:data<=-16'd4760;
      52403:data<=-16'd4769;
      52404:data<=-16'd6504;
      52405:data<=-16'd6760;
      52406:data<=-16'd6067;
      52407:data<=-16'd6352;
      52408:data<=-16'd5765;
      52409:data<=-16'd6050;
      52410:data<=-16'd7180;
      52411:data<=-16'd6945;
      52412:data<=-16'd7138;
      52413:data<=-16'd6787;
      52414:data<=-16'd6187;
      52415:data<=-16'd7018;
      52416:data<=-16'd6416;
      52417:data<=-16'd8947;
      52418:data<=-16'd17156;
      52419:data<=-16'd20392;
      52420:data<=-16'd18134;
      52421:data<=-16'd18033;
      52422:data<=-16'd18541;
      52423:data<=-16'd18442;
      52424:data<=-16'd18269;
      52425:data<=-16'd17170;
      52426:data<=-16'd16715;
      52427:data<=-16'd16061;
      52428:data<=-16'd14879;
      52429:data<=-16'd15432;
      52430:data<=-16'd15481;
      52431:data<=-16'd13579;
      52432:data<=-16'd11996;
      52433:data<=-16'd11095;
      52434:data<=-16'd10988;
      52435:data<=-16'd11505;
      52436:data<=-16'd11430;
      52437:data<=-16'd11015;
      52438:data<=-16'd10420;
      52439:data<=-16'd9544;
      52440:data<=-16'd9034;
      52441:data<=-16'd8648;
      52442:data<=-16'd7965;
      52443:data<=-16'd7394;
      52444:data<=-16'd7171;
      52445:data<=-16'd7003;
      52446:data<=-16'd6305;
      52447:data<=-16'd4872;
      52448:data<=-16'd3718;
      52449:data<=-16'd3660;
      52450:data<=-16'd3303;
      52451:data<=-16'd2435;
      52452:data<=-16'd2623;
      52453:data<=-16'd1861;
      52454:data<=16'd126;
      52455:data<=16'd38;
      52456:data<=16'd491;
      52457:data<=16'd1730;
      52458:data<=-16'd230;
      52459:data<=16'd2108;
      52460:data<=16'd11934;
      52461:data<=16'd16932;
      52462:data<=16'd15493;
      52463:data<=16'd15198;
      52464:data<=16'd14766;
      52465:data<=16'd14046;
      52466:data<=16'd15406;
      52467:data<=16'd15870;
      52468:data<=16'd14469;
      52469:data<=16'd13647;
      52470:data<=16'd13336;
      52471:data<=16'd12853;
      52472:data<=16'd13157;
      52473:data<=16'd13829;
      52474:data<=16'd13238;
      52475:data<=16'd12642;
      52476:data<=16'd12819;
      52477:data<=16'd12005;
      52478:data<=16'd11629;
      52479:data<=16'd12722;
      52480:data<=16'd12842;
      52481:data<=16'd11909;
      52482:data<=16'd10464;
      52483:data<=16'd8956;
      52484:data<=16'd9344;
      52485:data<=16'd10481;
      52486:data<=16'd10649;
      52487:data<=16'd10458;
      52488:data<=16'd9899;
      52489:data<=16'd9424;
      52490:data<=16'd9529;
      52491:data<=16'd10430;
      52492:data<=16'd11489;
      52493:data<=16'd10472;
      52494:data<=16'd9441;
      52495:data<=16'd9770;
      52496:data<=16'd8657;
      52497:data<=16'd9219;
      52498:data<=16'd11268;
      52499:data<=16'd9862;
      52500:data<=16'd9677;
      52501:data<=16'd8748;
      52502:data<=16'd391;
      52503:data<=-16'd4749;
      52504:data<=-16'd2458;
      52505:data<=-16'd2252;
      52506:data<=-16'd2696;
      52507:data<=-16'd1823;
      52508:data<=-16'd2543;
      52509:data<=-16'd1926;
      52510:data<=-16'd384;
      52511:data<=-16'd191;
      52512:data<=16'd237;
      52513:data<=16'd68;
      52514:data<=-16'd412;
      52515:data<=16'd162;
      52516:data<=16'd714;
      52517:data<=16'd1474;
      52518:data<=16'd1891;
      52519:data<=16'd1460;
      52520:data<=16'd1422;
      52521:data<=16'd1064;
      52522:data<=16'd1362;
      52523:data<=16'd3193;
      52524:data<=16'd3548;
      52525:data<=16'd2955;
      52526:data<=16'd3016;
      52527:data<=16'd2264;
      52528:data<=16'd2366;
      52529:data<=16'd4062;
      52530:data<=16'd4366;
      52531:data<=16'd4009;
      52532:data<=16'd4645;
      52533:data<=16'd4686;
      52534:data<=16'd4604;
      52535:data<=16'd5653;
      52536:data<=16'd5805;
      52537:data<=16'd5083;
      52538:data<=16'd5277;
      52539:data<=16'd4617;
      52540:data<=16'd3700;
      52541:data<=16'd4235;
      52542:data<=16'd3242;
      52543:data<=16'd3873;
      52544:data<=16'd10759;
      52545:data<=16'd16318;
      52546:data<=16'd16019;
      52547:data<=16'd14090;
      52548:data<=16'd11956;
      52549:data<=16'd11110;
      52550:data<=16'd11179;
      52551:data<=16'd9809;
      52552:data<=16'd9344;
      52553:data<=16'd8739;
      52554:data<=16'd6126;
      52555:data<=16'd5278;
      52556:data<=16'd5227;
      52557:data<=16'd4147;
      52558:data<=16'd4255;
      52559:data<=16'd3755;
      52560:data<=16'd1668;
      52561:data<=16'd481;
      52562:data<=16'd566;
      52563:data<=16'd878;
      52564:data<=16'd438;
      52565:data<=-16'd17;
      52566:data<=-16'd732;
      52567:data<=-16'd2667;
      52568:data<=-16'd2743;
      52569:data<=-16'd1756;
      52570:data<=-16'd2579;
      52571:data<=-16'd2490;
      52572:data<=-16'd2778;
      52573:data<=-16'd4535;
      52574:data<=-16'd4184;
      52575:data<=-16'd4256;
      52576:data<=-16'd5262;
      52577:data<=-16'd4423;
      52578:data<=-16'd4960;
      52579:data<=-16'd6457;
      52580:data<=-16'd6492;
      52581:data<=-16'd6869;
      52582:data<=-16'd7608;
      52583:data<=-16'd8426;
      52584:data<=-16'd8328;
      52585:data<=-16'd9265;
      52586:data<=-16'd16328;
      52587:data<=-16'd22738;
      52588:data<=-16'd22107;
      52589:data<=-16'd20733;
      52590:data<=-16'd20046;
      52591:data<=-16'd19634;
      52592:data<=-16'd21375;
      52593:data<=-16'd21176;
      52594:data<=-16'd19707;
      52595:data<=-16'd19682;
      52596:data<=-16'd18328;
      52597:data<=-16'd17785;
      52598:data<=-16'd19014;
      52599:data<=-16'd18503;
      52600:data<=-16'd17723;
      52601:data<=-16'd17159;
      52602:data<=-16'd15766;
      52603:data<=-16'd15693;
      52604:data<=-16'd16648;
      52605:data<=-16'd16710;
      52606:data<=-16'd15838;
      52607:data<=-16'd14882;
      52608:data<=-16'd14280;
      52609:data<=-16'd13502;
      52610:data<=-16'd13603;
      52611:data<=-16'd14736;
      52612:data<=-16'd14600;
      52613:data<=-16'd13825;
      52614:data<=-16'd13209;
      52615:data<=-16'd12187;
      52616:data<=-16'd12461;
      52617:data<=-16'd13503;
      52618:data<=-16'd13110;
      52619:data<=-16'd12228;
      52620:data<=-16'd11653;
      52621:data<=-16'd10862;
      52622:data<=-16'd10455;
      52623:data<=-16'd11712;
      52624:data<=-16'd12809;
      52625:data<=-16'd10939;
      52626:data<=-16'd9861;
      52627:data<=-16'd10232;
      52628:data<=-16'd4725;
      52629:data<=16'd2561;
      52630:data<=16'd2793;
      52631:data<=16'd1848;
      52632:data<=16'd4096;
      52633:data<=16'd4890;
      52634:data<=16'd4291;
      52635:data<=16'd3724;
      52636:data<=16'd2746;
      52637:data<=16'd2604;
      52638:data<=16'd2911;
      52639:data<=16'd2666;
      52640:data<=16'd2319;
      52641:data<=16'd2202;
      52642:data<=16'd2428;
      52643:data<=16'd2416;
      52644:data<=16'd2444;
      52645:data<=16'd2801;
      52646:data<=16'd2429;
      52647:data<=16'd2676;
      52648:data<=16'd4134;
      52649:data<=16'd4679;
      52650:data<=16'd4807;
      52651:data<=16'd4684;
      52652:data<=16'd3826;
      52653:data<=16'd4399;
      52654:data<=16'd6050;
      52655:data<=16'd6740;
      52656:data<=16'd6646;
      52657:data<=16'd6507;
      52658:data<=16'd6807;
      52659:data<=16'd6620;
      52660:data<=16'd6570;
      52661:data<=16'd7911;
      52662:data<=16'd8014;
      52663:data<=16'd7632;
      52664:data<=16'd8232;
      52665:data<=16'd7256;
      52666:data<=16'd7597;
      52667:data<=16'd9359;
      52668:data<=16'd8815;
      52669:data<=16'd9028;
      52670:data<=16'd5327;
      52671:data<=-16'd4232;
      52672:data<=-16'd5645;
      52673:data<=-16'd1249;
      52674:data<=-16'd2155;
      52675:data<=-16'd2499;
      52676:data<=-16'd1107;
      52677:data<=-16'd1929;
      52678:data<=-16'd1569;
      52679:data<=-16'd273;
      52680:data<=16'd617;
      52681:data<=16'd1048;
      52682:data<=16'd161;
      52683:data<=-16'd321;
      52684:data<=-16'd805;
      52685:data<=-16'd607;
      52686:data<=16'd1697;
      52687:data<=16'd2294;
      52688:data<=16'd1789;
      52689:data<=16'd2090;
      52690:data<=16'd1274;
      52691:data<=16'd2036;
      52692:data<=16'd4346;
      52693:data<=16'd4642;
      52694:data<=16'd4278;
      52695:data<=16'd3779;
      52696:data<=16'd3297;
      52697:data<=16'd4017;
      52698:data<=16'd5133;
      52699:data<=16'd5859;
      52700:data<=16'd5043;
      52701:data<=16'd4337;
      52702:data<=16'd5166;
      52703:data<=16'd4755;
      52704:data<=16'd5083;
      52705:data<=16'd6815;
      52706:data<=16'd6479;
      52707:data<=16'd6276;
      52708:data<=16'd6000;
      52709:data<=16'd5225;
      52710:data<=16'd6258;
      52711:data<=16'd6294;
      52712:data<=16'd10000;
      52713:data<=16'd18973;
      52714:data<=16'd20339;
      52715:data<=16'd17014;
      52716:data<=16'd18513;
      52717:data<=16'd19147;
      52718:data<=16'd18161;
      52719:data<=16'd17958;
      52720:data<=16'd16716;
      52721:data<=16'd16304;
      52722:data<=16'd16158;
      52723:data<=16'd16010;
      52724:data<=16'd16612;
      52725:data<=16'd15380;
      52726:data<=16'd14407;
      52727:data<=16'd14222;
      52728:data<=16'd12586;
      52729:data<=16'd12895;
      52730:data<=16'd14183;
      52731:data<=16'd13373;
      52732:data<=16'd13076;
      52733:data<=16'd13453;
      52734:data<=16'd13173;
      52735:data<=16'd12971;
      52736:data<=16'd13668;
      52737:data<=16'd14295;
      52738:data<=16'd12737;
      52739:data<=16'd11617;
      52740:data<=16'd12160;
      52741:data<=16'd11257;
      52742:data<=16'd10698;
      52743:data<=16'd10784;
      52744:data<=16'd9441;
      52745:data<=16'd8734;
      52746:data<=16'd8411;
      52747:data<=16'd7691;
      52748:data<=16'd6331;
      52749:data<=16'd4384;
      52750:data<=16'd5109;
      52751:data<=16'd4811;
      52752:data<=16'd2640;
      52753:data<=16'd4535;
      52754:data<=16'd644;
      52755:data<=-16'd10930;
      52756:data<=-16'd13402;
      52757:data<=-16'd10796;
      52758:data<=-16'd12137;
      52759:data<=-16'd11233;
      52760:data<=-16'd10887;
      52761:data<=-16'd13312;
      52762:data<=-16'd13016;
      52763:data<=-16'd12381;
      52764:data<=-16'd12333;
      52765:data<=-16'd11060;
      52766:data<=-16'd11224;
      52767:data<=-16'd12446;
      52768:data<=-16'd12654;
      52769:data<=-16'd11994;
      52770:data<=-16'd11133;
      52771:data<=-16'd10886;
      52772:data<=-16'd11103;
      52773:data<=-16'd11815;
      52774:data<=-16'd12357;
      52775:data<=-16'd11885;
      52776:data<=-16'd11819;
      52777:data<=-16'd11447;
      52778:data<=-16'd10358;
      52779:data<=-16'd11169;
      52780:data<=-16'd12381;
      52781:data<=-16'd12003;
      52782:data<=-16'd12181;
      52783:data<=-16'd12868;
      52784:data<=-16'd12634;
      52785:data<=-16'd12662;
      52786:data<=-16'd13767;
      52787:data<=-16'd14029;
      52788:data<=-16'd12927;
      52789:data<=-16'd12642;
      52790:data<=-16'd12091;
      52791:data<=-16'd11270;
      52792:data<=-16'd13159;
      52793:data<=-16'd13744;
      52794:data<=-16'd12223;
      52795:data<=-16'd13470;
      52796:data<=-16'd9661;
      52797:data<=16'd899;
      52798:data<=16'd3178;
      52799:data<=-16'd1040;
      52800:data<=-16'd629;
      52801:data<=16'd136;
      52802:data<=-16'd417;
      52803:data<=16'd966;
      52804:data<=16'd517;
      52805:data<=-16'd1509;
      52806:data<=-16'd1671;
      52807:data<=-16'd1504;
      52808:data<=-16'd1510;
      52809:data<=-16'd1110;
      52810:data<=-16'd1544;
      52811:data<=-16'd2930;
      52812:data<=-16'd3865;
      52813:data<=-16'd3398;
      52814:data<=-16'd2626;
      52815:data<=-16'd2784;
      52816:data<=-16'd3247;
      52817:data<=-16'd3786;
      52818:data<=-16'd4282;
      52819:data<=-16'd4100;
      52820:data<=-16'd3682;
      52821:data<=-16'd3253;
      52822:data<=-16'd2696;
      52823:data<=-16'd3039;
      52824:data<=-16'd4397;
      52825:data<=-16'd4673;
      52826:data<=-16'd3538;
      52827:data<=-16'd3298;
      52828:data<=-16'd3368;
      52829:data<=-16'd3045;
      52830:data<=-16'd4429;
      52831:data<=-16'd5160;
      52832:data<=-16'd3422;
      52833:data<=-16'd2299;
      52834:data<=-16'd1475;
      52835:data<=-16'd1898;
      52836:data<=-16'd3510;
      52837:data<=-16'd1970;
      52838:data<=-16'd4566;
      52839:data<=-16'd14061;
      52840:data<=-16'd16545;
      52841:data<=-16'd13549;
      52842:data<=-16'd13994;
      52843:data<=-16'd13204;
      52844:data<=-16'd11985;
      52845:data<=-16'd12354;
      52846:data<=-16'd11068;
      52847:data<=-16'd10936;
      52848:data<=-16'd10448;
      52849:data<=-16'd7486;
      52850:data<=-16'd6701;
      52851:data<=-16'd6264;
      52852:data<=-16'd5265;
      52853:data<=-16'd6173;
      52854:data<=-16'd4996;
      52855:data<=-16'd2535;
      52856:data<=-16'd2457;
      52857:data<=-16'd1773;
      52858:data<=-16'd661;
      52859:data<=-16'd1368;
      52860:data<=-16'd1162;
      52861:data<=16'd934;
      52862:data<=16'd1683;
      52863:data<=16'd910;
      52864:data<=16'd1165;
      52865:data<=16'd1353;
      52866:data<=16'd1274;
      52867:data<=16'd2675;
      52868:data<=16'd3247;
      52869:data<=16'd3112;
      52870:data<=16'd3908;
      52871:data<=16'd3495;
      52872:data<=16'd3174;
      52873:data<=16'd4159;
      52874:data<=16'd5180;
      52875:data<=16'd6284;
      52876:data<=16'd5662;
      52877:data<=16'd5480;
      52878:data<=16'd6438;
      52879:data<=16'd4913;
      52880:data<=16'd9489;
      52881:data<=16'd20233;
      52882:data<=16'd21413;
      52883:data<=16'd17390;
      52884:data<=16'd17453;
      52885:data<=16'd17023;
      52886:data<=16'd17579;
      52887:data<=16'd18621;
      52888:data<=16'd16918;
      52889:data<=16'd16703;
      52890:data<=16'd16336;
      52891:data<=16'd14721;
      52892:data<=16'd15729;
      52893:data<=16'd16515;
      52894:data<=16'd15978;
      52895:data<=16'd15659;
      52896:data<=16'd14240;
      52897:data<=16'd13226;
      52898:data<=16'd13782;
      52899:data<=16'd14603;
      52900:data<=16'd14386;
      52901:data<=16'd13157;
      52902:data<=16'd12962;
      52903:data<=16'd12922;
      52904:data<=16'd12593;
      52905:data<=16'd13664;
      52906:data<=16'd13787;
      52907:data<=16'd12707;
      52908:data<=16'd12302;
      52909:data<=16'd11714;
      52910:data<=16'd11761;
      52911:data<=16'd12091;
      52912:data<=16'd11940;
      52913:data<=16'd11991;
      52914:data<=16'd10840;
      52915:data<=16'd9979;
      52916:data<=16'd9908;
      52917:data<=16'd9461;
      52918:data<=16'd11273;
      52919:data<=16'd11307;
      52920:data<=16'd8724;
      52921:data<=16'd9947;
      52922:data<=16'd6619;
      52923:data<=-16'd3139;
      52924:data<=-16'd5178;
      52925:data<=-16'd3022;
      52926:data<=-16'd4103;
      52927:data<=-16'd3774;
      52928:data<=-16'd3530;
      52929:data<=-16'd3768;
      52930:data<=-16'd1983;
      52931:data<=-16'd1730;
      52932:data<=-16'd1911;
      52933:data<=-16'd238;
      52934:data<=16'd167;
      52935:data<=-16'd182;
      52936:data<=16'd940;
      52937:data<=16'd2117;
      52938:data<=16'd1801;
      52939:data<=16'd936;
      52940:data<=16'd1068;
      52941:data<=16'd1627;
      52942:data<=16'd1670;
      52943:data<=16'd1254;
      52944:data<=16'd488;
      52945:data<=-16'd158;
      52946:data<=-16'd196;
      52947:data<=16'd215;
      52948:data<=-16'd617;
      52949:data<=-16'd2779;
      52950:data<=-16'd3286;
      52951:data<=-16'd3265;
      52952:data<=-16'd4176;
      52953:data<=-16'd3430;
      52954:data<=-16'd3433;
      52955:data<=-16'd5297;
      52956:data<=-16'd5054;
      52957:data<=-16'd4872;
      52958:data<=-16'd5783;
      52959:data<=-16'd5369;
      52960:data<=-16'd5703;
      52961:data<=-16'd5849;
      52962:data<=-16'd5953;
      52963:data<=-16'd8257;
      52964:data<=-16'd4974;
      52965:data<=16'd4525;
      52966:data<=16'd8019;
      52967:data<=16'd5542;
      52968:data<=16'd3983;
      52969:data<=16'd3077;
      52970:data<=16'd2955;
      52971:data<=16'd3450;
      52972:data<=16'd2933;
      52973:data<=16'd1924;
      52974:data<=16'd523;
      52975:data<=-16'd328;
      52976:data<=-16'd44;
      52977:data<=-16'd290;
      52978:data<=-16'd343;
      52979:data<=-16'd566;
      52980:data<=-16'd2689;
      52981:data<=-16'd3789;
      52982:data<=-16'd3597;
      52983:data<=-16'd5215;
      52984:data<=-16'd6214;
      52985:data<=-16'd5275;
      52986:data<=-16'd5843;
      52987:data<=-16'd7506;
      52988:data<=-16'd7653;
      52989:data<=-16'd6953;
      52990:data<=-16'd6440;
      52991:data<=-16'd6115;
      52992:data<=-16'd6936;
      52993:data<=-16'd8299;
      52994:data<=-16'd8087;
      52995:data<=-16'd7809;
      52996:data<=-16'd8358;
      52997:data<=-16'd7664;
      52998:data<=-16'd7689;
      52999:data<=-16'd9206;
      53000:data<=-16'd9160;
      53001:data<=-16'd8630;
      53002:data<=-16'd8338;
      53003:data<=-16'd7818;
      53004:data<=-16'd8038;
      53005:data<=-16'd7756;
      53006:data<=-16'd10959;
      53007:data<=-16'd19643;
      53008:data<=-16'd23335;
      53009:data<=-16'd20812;
      53010:data<=-16'd20086;
      53011:data<=-16'd20190;
      53012:data<=-16'd20369;
      53013:data<=-16'd20706;
      53014:data<=-16'd19108;
      53015:data<=-16'd18075;
      53016:data<=-16'd17643;
      53017:data<=-16'd17097;
      53018:data<=-16'd17952;
      53019:data<=-16'd17327;
      53020:data<=-16'd16029;
      53021:data<=-16'd16096;
      53022:data<=-16'd14624;
      53023:data<=-16'd13897;
      53024:data<=-16'd14957;
      53025:data<=-16'd14184;
      53026:data<=-16'd13420;
      53027:data<=-16'd13433;
      53028:data<=-16'd12427;
      53029:data<=-16'd11913;
      53030:data<=-16'd12592;
      53031:data<=-16'd13221;
      53032:data<=-16'd12210;
      53033:data<=-16'd10213;
      53034:data<=-16'd9313;
      53035:data<=-16'd8674;
      53036:data<=-16'd8595;
      53037:data<=-16'd9450;
      53038:data<=-16'd9092;
      53039:data<=-16'd8238;
      53040:data<=-16'd7893;
      53041:data<=-16'd7756;
      53042:data<=-16'd7400;
      53043:data<=-16'd6041;
      53044:data<=-16'd5768;
      53045:data<=-16'd5456;
      53046:data<=-16'd4088;
      53047:data<=-16'd5542;
      53048:data<=-16'd2625;
      53049:data<=16'd8153;
      53050:data<=16'd12792;
      53051:data<=16'd10980;
      53052:data<=16'd11356;
      53053:data<=16'd10634;
      53054:data<=16'd9559;
      53055:data<=16'd10931;
      53056:data<=16'd11828;
      53057:data<=16'd12000;
      53058:data<=16'd11629;
      53059:data<=16'd11239;
      53060:data<=16'd11341;
      53061:data<=16'd11179;
      53062:data<=16'd12160;
      53063:data<=16'd12545;
      53064:data<=16'd11450;
      53065:data<=16'd11609;
      53066:data<=16'd11201;
      53067:data<=16'd10921;
      53068:data<=16'd12225;
      53069:data<=16'd11897;
      53070:data<=16'd11896;
      53071:data<=16'd12372;
      53072:data<=16'd10833;
      53073:data<=16'd11257;
      53074:data<=16'd12795;
      53075:data<=16'd12232;
      53076:data<=16'd12094;
      53077:data<=16'd12290;
      53078:data<=16'd11715;
      53079:data<=16'd10757;
      53080:data<=16'd10674;
      53081:data<=16'd12528;
      53082:data<=16'd12627;
      53083:data<=16'd10853;
      53084:data<=16'd9943;
      53085:data<=16'd8611;
      53086:data<=16'd9127;
      53087:data<=16'd10549;
      53088:data<=16'd9862;
      53089:data<=16'd11053;
      53090:data<=16'd8805;
      53091:data<=-16'd519;
      53092:data<=-16'd4249;
      53093:data<=-16'd1560;
      53094:data<=-16'd981;
      53095:data<=-16'd802;
      53096:data<=-16'd611;
      53097:data<=-16'd1287;
      53098:data<=-16'd720;
      53099:data<=16'd631;
      53100:data<=16'd1945;
      53101:data<=16'd1956;
      53102:data<=16'd1089;
      53103:data<=16'd1445;
      53104:data<=16'd1491;
      53105:data<=16'd1713;
      53106:data<=16'd3248;
      53107:data<=16'd3385;
      53108:data<=16'd2936;
      53109:data<=16'd3328;
      53110:data<=16'd3324;
      53111:data<=16'd3788;
      53112:data<=16'd4451;
      53113:data<=16'd4144;
      53114:data<=16'd3756;
      53115:data<=16'd3453;
      53116:data<=16'd3269;
      53117:data<=16'd3771;
      53118:data<=16'd4852;
      53119:data<=16'd5297;
      53120:data<=16'd4434;
      53121:data<=16'd4322;
      53122:data<=16'd4758;
      53123:data<=16'd4027;
      53124:data<=16'd4469;
      53125:data<=16'd5568;
      53126:data<=16'd5140;
      53127:data<=16'd5368;
      53128:data<=16'd5162;
      53129:data<=16'd3980;
      53130:data<=16'd5124;
      53131:data<=16'd5991;
      53132:data<=16'd7532;
      53133:data<=16'd15104;
      53134:data<=16'd21006;
      53135:data<=16'd19384;
      53136:data<=16'd18550;
      53137:data<=16'd20198;
      53138:data<=16'd19620;
      53139:data<=16'd18334;
      53140:data<=16'd17438;
      53141:data<=16'd16568;
      53142:data<=16'd16252;
      53143:data<=16'd15138;
      53144:data<=16'd13756;
      53145:data<=16'd13110;
      53146:data<=16'd11734;
      53147:data<=16'd10848;
      53148:data<=16'd11145;
      53149:data<=16'd9923;
      53150:data<=16'd8038;
      53151:data<=16'd7389;
      53152:data<=16'd6405;
      53153:data<=16'd5653;
      53154:data<=16'd6269;
      53155:data<=16'd5330;
      53156:data<=16'd2914;
      53157:data<=16'd2500;
      53158:data<=16'd2554;
      53159:data<=16'd1592;
      53160:data<=16'd1726;
      53161:data<=16'd1412;
      53162:data<=-16'd282;
      53163:data<=-16'd936;
      53164:data<=-16'd1575;
      53165:data<=-16'd2444;
      53166:data<=-16'd1867;
      53167:data<=-16'd1803;
      53168:data<=-16'd3156;
      53169:data<=-16'd4077;
      53170:data<=-16'd4015;
      53171:data<=-16'd4091;
      53172:data<=-16'd4555;
      53173:data<=-16'd3891;
      53174:data<=-16'd6334;
      53175:data<=-16'd15004;
      53176:data<=-16'd20014;
      53177:data<=-16'd18437;
      53178:data<=-16'd18104;
      53179:data<=-16'd17758;
      53180:data<=-16'd17288;
      53181:data<=-16'd19074;
      53182:data<=-16'd18480;
      53183:data<=-16'd17854;
      53184:data<=-16'd19570;
      53185:data<=-16'd18545;
      53186:data<=-16'd17769;
      53187:data<=-16'd19018;
      53188:data<=-16'd18269;
      53189:data<=-16'd17705;
      53190:data<=-16'd17609;
      53191:data<=-16'd16290;
      53192:data<=-16'd16211;
      53193:data<=-16'd17071;
      53194:data<=-16'd17302;
      53195:data<=-16'd16707;
      53196:data<=-16'd15816;
      53197:data<=-16'd15666;
      53198:data<=-16'd14844;
      53199:data<=-16'd14372;
      53200:data<=-16'd15673;
      53201:data<=-16'd15241;
      53202:data<=-16'd13907;
      53203:data<=-16'd13899;
      53204:data<=-16'd12866;
      53205:data<=-16'd12223;
      53206:data<=-16'd13186;
      53207:data<=-16'd13088;
      53208:data<=-16'd12302;
      53209:data<=-16'd11913;
      53210:data<=-16'd11409;
      53211:data<=-16'd11320;
      53212:data<=-16'd12290;
      53213:data<=-16'd12674;
      53214:data<=-16'd11239;
      53215:data<=-16'd10827;
      53216:data<=-16'd9432;
      53217:data<=-16'd2179;
      53218:data<=16'd3626;
      53219:data<=16'd2833;
      53220:data<=16'd2332;
      53221:data<=16'd2660;
      53222:data<=16'd1765;
      53223:data<=16'd2379;
      53224:data<=16'd2594;
      53225:data<=16'd1342;
      53226:data<=16'd936;
      53227:data<=16'd490;
      53228:data<=16'd140;
      53229:data<=16'd784;
      53230:data<=16'd526;
      53231:data<=-16'd1107;
      53232:data<=-16'd1557;
      53233:data<=16'd135;
      53234:data<=16'd1481;
      53235:data<=16'd1757;
      53236:data<=16'd1448;
      53237:data<=-16'd311;
      53238:data<=-16'd910;
      53239:data<=16'd520;
      53240:data<=16'd281;
      53241:data<=-16'd553;
      53242:data<=-16'd375;
      53243:data<=-16'd385;
      53244:data<=16'd167;
      53245:data<=16'd604;
      53246:data<=16'd913;
      53247:data<=16'd1483;
      53248:data<=16'd528;
      53249:data<=16'd896;
      53250:data<=16'd3033;
      53251:data<=16'd3043;
      53252:data<=16'd3526;
      53253:data<=16'd4349;
      53254:data<=16'd3146;
      53255:data<=16'd3808;
      53256:data<=16'd5304;
      53257:data<=16'd5547;
      53258:data<=16'd5122;
      53259:data<=-16'd441;
      53260:data<=-16'd7439;
      53261:data<=-16'd7712;
      53262:data<=-16'd5551;
      53263:data<=-16'd4488;
      53264:data<=-16'd2999;
      53265:data<=-16'd2783;
      53266:data<=-16'd3353;
      53267:data<=-16'd3162;
      53268:data<=-16'd2220;
      53269:data<=-16'd505;
      53270:data<=16'd426;
      53271:data<=16'd523;
      53272:data<=16'd437;
      53273:data<=16'd9;
      53274:data<=16'd1098;
      53275:data<=16'd2972;
      53276:data<=16'd3503;
      53277:data<=16'd3879;
      53278:data<=16'd3892;
      53279:data<=16'd3122;
      53280:data<=16'd3233;
      53281:data<=16'd4476;
      53282:data<=16'd5862;
      53283:data<=16'd5614;
      53284:data<=16'd3932;
      53285:data<=16'd3389;
      53286:data<=16'd3674;
      53287:data<=16'd4264;
      53288:data<=16'd5316;
      53289:data<=16'd5151;
      53290:data<=16'd4907;
      53291:data<=16'd5777;
      53292:data<=16'd6100;
      53293:data<=16'd6637;
      53294:data<=16'd7780;
      53295:data<=16'd8023;
      53296:data<=16'd7450;
      53297:data<=16'd6561;
      53298:data<=16'd6287;
      53299:data<=16'd6441;
      53300:data<=16'd7624;
      53301:data<=16'd13860;
      53302:data<=16'd21291;
      53303:data<=16'd21552;
      53304:data<=16'd19039;
      53305:data<=16'd19816;
      53306:data<=16'd20306;
      53307:data<=16'd19738;
      53308:data<=16'd19808;
      53309:data<=16'd18480;
      53310:data<=16'd16669;
      53311:data<=16'd16483;
      53312:data<=16'd16237;
      53313:data<=16'd15644;
      53314:data<=16'd15559;
      53315:data<=16'd15097;
      53316:data<=16'd14499;
      53317:data<=16'd13749;
      53318:data<=16'd12939;
      53319:data<=16'd13917;
      53320:data<=16'd14628;
      53321:data<=16'd13261;
      53322:data<=16'd13057;
      53323:data<=16'd13079;
      53324:data<=16'd11938;
      53325:data<=16'd12596;
      53326:data<=16'd12798;
      53327:data<=16'd11095;
      53328:data<=16'd10627;
      53329:data<=16'd10138;
      53330:data<=16'd10442;
      53331:data<=16'd12730;
      53332:data<=16'd12228;
      53333:data<=16'd10693;
      53334:data<=16'd11700;
      53335:data<=16'd11546;
      53336:data<=16'd10713;
      53337:data<=16'd11135;
      53338:data<=16'd11091;
      53339:data<=16'd11022;
      53340:data<=16'd10081;
      53341:data<=16'd9021;
      53342:data<=16'd9392;
      53343:data<=16'd5081;
      53344:data<=-16'd2940;
      53345:data<=-16'd5285;
      53346:data<=-16'd4538;
      53347:data<=-16'd5413;
      53348:data<=-16'd5004;
      53349:data<=-16'd4819;
      53350:data<=-16'd6429;
      53351:data<=-16'd7004;
      53352:data<=-16'd6771;
      53353:data<=-16'd6558;
      53354:data<=-16'd6225;
      53355:data<=-16'd6907;
      53356:data<=-16'd8414;
      53357:data<=-16'd9394;
      53358:data<=-16'd9200;
      53359:data<=-16'd8625;
      53360:data<=-16'd8440;
      53361:data<=-16'd7718;
      53362:data<=-16'd7407;
      53363:data<=-16'd8687;
      53364:data<=-16'd9520;
      53365:data<=-16'd9605;
      53366:data<=-16'd9441;
      53367:data<=-16'd8223;
      53368:data<=-16'd7595;
      53369:data<=-16'd8102;
      53370:data<=-16'd8357;
      53371:data<=-16'd8913;
      53372:data<=-16'd9354;
      53373:data<=-16'd8825;
      53374:data<=-16'd8590;
      53375:data<=-16'd9444;
      53376:data<=-16'd10516;
      53377:data<=-16'd10686;
      53378:data<=-16'd10326;
      53379:data<=-16'd9529;
      53380:data<=-16'd8796;
      53381:data<=-16'd10302;
      53382:data<=-16'd11195;
      53383:data<=-16'd10366;
      53384:data<=-16'd11914;
      53385:data<=-16'd8977;
      53386:data<=16'd519;
      53387:data<=16'd2535;
      53388:data<=-16'd969;
      53389:data<=-16'd329;
      53390:data<=-16'd870;
      53391:data<=-16'd1847;
      53392:data<=-16'd144;
      53393:data<=-16'd1683;
      53394:data<=-16'd4084;
      53395:data<=-16'd3739;
      53396:data<=-16'd4137;
      53397:data<=-16'd4067;
      53398:data<=-16'd2928;
      53399:data<=-16'd3723;
      53400:data<=-16'd5344;
      53401:data<=-16'd5821;
      53402:data<=-16'd5629;
      53403:data<=-16'd5251;
      53404:data<=-16'd4502;
      53405:data<=-16'd4476;
      53406:data<=-16'd6158;
      53407:data<=-16'd7272;
      53408:data<=-16'd6761;
      53409:data<=-16'd6322;
      53410:data<=-16'd6034;
      53411:data<=-16'd5662;
      53412:data<=-16'd5899;
      53413:data<=-16'd7092;
      53414:data<=-16'd8064;
      53415:data<=-16'd7376;
      53416:data<=-16'd6701;
      53417:data<=-16'd6824;
      53418:data<=-16'd7059;
      53419:data<=-16'd8290;
      53420:data<=-16'd8643;
      53421:data<=-16'd7911;
      53422:data<=-16'd8108;
      53423:data<=-16'd6987;
      53424:data<=-16'd6555;
      53425:data<=-16'd8229;
      53426:data<=-16'd7576;
      53427:data<=-16'd9999;
      53428:data<=-16'd17515;
      53429:data<=-16'd19241;
      53430:data<=-16'd16712;
      53431:data<=-16'd17406;
      53432:data<=-16'd17981;
      53433:data<=-16'd17179;
      53434:data<=-16'd17004;
      53435:data<=-16'd16049;
      53436:data<=-16'd14475;
      53437:data<=-16'd14744;
      53438:data<=-16'd16362;
      53439:data<=-16'd15858;
      53440:data<=-16'd13870;
      53441:data<=-16'd13241;
      53442:data<=-16'd12969;
      53443:data<=-16'd12897;
      53444:data<=-16'd12848;
      53445:data<=-16'd11418;
      53446:data<=-16'd10430;
      53447:data<=-16'd10117;
      53448:data<=-16'd9341;
      53449:data<=-16'd8381;
      53450:data<=-16'd6502;
      53451:data<=-16'd5600;
      53452:data<=-16'd5802;
      53453:data<=-16'd4297;
      53454:data<=-16'd3864;
      53455:data<=-16'd4391;
      53456:data<=-16'd2541;
      53457:data<=-16'd1190;
      53458:data<=-16'd887;
      53459:data<=-16'd306;
      53460:data<=-16'd814;
      53461:data<=-16'd758;
      53462:data<=16'd617;
      53463:data<=16'd2182;
      53464:data<=16'd3124;
      53465:data<=16'd2484;
      53466:data<=16'd2874;
      53467:data<=16'd3275;
      53468:data<=16'd1888;
      53469:data<=16'd6357;
      53470:data<=16'd14815;
      53471:data<=16'd16360;
      53472:data<=16'd14651;
      53473:data<=16'd14959;
      53474:data<=16'd14569;
      53475:data<=16'd14895;
      53476:data<=16'd15719;
      53477:data<=16'd14569;
      53478:data<=16'd14092;
      53479:data<=16'd14317;
      53480:data<=16'd13182;
      53481:data<=16'd12974;
      53482:data<=16'd13888;
      53483:data<=16'd13643;
      53484:data<=16'd13396;
      53485:data<=16'd13239;
      53486:data<=16'd11931;
      53487:data<=16'd12029;
      53488:data<=16'd13364;
      53489:data<=16'd12645;
      53490:data<=16'd11931;
      53491:data<=16'd12088;
      53492:data<=16'd10934;
      53493:data<=16'd11341;
      53494:data<=16'd13189;
      53495:data<=16'd12135;
      53496:data<=16'd10821;
      53497:data<=16'd11723;
      53498:data<=16'd11735;
      53499:data<=16'd10998;
      53500:data<=16'd11350;
      53501:data<=16'd11565;
      53502:data<=16'd10983;
      53503:data<=16'd10787;
      53504:data<=16'd10574;
      53505:data<=16'd9133;
      53506:data<=16'd9242;
      53507:data<=16'd11825;
      53508:data<=16'd11473;
      53509:data<=16'd9409;
      53510:data<=16'd9875;
      53511:data<=16'd6598;
      53512:data<=-16'd576;
      53513:data<=-16'd1885;
      53514:data<=16'd234;
      53515:data<=-16'd613;
      53516:data<=-16'd1389;
      53517:data<=-16'd1115;
      53518:data<=-16'd828;
      53519:data<=16'd644;
      53520:data<=16'd1403;
      53521:data<=16'd822;
      53522:data<=16'd1134;
      53523:data<=16'd1438;
      53524:data<=16'd928;
      53525:data<=16'd1554;
      53526:data<=16'd2898;
      53527:data<=16'd2783;
      53528:data<=16'd2391;
      53529:data<=16'd2689;
      53530:data<=16'd2033;
      53531:data<=16'd2096;
      53532:data<=16'd3712;
      53533:data<=16'd3607;
      53534:data<=16'd2961;
      53535:data<=16'd3154;
      53536:data<=16'd2085;
      53537:data<=16'd2020;
      53538:data<=16'd3764;
      53539:data<=16'd3946;
      53540:data<=16'd3127;
      53541:data<=16'd3268;
      53542:data<=16'd4578;
      53543:data<=16'd5015;
      53544:data<=16'd2907;
      53545:data<=16'd2077;
      53546:data<=16'd3328;
      53547:data<=16'd2863;
      53548:data<=16'd1629;
      53549:data<=16'd1028;
      53550:data<=16'd829;
      53551:data<=16'd106;
      53552:data<=-16'd2036;
      53553:data<=16'd187;
      53554:data<=16'd7297;
      53555:data<=16'd9498;
      53556:data<=16'd7060;
      53557:data<=16'd6258;
      53558:data<=16'd6143;
      53559:data<=16'd5513;
      53560:data<=16'd4993;
      53561:data<=16'd5121;
      53562:data<=16'd4654;
      53563:data<=16'd2137;
      53564:data<=16'd1030;
      53565:data<=16'd1535;
      53566:data<=16'd732;
      53567:data<=16'd720;
      53568:data<=16'd726;
      53569:data<=-16'd851;
      53570:data<=-16'd1401;
      53571:data<=-16'd1795;
      53572:data<=-16'd2692;
      53573:data<=-16'd2413;
      53574:data<=-16'd2027;
      53575:data<=-16'd3016;
      53576:data<=-16'd5260;
      53577:data<=-16'd5799;
      53578:data<=-16'd4507;
      53579:data<=-16'd5110;
      53580:data<=-16'd4946;
      53581:data<=-16'd3889;
      53582:data<=-16'd5930;
      53583:data<=-16'd6725;
      53584:data<=-16'd6187;
      53585:data<=-16'd7286;
      53586:data<=-16'd5692;
      53587:data<=-16'd4481;
      53588:data<=-16'd6880;
      53589:data<=-16'd7360;
      53590:data<=-16'd6396;
      53591:data<=-16'd5846;
      53592:data<=-16'd5527;
      53593:data<=-16'd6173;
      53594:data<=-16'd5603;
      53595:data<=-16'd8216;
      53596:data<=-16'd16089;
      53597:data<=-16'd19021;
      53598:data<=-16'd17076;
      53599:data<=-16'd16926;
      53600:data<=-16'd16948;
      53601:data<=-16'd17274;
      53602:data<=-16'd17368;
      53603:data<=-16'd15781;
      53604:data<=-16'd15329;
      53605:data<=-16'd15126;
      53606:data<=-16'd15032;
      53607:data<=-16'd16237;
      53608:data<=-16'd15380;
      53609:data<=-16'd13958;
      53610:data<=-16'd13979;
      53611:data<=-16'd12565;
      53612:data<=-16'd11779;
      53613:data<=-16'd12888;
      53614:data<=-16'd13006;
      53615:data<=-16'd12630;
      53616:data<=-16'd12295;
      53617:data<=-16'd11665;
      53618:data<=-16'd11298;
      53619:data<=-16'd11497;
      53620:data<=-16'd12656;
      53621:data<=-16'd12678;
      53622:data<=-16'd11016;
      53623:data<=-16'd10610;
      53624:data<=-16'd10448;
      53625:data<=-16'd9993;
      53626:data<=-16'd10995;
      53627:data<=-16'd10981;
      53628:data<=-16'd9658;
      53629:data<=-16'd9382;
      53630:data<=-16'd8851;
      53631:data<=-16'd8316;
      53632:data<=-16'd9291;
      53633:data<=-16'd9988;
      53634:data<=-16'd9232;
      53635:data<=-16'd8669;
      53636:data<=-16'd8739;
      53637:data<=-16'd5741;
      53638:data<=16'd443;
      53639:data<=16'd3310;
      53640:data<=16'd2854;
      53641:data<=16'd3395;
      53642:data<=16'd3081;
      53643:data<=16'd2466;
      53644:data<=16'd3818;
      53645:data<=16'd3902;
      53646:data<=16'd3218;
      53647:data<=16'd4410;
      53648:data<=16'd4373;
      53649:data<=16'd2836;
      53650:data<=16'd3712;
      53651:data<=16'd6229;
      53652:data<=16'd7262;
      53653:data<=16'd7212;
      53654:data<=16'd7257;
      53655:data<=16'd6971;
      53656:data<=16'd7636;
      53657:data<=16'd9653;
      53658:data<=16'd9712;
      53659:data<=16'd8554;
      53660:data<=16'd9121;
      53661:data<=16'd8845;
      53662:data<=16'd7580;
      53663:data<=16'd8830;
      53664:data<=16'd10486;
      53665:data<=16'd10084;
      53666:data<=16'd9750;
      53667:data<=16'd9935;
      53668:data<=16'd9803;
      53669:data<=16'd10649;
      53670:data<=16'd12000;
      53671:data<=16'd11502;
      53672:data<=16'd10355;
      53673:data<=16'd10296;
      53674:data<=16'd10266;
      53675:data<=16'd10912;
      53676:data<=16'd11888;
      53677:data<=16'd11729;
      53678:data<=16'd12190;
      53679:data<=16'd9955;
      53680:data<=16'd2760;
      53681:data<=-16'd391;
      53682:data<=16'd1107;
      53683:data<=16'd130;
      53684:data<=16'd61;
      53685:data<=16'd1325;
      53686:data<=16'd58;
      53687:data<=16'd270;
      53688:data<=16'd2393;
      53689:data<=16'd3239;
      53690:data<=16'd3726;
      53691:data<=16'd3521;
      53692:data<=16'd2961;
      53693:data<=16'd2998;
      53694:data<=16'd3200;
      53695:data<=16'd4695;
      53696:data<=16'd5767;
      53697:data<=16'd4475;
      53698:data<=16'd3618;
      53699:data<=16'd4199;
      53700:data<=16'd4777;
      53701:data<=16'd4554;
      53702:data<=16'd4293;
      53703:data<=16'd5385;
      53704:data<=16'd5883;
      53705:data<=16'd5529;
      53706:data<=16'd6382;
      53707:data<=16'd6607;
      53708:data<=16'd6452;
      53709:data<=16'd7282;
      53710:data<=16'd6959;
      53711:data<=16'd6114;
      53712:data<=16'd5841;
      53713:data<=16'd6152;
      53714:data<=16'd7999;
      53715:data<=16'd8900;
      53716:data<=16'd7771;
      53717:data<=16'd7031;
      53718:data<=16'd7166;
      53719:data<=16'd7932;
      53720:data<=16'd8684;
      53721:data<=16'd11462;
      53722:data<=16'd17282;
      53723:data<=16'd19341;
      53724:data<=16'd17755;
      53725:data<=16'd18627;
      53726:data<=16'd18992;
      53727:data<=16'd18239;
      53728:data<=16'd18654;
      53729:data<=16'd17141;
      53730:data<=16'd15487;
      53731:data<=16'd16230;
      53732:data<=16'd16680;
      53733:data<=16'd16299;
      53734:data<=16'd15227;
      53735:data<=16'd14296;
      53736:data<=16'd14343;
      53737:data<=16'd13232;
      53738:data<=16'd12366;
      53739:data<=16'd13808;
      53740:data<=16'd14322;
      53741:data<=16'd12762;
      53742:data<=16'd12035;
      53743:data<=16'd12480;
      53744:data<=16'd11329;
      53745:data<=16'd9344;
      53746:data<=16'd9370;
      53747:data<=16'd9407;
      53748:data<=16'd8627;
      53749:data<=16'd8546;
      53750:data<=16'd6949;
      53751:data<=16'd4555;
      53752:data<=16'd4114;
      53753:data<=16'd3855;
      53754:data<=16'd2958;
      53755:data<=16'd2247;
      53756:data<=16'd1532;
      53757:data<=16'd390;
      53758:data<=-16'd787;
      53759:data<=-16'd602;
      53760:data<=-16'd1105;
      53761:data<=-16'd2059;
      53762:data<=-16'd96;
      53763:data<=-16'd2432;
      53764:data<=-16'd11615;
      53765:data<=-16'd15802;
      53766:data<=-16'd14797;
      53767:data<=-16'd15215;
      53768:data<=-16'd14803;
      53769:data<=-16'd14619;
      53770:data<=-16'd15884;
      53771:data<=-16'd15273;
      53772:data<=-16'd14254;
      53773:data<=-16'd14469;
      53774:data<=-16'd14387;
      53775:data<=-16'd14017;
      53776:data<=-16'd14085;
      53777:data<=-16'd14586;
      53778:data<=-16'd14628;
      53779:data<=-16'd13987;
      53780:data<=-16'd13324;
      53781:data<=-16'd13044;
      53782:data<=-16'd13709;
      53783:data<=-16'd14037;
      53784:data<=-16'd13426;
      53785:data<=-16'd13490;
      53786:data<=-16'd12724;
      53787:data<=-16'd11036;
      53788:data<=-16'd11608;
      53789:data<=-16'd13036;
      53790:data<=-16'd12809;
      53791:data<=-16'd11499;
      53792:data<=-16'd10272;
      53793:data<=-16'd10417;
      53794:data<=-16'd11210;
      53795:data<=-16'd11696;
      53796:data<=-16'd12395;
      53797:data<=-16'd11922;
      53798:data<=-16'd10310;
      53799:data<=-16'd10132;
      53800:data<=-16'd11136;
      53801:data<=-16'd11456;
      53802:data<=-16'd10937;
      53803:data<=-16'd10941;
      53804:data<=-16'd11179;
      53805:data<=-16'd8225;
      53806:data<=-16'd2685;
      53807:data<=-16'd188;
      53808:data<=-16'd840;
      53809:data<=-16'd711;
      53810:data<=-16'd567;
      53811:data<=-16'd863;
      53812:data<=16'd150;
      53813:data<=-16'd133;
      53814:data<=-16'd2021;
      53815:data<=-16'd1726;
      53816:data<=-16'd1403;
      53817:data<=-16'd2487;
      53818:data<=-16'd2435;
      53819:data<=-16'd3203;
      53820:data<=-16'd4548;
      53821:data<=-16'd4029;
      53822:data<=-16'd3864;
      53823:data<=-16'd3794;
      53824:data<=-16'd3427;
      53825:data<=-16'd4743;
      53826:data<=-16'd5597;
      53827:data<=-16'd5485;
      53828:data<=-16'd5829;
      53829:data<=-16'd5439;
      53830:data<=-16'd5136;
      53831:data<=-16'd5165;
      53832:data<=-16'd4996;
      53833:data<=-16'd5938;
      53834:data<=-16'd6311;
      53835:data<=-16'd5224;
      53836:data<=-16'd4672;
      53837:data<=-16'd4802;
      53838:data<=-16'd5489;
      53839:data<=-16'd5827;
      53840:data<=-16'd5524;
      53841:data<=-16'd6382;
      53842:data<=-16'd6834;
      53843:data<=-16'd5941;
      53844:data<=-16'd6190;
      53845:data<=-16'd6162;
      53846:data<=-16'd4278;
      53847:data<=-16'd4910;
      53848:data<=-16'd10317;
      53849:data<=-16'd14569;
      53850:data<=-16'd13709;
      53851:data<=-16'd11705;
      53852:data<=-16'd10334;
      53853:data<=-16'd8959;
      53854:data<=-16'd9327;
      53855:data<=-16'd9826;
      53856:data<=-16'd8611;
      53857:data<=-16'd6898;
      53858:data<=-16'd5221;
      53859:data<=-16'd5081;
      53860:data<=-16'd5162;
      53861:data<=-16'd3507;
      53862:data<=-16'd3322;
      53863:data<=-16'd3142;
      53864:data<=-16'd534;
      53865:data<=16'd259;
      53866:data<=-16'd488;
      53867:data<=-16'd156;
      53868:data<=16'd352;
      53869:data<=16'd1644;
      53870:data<=16'd3224;
      53871:data<=16'd3835;
      53872:data<=16'd3802;
      53873:data<=16'd3281;
      53874:data<=16'd3365;
      53875:data<=16'd3926;
      53876:data<=16'd4918;
      53877:data<=16'd6730;
      53878:data<=16'd6642;
      53879:data<=16'd5510;
      53880:data<=16'd5723;
      53881:data<=16'd5253;
      53882:data<=16'd5227;
      53883:data<=16'd6370;
      53884:data<=16'd6094;
      53885:data<=16'd5903;
      53886:data<=16'd6434;
      53887:data<=16'd6187;
      53888:data<=16'd6449;
      53889:data<=16'd8851;
      53890:data<=16'd13746;
      53891:data<=16'd17656;
      53892:data<=16'd17387;
      53893:data<=16'd16107;
      53894:data<=16'd16146;
      53895:data<=16'd16904;
      53896:data<=16'd17482;
      53897:data<=16'd16483;
      53898:data<=16'd15558;
      53899:data<=16'd15147;
      53900:data<=16'd13951;
      53901:data<=16'd14395;
      53902:data<=16'd15280;
      53903:data<=16'd13916;
      53904:data<=16'd13118;
      53905:data<=16'd12953;
      53906:data<=16'd12198;
      53907:data<=16'd12619;
      53908:data<=16'd12951;
      53909:data<=16'd12178;
      53910:data<=16'd11947;
      53911:data<=16'd11429;
      53912:data<=16'd10146;
      53913:data<=16'd10513;
      53914:data<=16'd12361;
      53915:data<=16'd12452;
      53916:data<=16'd11100;
      53917:data<=16'd10657;
      53918:data<=16'd10125;
      53919:data<=16'd9717;
      53920:data<=16'd11013;
      53921:data<=16'd11388;
      53922:data<=16'd9520;
      53923:data<=16'd8355;
      53924:data<=16'd8332;
      53925:data<=16'd7711;
      53926:data<=16'd7577;
      53927:data<=16'd9041;
      53928:data<=16'd9558;
      53929:data<=16'd8586;
      53930:data<=16'd8853;
      53931:data<=16'd7926;
      53932:data<=16'd2643;
      53933:data<=-16'd1955;
      53934:data<=-16'd1829;
      53935:data<=-16'd669;
      53936:data<=-16'd1110;
      53937:data<=-16'd1612;
      53938:data<=-16'd1491;
      53939:data<=-16'd628;
      53940:data<=16'd896;
      53941:data<=16'd908;
      53942:data<=-16'd270;
      53943:data<=16'd127;
      53944:data<=16'd840;
      53945:data<=16'd218;
      53946:data<=-16'd781;
      53947:data<=-16'd1579;
      53948:data<=-16'd1418;
      53949:data<=-16'd1240;
      53950:data<=-16'd2018;
      53951:data<=-16'd2273;
      53952:data<=-16'd2908;
      53953:data<=-16'd3987;
      53954:data<=-16'd3706;
      53955:data<=-16'd3586;
      53956:data<=-16'd3565;
      53957:data<=-16'd3428;
      53958:data<=-16'd4922;
      53959:data<=-16'd5655;
      53960:data<=-16'd5148;
      53961:data<=-16'd5691;
      53962:data<=-16'd5796;
      53963:data<=-16'd5821;
      53964:data<=-16'd7286;
      53965:data<=-16'd8555;
      53966:data<=-16'd8622;
      53967:data<=-16'd7665;
      53968:data<=-16'd6190;
      53969:data<=-16'd5630;
      53970:data<=-16'd9059;
      53971:data<=-16'd15023;
      53972:data<=-16'd16081;
      53973:data<=-16'd14637;
      53974:data<=-16'd15687;
      53975:data<=-16'd13755;
      53976:data<=-16'd12366;
      53977:data<=-16'd15923;
      53978:data<=-16'd11583;
      53979:data<=16'd3686;
      53980:data<=16'd14548;
      53981:data<=16'd12348;
      53982:data<=16'd5495;
      53983:data<=16'd4493;
      53984:data<=16'd4454;
      53985:data<=16'd2319;
      53986:data<=16'd3598;
      53987:data<=16'd2234;
      53988:data<=-16'd3395;
      53989:data<=-16'd5873;
      53990:data<=-16'd6508;
      53991:data<=-16'd5442;
      53992:data<=-16'd7894;
      53993:data<=-16'd17517;
      53994:data<=-16'd18971;
      53995:data<=-16'd13561;
      53996:data<=-16'd14051;
      53997:data<=-16'd13261;
      53998:data<=-16'd11353;
      53999:data<=-16'd12424;
      54000:data<=-16'd10613;
      54001:data<=-16'd9834;
      54002:data<=-16'd10771;
      54003:data<=-16'd9585;
      54004:data<=-16'd9950;
      54005:data<=-16'd9673;
      54006:data<=-16'd8834;
      54007:data<=-16'd9450;
      54008:data<=-16'd8135;
      54009:data<=-16'd9542;
      54010:data<=-16'd11461;
      54011:data<=-16'd8596;
      54012:data<=-16'd13241;
      54013:data<=-16'd24209;
      54014:data<=-16'd26426;
      54015:data<=-16'd23581;
      54016:data<=-16'd22718;
      54017:data<=-16'd21698;
      54018:data<=-16'd20433;
      54019:data<=-16'd20456;
      54020:data<=-16'd20895;
      54021:data<=-16'd20069;
      54022:data<=-16'd19511;
      54023:data<=-16'd19052;
      54024:data<=-16'd16980;
      54025:data<=-16'd16507;
      54026:data<=-16'd15905;
      54027:data<=-16'd13470;
      54028:data<=-16'd14017;
      54029:data<=-16'd12518;
      54030:data<=-16'd6282;
      54031:data<=-16'd3938;
      54032:data<=-16'd4946;
      54033:data<=-16'd5186;
      54034:data<=-16'd4629;
      54035:data<=-16'd3257;
      54036:data<=-16'd3485;
      54037:data<=-16'd3641;
      54038:data<=-16'd2484;
      54039:data<=-16'd2535;
      54040:data<=-16'd2267;
      54041:data<=-16'd2538;
      54042:data<=-16'd1967;
      54043:data<=16'd132;
      54044:data<=-16'd2610;
      54045:data<=-16'd376;
      54046:data<=16'd12413;
      54047:data<=16'd17206;
      54048:data<=16'd14178;
      54049:data<=16'd14882;
      54050:data<=16'd15186;
      54051:data<=16'd14912;
      54052:data<=16'd14815;
      54053:data<=16'd13593;
      54054:data<=16'd14020;
      54055:data<=16'd13421;
      54056:data<=16'd12094;
      54057:data<=16'd11640;
      54058:data<=16'd9828;
      54059:data<=16'd10084;
      54060:data<=16'd10733;
      54061:data<=16'd9323;
      54062:data<=16'd9709;
      54063:data<=16'd9262;
      54064:data<=16'd9081;
      54065:data<=16'd10577;
      54066:data<=16'd9147;
      54067:data<=16'd9348;
      54068:data<=16'd10161;
      54069:data<=16'd7291;
      54070:data<=16'd7157;
      54071:data<=16'd6159;
      54072:data<=16'd949;
      54073:data<=-16'd1624;
      54074:data<=-16'd1779;
      54075:data<=-16'd587;
      54076:data<=-16'd907;
      54077:data<=-16'd2770;
      54078:data<=-16'd981;
      54079:data<=-16'd6211;
      54080:data<=-16'd18638;
      54081:data<=-16'd20923;
      54082:data<=-16'd18883;
      54083:data<=-16'd20078;
      54084:data<=-16'd18606;
      54085:data<=-16'd17344;
      54086:data<=-16'd16498;
      54087:data<=-16'd14630;
      54088:data<=-16'd14621;
      54089:data<=-16'd13944;
      54090:data<=-16'd12731;
      54091:data<=-16'd12000;
      54092:data<=-16'd10928;
      54093:data<=-16'd11050;
      54094:data<=-16'd10464;
      54095:data<=-16'd9979;
      54096:data<=-16'd10766;
      54097:data<=-16'd9538;
      54098:data<=-16'd8798;
      54099:data<=-16'd8992;
      54100:data<=-16'd7829;
      54101:data<=-16'd7479;
      54102:data<=-16'd6352;
      54103:data<=-16'd4981;
      54104:data<=-16'd5532;
      54105:data<=-16'd5272;
      54106:data<=-16'd5335;
      54107:data<=-16'd6347;
      54108:data<=-16'd6748;
      54109:data<=-16'd6437;
      54110:data<=-16'd5065;
      54111:data<=-16'd5659;
      54112:data<=-16'd2209;
      54113:data<=16'd11952;
      54114:data<=16'd22374;
      54115:data<=16'd23099;
      54116:data<=16'd23372;
      54117:data<=16'd22541;
      54118:data<=16'd21405;
      54119:data<=16'd21221;
      54120:data<=16'd18813;
      54121:data<=16'd18190;
      54122:data<=16'd19146;
      54123:data<=16'd17888;
      54124:data<=16'd16853;
      54125:data<=16'd16431;
      54126:data<=16'd16072;
      54127:data<=16'd15350;
      54128:data<=16'd13984;
      54129:data<=16'd13903;
      54130:data<=16'd13726;
      54131:data<=16'd13074;
      54132:data<=16'd12693;
      54133:data<=16'd11168;
      54134:data<=16'd10912;
      54135:data<=16'd11741;
      54136:data<=16'd11179;
      54137:data<=16'd10942;
      54138:data<=16'd10542;
      54139:data<=16'd10272;
      54140:data<=16'd10765;
      54141:data<=16'd10128;
      54142:data<=16'd9959;
      54143:data<=16'd9482;
      54144:data<=16'd8002;
      54145:data<=16'd6558;
      54146:data<=-16'd1063;
      54147:data<=-16'd11524;
      54148:data<=-16'd12979;
      54149:data<=-16'd10093;
      54150:data<=-16'd10422;
      54151:data<=-16'd10551;
      54152:data<=-16'd9492;
      54153:data<=-16'd9395;
      54154:data<=-16'd9009;
      54155:data<=-16'd8737;
      54156:data<=-16'd12718;
      54157:data<=-16'd18177;
      54158:data<=-16'd18553;
      54159:data<=-16'd16642;
      54160:data<=-16'd15676;
      54161:data<=-16'd14692;
      54162:data<=-16'd14460;
      54163:data<=-16'd13608;
      54164:data<=-16'd12122;
      54165:data<=-16'd11438;
      54166:data<=-16'd10601;
      54167:data<=-16'd10229;
      54168:data<=-16'd9417;
      54169:data<=-16'd9222;
      54170:data<=-16'd10968;
      54171:data<=-16'd9820;
      54172:data<=-16'd8633;
      54173:data<=-16'd9999;
      54174:data<=-16'd8745;
      54175:data<=-16'd7993;
      54176:data<=-16'd7342;
      54177:data<=-16'd5932;
      54178:data<=-16'd8751;
      54179:data<=-16'd3667;
      54180:data<=16'd10724;
      54181:data<=16'd14668;
      54182:data<=16'd11917;
      54183:data<=16'd13024;
      54184:data<=16'd13535;
      54185:data<=16'd13626;
      54186:data<=16'd13621;
      54187:data<=16'd12157;
      54188:data<=16'd11406;
      54189:data<=16'd11884;
      54190:data<=16'd12700;
      54191:data<=16'd11811;
      54192:data<=16'd11082;
      54193:data<=16'd11775;
      54194:data<=16'd10857;
      54195:data<=16'd11570;
      54196:data<=16'd12748;
      54197:data<=16'd12082;
      54198:data<=16'd16368;
      54199:data<=16'd20054;
      54200:data<=16'd18269;
      54201:data<=16'd19026;
      54202:data<=16'd19431;
      54203:data<=16'd17590;
      54204:data<=16'd17424;
      54205:data<=16'd16263;
      54206:data<=16'd15838;
      54207:data<=16'd16677;
      54208:data<=16'd17215;
      54209:data<=16'd18351;
      54210:data<=16'd16222;
      54211:data<=16'd15017;
      54212:data<=16'd15529;
      54213:data<=16'd6639;
      54214:data<=-16'd3551;
      54215:data<=-16'd4438;
      54216:data<=-16'd3615;
      54217:data<=-16'd3474;
      54218:data<=-16'd2977;
      54219:data<=-16'd2231;
      54220:data<=16'd36;
      54221:data<=16'd18;
      54222:data<=-16'd1219;
      54223:data<=-16'd297;
      54224:data<=16'd21;
      54225:data<=-16'd378;
      54226:data<=-16'd491;
      54227:data<=-16'd476;
      54228:data<=-16'd513;
      54229:data<=-16'd934;
      54230:data<=-16'd229;
      54231:data<=-16'd115;
      54232:data<=-16'd194;
      54233:data<=16'd2347;
      54234:data<=16'd2751;
      54235:data<=16'd1582;
      54236:data<=16'd2943;
      54237:data<=16'd3298;
      54238:data<=16'd3401;
      54239:data<=16'd2974;
      54240:data<=-16'd1157;
      54241:data<=-16'd4966;
      54242:data<=-16'd6827;
      54243:data<=-16'd6187;
      54244:data<=-16'd4429;
      54245:data<=-16'd5383;
      54246:data<=16'd594;
      54247:data<=16'd13637;
      54248:data<=16'd16876;
      54249:data<=16'd14163;
      54250:data<=16'd15186;
      54251:data<=16'd14522;
      54252:data<=16'd12897;
      54253:data<=16'd13145;
      54254:data<=16'd12693;
      54255:data<=16'd12113;
      54256:data<=16'd11511;
      54257:data<=16'd11050;
      54258:data<=16'd11829;
      54259:data<=16'd12346;
      54260:data<=16'd12152;
      54261:data<=16'd11599;
      54262:data<=16'd10272;
      54263:data<=16'd8919;
      54264:data<=16'd8631;
      54265:data<=16'd9186;
      54266:data<=16'd9235;
      54267:data<=16'd8887;
      54268:data<=16'd8809;
      54269:data<=16'd8918;
      54270:data<=16'd9887;
      54271:data<=16'd10184;
      54272:data<=16'd8889;
      54273:data<=16'd8379;
      54274:data<=16'd7929;
      54275:data<=16'd7545;
      54276:data<=16'd8255;
      54277:data<=16'd7110;
      54278:data<=16'd6361;
      54279:data<=16'd6008;
      54280:data<=-16'd2629;
      54281:data<=-16'd12671;
      54282:data<=-16'd9777;
      54283:data<=-16'd1795;
      54284:data<=-16'd409;
      54285:data<=-16'd1325;
      54286:data<=-16'd845;
      54287:data<=-16'd1118;
      54288:data<=-16'd1225;
      54289:data<=-16'd896;
      54290:data<=-16'd1597;
      54291:data<=-16'd1751;
      54292:data<=-16'd1530;
      54293:data<=-16'd2315;
      54294:data<=-16'd1313;
      54295:data<=16'd922;
      54296:data<=16'd913;
      54297:data<=16'd658;
      54298:data<=16'd1421;
      54299:data<=16'd1403;
      54300:data<=16'd784;
      54301:data<=16'd49;
      54302:data<=-16'd470;
      54303:data<=-16'd754;
      54304:data<=-16'd731;
      54305:data<=-16'd461;
      54306:data<=-16'd1296;
      54307:data<=-16'd509;
      54308:data<=16'd1842;
      54309:data<=16'd111;
      54310:data<=-16'd623;
      54311:data<=16'd1231;
      54312:data<=-16'd1695;
      54313:data<=16'd1701;
      54314:data<=16'd14912;
      54315:data<=16'd18198;
      54316:data<=16'd14145;
      54317:data<=16'd15394;
      54318:data<=16'd15144;
      54319:data<=16'd13220;
      54320:data<=16'd14301;
      54321:data<=16'd13808;
      54322:data<=16'd12932;
      54323:data<=16'd13594;
      54324:data<=16'd10258;
      54325:data<=16'd3607;
      54326:data<=16'd1005;
      54327:data<=16'd2155;
      54328:data<=16'd1710;
      54329:data<=16'd1183;
      54330:data<=16'd1438;
      54331:data<=-16'd27;
      54332:data<=16'd264;
      54333:data<=16'd2370;
      54334:data<=16'd2297;
      54335:data<=16'd1974;
      54336:data<=16'd1562;
      54337:data<=16'd584;
      54338:data<=16'd792;
      54339:data<=16'd705;
      54340:data<=16'd422;
      54341:data<=16'd282;
      54342:data<=-16'd21;
      54343:data<=16'd109;
      54344:data<=-16'd898;
      54345:data<=16'd277;
      54346:data<=16'd1046;
      54347:data<=-16'd8884;
      54348:data<=-16'd18864;
      54349:data<=-16'd17867;
      54350:data<=-16'd16484;
      54351:data<=-16'd16795;
      54352:data<=-16'd14991;
      54353:data<=-16'd14440;
      54354:data<=-16'd13893;
      54355:data<=-16'd13056;
      54356:data<=-16'd13206;
      54357:data<=-16'd12302;
      54358:data<=-16'd10930;
      54359:data<=-16'd10149;
      54360:data<=-16'd9824;
      54361:data<=-16'd9527;
      54362:data<=-16'd9204;
      54363:data<=-16'd8995;
      54364:data<=-16'd8282;
      54365:data<=-16'd8828;
      54366:data<=-16'd6892;
      54367:data<=-16'd96;
      54368:data<=16'd1199;
      54369:data<=-16'd792;
      54370:data<=16'd1733;
      54371:data<=16'd1971;
      54372:data<=16'd1397;
      54373:data<=16'd1989;
      54374:data<=16'd143;
      54375:data<=16'd846;
      54376:data<=16'd784;
      54377:data<=-16'd394;
      54378:data<=16'd1491;
      54379:data<=-16'd1139;
      54380:data<=16'd2367;
      54381:data<=16'd16548;
      54382:data<=16'd19223;
      54383:data<=16'd15341;
      54384:data<=16'd16146;
      54385:data<=16'd13744;
      54386:data<=16'd12157;
      54387:data<=16'd11925;
      54388:data<=16'd10110;
      54389:data<=16'd11174;
      54390:data<=16'd10931;
      54391:data<=16'd9934;
      54392:data<=16'd9958;
      54393:data<=16'd7568;
      54394:data<=16'd7457;
      54395:data<=16'd7206;
      54396:data<=16'd3962;
      54397:data<=16'd3583;
      54398:data<=16'd3491;
      54399:data<=16'd2798;
      54400:data<=16'd2866;
      54401:data<=16'd1706;
      54402:data<=16'd1618;
      54403:data<=16'd1351;
      54404:data<=16'd966;
      54405:data<=16'd1303;
      54406:data<=16'd47;
      54407:data<=16'd678;
      54408:data<=-16'd2256;
      54409:data<=-16'd10534;
      54410:data<=-16'd11862;
      54411:data<=-16'd10860;
      54412:data<=-16'd10974;
      54413:data<=-16'd10384;
      54414:data<=-16'd19684;
      54415:data<=-16'd28241;
      54416:data<=-16'd25535;
      54417:data<=-16'd25175;
      54418:data<=-16'd25431;
      54419:data<=-16'd23135;
      54420:data<=-16'd24529;
      54421:data<=-16'd25241;
      54422:data<=-16'd24650;
      54423:data<=-16'd23908;
      54424:data<=-16'd22632;
      54425:data<=-16'd23108;
      54426:data<=-16'd21705;
      54427:data<=-16'd20013;
      54428:data<=-16'd19910;
      54429:data<=-16'd17499;
      54430:data<=-16'd16492;
      54431:data<=-16'd16938;
      54432:data<=-16'd16868;
      54433:data<=-16'd18064;
      54434:data<=-16'd17461;
      54435:data<=-16'd16824;
      54436:data<=-16'd16630;
      54437:data<=-16'd14656;
      54438:data<=-16'd14662;
      54439:data<=-16'd14222;
      54440:data<=-16'd13869;
      54441:data<=-16'd14654;
      54442:data<=-16'd11626;
      54443:data<=-16'd11450;
      54444:data<=-16'd12087;
      54445:data<=-16'd10143;
      54446:data<=-16'd14642;
      54447:data<=-16'd9673;
      54448:data<=16'd6307;
      54449:data<=16'd7608;
      54450:data<=16'd6904;
      54451:data<=16'd14722;
      54452:data<=16'd15320;
      54453:data<=16'd13914;
      54454:data<=16'd14230;
      54455:data<=16'd12575;
      54456:data<=16'd13133;
      54457:data<=16'd12615;
      54458:data<=16'd11130;
      54459:data<=16'd10241;
      54460:data<=16'd7991;
      54461:data<=16'd8439;
      54462:data<=16'd8727;
      54463:data<=16'd6822;
      54464:data<=16'd6714;
      54465:data<=16'd6407;
      54466:data<=16'd6805;
      54467:data<=16'd6959;
      54468:data<=16'd5210;
      54469:data<=16'd6156;
      54470:data<=16'd6240;
      54471:data<=16'd3823;
      54472:data<=16'd3307;
      54473:data<=16'd3385;
      54474:data<=16'd4411;
      54475:data<=16'd4625;
      54476:data<=16'd3472;
      54477:data<=16'd4276;
      54478:data<=16'd3580;
      54479:data<=16'd3415;
      54480:data<=16'd2155;
      54481:data<=-16'd8272;
      54482:data<=-16'd16354;
      54483:data<=-16'd16719;
      54484:data<=-16'd18054;
      54485:data<=-16'd16759;
      54486:data<=-16'd14792;
      54487:data<=-16'd15647;
      54488:data<=-16'd14005;
      54489:data<=-16'd13544;
      54490:data<=-16'd13439;
      54491:data<=-16'd10677;
      54492:data<=-16'd13382;
      54493:data<=-16'd19296;
      54494:data<=-16'd20168;
      54495:data<=-16'd18639;
      54496:data<=-16'd18698;
      54497:data<=-16'd18804;
      54498:data<=-16'd17061;
      54499:data<=-16'd16572;
      54500:data<=-16'd17017;
      54501:data<=-16'd14666;
      54502:data<=-16'd13024;
      54503:data<=-16'd13112;
      54504:data<=-16'd13035;
      54505:data<=-16'd13179;
      54506:data<=-16'd11632;
      54507:data<=-16'd11797;
      54508:data<=-16'd13624;
      54509:data<=-16'd12019;
      54510:data<=-16'd12105;
      54511:data<=-16'd12252;
      54512:data<=-16'd10245;
      54513:data<=-16'd12436;
      54514:data<=-16'd6775;
      54515:data<=16'd8364;
      54516:data<=16'd11711;
      54517:data<=16'd8161;
      54518:data<=16'd9536;
      54519:data<=16'd9527;
      54520:data<=16'd8896;
      54521:data<=16'd8489;
      54522:data<=16'd6510;
      54523:data<=16'd7063;
      54524:data<=16'd7856;
      54525:data<=16'd7330;
      54526:data<=16'd7912;
      54527:data<=16'd7524;
      54528:data<=16'd7524;
      54529:data<=16'd8059;
      54530:data<=16'd6161;
      54531:data<=16'd6122;
      54532:data<=16'd7530;
      54533:data<=16'd5325;
      54534:data<=16'd6008;
      54535:data<=16'd11902;
      54536:data<=16'd13474;
      54537:data<=16'd11597;
      54538:data<=16'd12090;
      54539:data<=16'd12013;
      54540:data<=16'd11856;
      54541:data<=16'd12613;
      54542:data<=16'd11145;
      54543:data<=16'd10901;
      54544:data<=16'd11667;
      54545:data<=16'd9712;
      54546:data<=16'd9741;
      54547:data<=16'd7410;
      54548:data<=-16'd3597;
      54549:data<=-16'd10901;
      54550:data<=-16'd9542;
      54551:data<=-16'd8787;
      54552:data<=-16'd8936;
      54553:data<=-16'd8053;
      54554:data<=-16'd7847;
      54555:data<=-16'd7253;
      54556:data<=-16'd6408;
      54557:data<=-16'd6011;
      54558:data<=-16'd5996;
      54559:data<=-16'd6799;
      54560:data<=-16'd6886;
      54561:data<=-16'd6253;
      54562:data<=-16'd6605;
      54563:data<=-16'd6373;
      54564:data<=-16'd4983;
      54565:data<=-16'd4672;
      54566:data<=-16'd4921;
      54567:data<=-16'd4282;
      54568:data<=-16'd3720;
      54569:data<=-16'd3388;
      54570:data<=-16'd3636;
      54571:data<=-16'd5037;
      54572:data<=-16'd4470;
      54573:data<=-16'd2908;
      54574:data<=-16'd4173;
      54575:data<=-16'd4103;
      54576:data<=-16'd4502;
      54577:data<=-16'd10578;
      54578:data<=-16'd12678;
      54579:data<=-16'd10793;
      54580:data<=-16'd13106;
      54581:data<=-16'd7090;
      54582:data<=16'd7203;
      54583:data<=16'd10792;
      54584:data<=16'd8716;
      54585:data<=16'd10379;
      54586:data<=16'd10188;
      54587:data<=16'd9656;
      54588:data<=16'd10097;
      54589:data<=16'd8749;
      54590:data<=16'd8382;
      54591:data<=16'd8727;
      54592:data<=16'd8416;
      54593:data<=16'd8337;
      54594:data<=16'd7758;
      54595:data<=16'd8425;
      54596:data<=16'd10332;
      54597:data<=16'd10396;
      54598:data<=16'd9639;
      54599:data<=16'd9397;
      54600:data<=16'd9045;
      54601:data<=16'd8795;
      54602:data<=16'd8549;
      54603:data<=16'd8005;
      54604:data<=16'd7830;
      54605:data<=16'd8395;
      54606:data<=16'd8246;
      54607:data<=16'd7785;
      54608:data<=16'd9068;
      54609:data<=16'd10924;
      54610:data<=16'd12172;
      54611:data<=16'd11477;
      54612:data<=16'd9928;
      54613:data<=16'd11825;
      54614:data<=16'd8771;
      54615:data<=-16'd3798;
      54616:data<=-16'd10246;
      54617:data<=-16'd8763;
      54618:data<=-16'd6940;
      54619:data<=-16'd1105;
      54620:data<=16'd2983;
      54621:data<=16'd2165;
      54622:data<=16'd3715;
      54623:data<=16'd4029;
      54624:data<=16'd2958;
      54625:data<=16'd4255;
      54626:data<=16'd3852;
      54627:data<=16'd3057;
      54628:data<=16'd2773;
      54629:data<=16'd1898;
      54630:data<=16'd3118;
      54631:data<=16'd3712;
      54632:data<=16'd2904;
      54633:data<=16'd3633;
      54634:data<=16'd5048;
      54635:data<=16'd6235;
      54636:data<=16'd5773;
      54637:data<=16'd5210;
      54638:data<=16'd5300;
      54639:data<=16'd4009;
      54640:data<=16'd4899;
      54641:data<=16'd5206;
      54642:data<=16'd2866;
      54643:data<=16'd4014;
      54644:data<=16'd3629;
      54645:data<=16'd2317;
      54646:data<=16'd4040;
      54647:data<=16'd2017;
      54648:data<=16'd7664;
      54649:data<=16'd21937;
      54650:data<=16'd23138;
      54651:data<=16'd19337;
      54652:data<=16'd20521;
      54653:data<=16'd18788;
      54654:data<=16'd18586;
      54655:data<=16'd18810;
      54656:data<=16'd16621;
      54657:data<=16'd16565;
      54658:data<=16'd15973;
      54659:data<=16'd16923;
      54660:data<=16'd15834;
      54661:data<=16'd7808;
      54662:data<=16'd5239;
      54663:data<=16'd6495;
      54664:data<=16'd4106;
      54665:data<=16'd4449;
      54666:data<=16'd4761;
      54667:data<=16'd3900;
      54668:data<=16'd4878;
      54669:data<=16'd3630;
      54670:data<=16'd3307;
      54671:data<=16'd5218;
      54672:data<=16'd5398;
      54673:data<=16'd5171;
      54674:data<=16'd4775;
      54675:data<=16'd4675;
      54676:data<=16'd4528;
      54677:data<=16'd4008;
      54678:data<=16'd4243;
      54679:data<=16'd3472;
      54680:data<=16'd4610;
      54681:data<=16'd2361;
      54682:data<=-16'd10254;
      54683:data<=-16'd16102;
      54684:data<=-16'd12022;
      54685:data<=-16'd12393;
      54686:data<=-16'd11960;
      54687:data<=-16'd10161;
      54688:data<=-16'd10992;
      54689:data<=-16'd9547;
      54690:data<=-16'd9868;
      54691:data<=-16'd10469;
      54692:data<=-16'd8034;
      54693:data<=-16'd8205;
      54694:data<=-16'd8129;
      54695:data<=-16'd7356;
      54696:data<=-16'd7087;
      54697:data<=-16'd4563;
      54698:data<=-16'd4907;
      54699:data<=-16'd6047;
      54700:data<=-16'd5048;
      54701:data<=-16'd6152;
      54702:data<=-16'd3447;
      54703:data<=16'd2344;
      54704:data<=16'd3906;
      54705:data<=16'd3952;
      54706:data<=16'd3444;
      54707:data<=16'd3404;
      54708:data<=16'd3894;
      54709:data<=16'd3366;
      54710:data<=16'd4541;
      54711:data<=16'd4047;
      54712:data<=16'd3092;
      54713:data<=16'd3624;
      54714:data<=16'd79;
      54715:data<=16'd4874;
      54716:data<=16'd19108;
      54717:data<=16'd21455;
      54718:data<=16'd18249;
      54719:data<=16'd19092;
      54720:data<=16'd17188;
      54721:data<=16'd17126;
      54722:data<=16'd18228;
      54723:data<=16'd16389;
      54724:data<=16'd16172;
      54725:data<=16'd15555;
      54726:data<=16'd14433;
      54727:data<=16'd14123;
      54728:data<=16'd12187;
      54729:data<=16'd11333;
      54730:data<=16'd10807;
      54731:data<=16'd9341;
      54732:data<=16'd9567;
      54733:data<=16'd9881;
      54734:data<=16'd10201;
      54735:data<=16'd10110;
      54736:data<=16'd8643;
      54737:data<=16'd8707;
      54738:data<=16'd8478;
      54739:data<=16'd6843;
      54740:data<=16'd6658;
      54741:data<=16'd6534;
      54742:data<=16'd5915;
      54743:data<=16'd6053;
      54744:data<=16'd4643;
      54745:data<=-16'd1008;
      54746:data<=-16'd4707;
      54747:data<=-16'd986;
      54748:data<=-16'd3479;
      54749:data<=-16'd16070;
      54750:data<=-16'd21035;
      54751:data<=-16'd19579;
      54752:data<=-16'd20592;
      54753:data<=-16'd19373;
      54754:data<=-16'd17819;
      54755:data<=-16'd17638;
      54756:data<=-16'd16809;
      54757:data<=-16'd17543;
      54758:data<=-16'd16933;
      54759:data<=-16'd14616;
      54760:data<=-16'd13782;
      54761:data<=-16'd13385;
      54762:data<=-16'd13602;
      54763:data<=-16'd12750;
      54764:data<=-16'd11298;
      54765:data<=-16'd11956;
      54766:data<=-16'd11825;
      54767:data<=-16'd11740;
      54768:data<=-16'd12025;
      54769:data<=-16'd10637;
      54770:data<=-16'd10716;
      54771:data<=-16'd9784;
      54772:data<=-16'd7206;
      54773:data<=-16'd7268;
      54774:data<=-16'd6913;
      54775:data<=-16'd7048;
      54776:data<=-16'd7941;
      54777:data<=-16'd6452;
      54778:data<=-16'd6978;
      54779:data<=-16'd6840;
      54780:data<=-16'd5947;
      54781:data<=-16'd9665;
      54782:data<=-16'd4896;
      54783:data<=16'd8916;
      54784:data<=16'd12513;
      54785:data<=16'd9333;
      54786:data<=16'd11057;
      54787:data<=16'd15264;
      54788:data<=16'd17564;
      54789:data<=16'd16631;
      54790:data<=16'd15362;
      54791:data<=16'd15136;
      54792:data<=16'd14287;
      54793:data<=16'd13712;
      54794:data<=16'd12972;
      54795:data<=16'd12005;
      54796:data<=16'd10824;
      54797:data<=16'd8335;
      54798:data<=16'd7371;
      54799:data<=16'd7580;
      54800:data<=16'd6658;
      54801:data<=16'd6398;
      54802:data<=16'd6053;
      54803:data<=16'd5436;
      54804:data<=16'd5200;
      54805:data<=16'd4049;
      54806:data<=16'd3659;
      54807:data<=16'd3751;
      54808:data<=16'd2867;
      54809:data<=16'd1892;
      54810:data<=16'd781;
      54811:data<=16'd1092;
      54812:data<=16'd1036;
      54813:data<=-16'd146;
      54814:data<=16'd1626;
      54815:data<=-16'd1921;
      54816:data<=-16'd13770;
      54817:data<=-16'd18959;
      54818:data<=-16'd17626;
      54819:data<=-16'd18066;
      54820:data<=-16'd17371;
      54821:data<=-16'd16782;
      54822:data<=-16'd17885;
      54823:data<=-16'd17775;
      54824:data<=-16'd17249;
      54825:data<=-16'd16845;
      54826:data<=-16'd16246;
      54827:data<=-16'd15441;
      54828:data<=-16'd15969;
      54829:data<=-16'd19817;
      54830:data<=-16'd22582;
      54831:data<=-16'd22013;
      54832:data<=-16'd21312;
      54833:data<=-16'd20762;
      54834:data<=-16'd21043;
      54835:data<=-16'd21149;
      54836:data<=-16'd19672;
      54837:data<=-16'd19368;
      54838:data<=-16'd18703;
      54839:data<=-16'd17246;
      54840:data<=-16'd17399;
      54841:data<=-16'd16452;
      54842:data<=-16'd15913;
      54843:data<=-16'd16622;
      54844:data<=-16'd15156;
      54845:data<=-16'd14709;
      54846:data<=-16'd14580;
      54847:data<=-16'd14442;
      54848:data<=-16'd17656;
      54849:data<=-16'd12229;
      54850:data<=16'd2507;
      54851:data<=16'd6760;
      54852:data<=16'd3580;
      54853:data<=16'd4631;
      54854:data<=16'd4608;
      54855:data<=16'd3301;
      54856:data<=16'd3920;
      54857:data<=16'd3952;
      54858:data<=16'd3598;
      54859:data<=16'd2648;
      54860:data<=16'd1192;
      54861:data<=16'd969;
      54862:data<=16'd725;
      54863:data<=16'd464;
      54864:data<=16'd1086;
      54865:data<=16'd1124;
      54866:data<=16'd505;
      54867:data<=16'd367;
      54868:data<=16'd346;
      54869:data<=-16'd35;
      54870:data<=16'd1404;
      54871:data<=16'd5668;
      54872:data<=16'd8325;
      54873:data<=16'd7359;
      54874:data<=16'd6563;
      54875:data<=16'd7389;
      54876:data<=16'd7313;
      54877:data<=16'd6091;
      54878:data<=16'd6323;
      54879:data<=16'd6256;
      54880:data<=16'd5068;
      54881:data<=16'd6778;
      54882:data<=16'd4208;
      54883:data<=-16'd7862;
      54884:data<=-16'd15139;
      54885:data<=-16'd14361;
      54886:data<=-16'd14665;
      54887:data<=-16'd13667;
      54888:data<=-16'd12193;
      54889:data<=-16'd12945;
      54890:data<=-16'd11603;
      54891:data<=-16'd10543;
      54892:data<=-16'd10809;
      54893:data<=-16'd9391;
      54894:data<=-16'd8648;
      54895:data<=-16'd8354;
      54896:data<=-16'd8255;
      54897:data<=-16'd9518;
      54898:data<=-16'd9583;
      54899:data<=-16'd8924;
      54900:data<=-16'd8507;
      54901:data<=-16'd7928;
      54902:data<=-16'd7973;
      54903:data<=-16'd7339;
      54904:data<=-16'd6789;
      54905:data<=-16'd6660;
      54906:data<=-16'd5667;
      54907:data<=-16'd5457;
      54908:data<=-16'd4634;
      54909:data<=-16'd4549;
      54910:data<=-16'd7251;
      54911:data<=-16'd6928;
      54912:data<=-16'd6161;
      54913:data<=-16'd9453;
      54914:data<=-16'd13253;
      54915:data<=-16'd16246;
      54916:data<=-16'd9832;
      54917:data<=16'd4639;
      54918:data<=16'd8070;
      54919:data<=16'd5168;
      54920:data<=16'd6925;
      54921:data<=16'd5802;
      54922:data<=16'd4064;
      54923:data<=16'd4689;
      54924:data<=16'd3424;
      54925:data<=16'd3259;
      54926:data<=16'd3189;
      54927:data<=16'd2437;
      54928:data<=16'd3771;
      54929:data<=16'd3802;
      54930:data<=16'd3315;
      54931:data<=16'd3861;
      54932:data<=16'd2986;
      54933:data<=16'd2858;
      54934:data<=16'd2974;
      54935:data<=16'd1421;
      54936:data<=16'd975;
      54937:data<=16'd1698;
      54938:data<=16'd2064;
      54939:data<=16'd2047;
      54940:data<=16'd1855;
      54941:data<=16'd2221;
      54942:data<=16'd2772;
      54943:data<=16'd2685;
      54944:data<=16'd2816;
      54945:data<=16'd3965;
      54946:data<=16'd3224;
      54947:data<=16'd1171;
      54948:data<=16'd2767;
      54949:data<=-16'd224;
      54950:data<=-16'd12495;
      54951:data<=-16'd18070;
      54952:data<=-16'd15256;
      54953:data<=-16'd15458;
      54954:data<=-16'd14957;
      54955:data<=-16'd10583;
      54956:data<=-16'd5773;
      54957:data<=-16'd2781;
      54958:data<=-16'd3181;
      54959:data<=-16'd3615;
      54960:data<=-16'd3820;
      54961:data<=-16'd4834;
      54962:data<=-16'd3427;
      54963:data<=-16'd2541;
      54964:data<=-16'd3146;
      54965:data<=-16'd2476;
      54966:data<=-16'd2079;
      54967:data<=-16'd1024;
      54968:data<=-16'd878;
      54969:data<=-16'd2065;
      54970:data<=-16'd409;
      54971:data<=-16'd9;
      54972:data<=-16'd1651;
      54973:data<=-16'd1676;
      54974:data<=-16'd1914;
      54975:data<=-16'd852;
      54976:data<=-16'd610;
      54977:data<=-16'd2165;
      54978:data<=-16'd362;
      54979:data<=16'd250;
      54980:data<=-16'd129;
      54981:data<=16'd857;
      54982:data<=-16'd1300;
      54983:data<=16'd4508;
      54984:data<=16'd18049;
      54985:data<=16'd20450;
      54986:data<=16'd17616;
      54987:data<=16'd18313;
      54988:data<=16'd16853;
      54989:data<=16'd16067;
      54990:data<=16'd16786;
      54991:data<=16'd16180;
      54992:data<=16'd15932;
      54993:data<=16'd15320;
      54994:data<=16'd14164;
      54995:data<=16'd13681;
      54996:data<=16'd13946;
      54997:data<=16'd12091;
      54998:data<=16'd6916;
      54999:data<=16'd4825;
      55000:data<=16'd5530;
      55001:data<=16'd4758;
      55002:data<=16'd5198;
      55003:data<=16'd5342;
      55004:data<=16'd4827;
      55005:data<=16'd5705;
      55006:data<=16'd5251;
      55007:data<=16'd4893;
      55008:data<=16'd4871;
      55009:data<=16'd4933;
      55010:data<=16'd6956;
      55011:data<=16'd6699;
      55012:data<=16'd6352;
      55013:data<=16'd7225;
      55014:data<=16'd5526;
      55015:data<=16'd7242;
      55016:data<=16'd4460;
      55017:data<=-16'd9148;
      55018:data<=-16'd14045;
      55019:data<=-16'd11267;
      55020:data<=-16'd12703;
      55021:data<=-16'd11376;
      55022:data<=-16'd9306;
      55023:data<=-16'd9159;
      55024:data<=-16'd7256;
      55025:data<=-16'd6968;
      55026:data<=-16'd6749;
      55027:data<=-16'd5855;
      55028:data<=-16'd5709;
      55029:data<=-16'd4267;
      55030:data<=-16'd4161;
      55031:data<=-16'd4300;
      55032:data<=-16'd3780;
      55033:data<=-16'd4367;
      55034:data<=-16'd2281;
      55035:data<=-16'd796;
      55036:data<=-16'd1111;
      55037:data<=16'd325;
      55038:data<=-16'd594;
      55039:data<=16'd1498;
      55040:data<=16'd8153;
      55041:data<=16'd9262;
      55042:data<=16'd8937;
      55043:data<=16'd9180;
      55044:data<=16'd7109;
      55045:data<=16'd7086;
      55046:data<=16'd7071;
      55047:data<=16'd8308;
      55048:data<=16'd9767;
      55049:data<=16'd7118;
      55050:data<=16'd13735;
      55051:data<=16'd26373;
      55052:data<=16'd26823;
      55053:data<=16'd23962;
      55054:data<=16'd24647;
      55055:data<=16'd23344;
      55056:data<=16'd22903;
      55057:data<=16'd21961;
      55058:data<=16'd19936;
      55059:data<=16'd20363;
      55060:data<=16'd20566;
      55061:data<=16'd20024;
      55062:data<=16'd19839;
      55063:data<=16'd19035;
      55064:data<=16'd17872;
      55065:data<=16'd17035;
      55066:data<=16'd16921;
      55067:data<=16'd15763;
      55068:data<=16'd14292;
      55069:data<=16'd14070;
      55070:data<=16'd12800;
      55071:data<=16'd12609;
      55072:data<=16'd13631;
      55073:data<=16'd12740;
      55074:data<=16'd12928;
      55075:data<=16'd12953;
      55076:data<=16'd11847;
      55077:data<=16'd12257;
      55078:data<=16'd10933;
      55079:data<=16'd10507;
      55080:data<=16'd11477;
      55081:data<=16'd7661;
      55082:data<=16'd3570;
      55083:data<=-16'd2820;
      55084:data<=-16'd14457;
      55085:data<=-16'd17829;
      55086:data<=-16'd14468;
      55087:data<=-16'd14557;
      55088:data<=-16'd13928;
      55089:data<=-16'd13259;
      55090:data<=-16'd14095;
      55091:data<=-16'd12792;
      55092:data<=-16'd12199;
      55093:data<=-16'd12521;
      55094:data<=-16'd11320;
      55095:data<=-16'd10754;
      55096:data<=-16'd10746;
      55097:data<=-16'd9538;
      55098:data<=-16'd8066;
      55099:data<=-16'd7843;
      55100:data<=-16'd7682;
      55101:data<=-16'd6807;
      55102:data<=-16'd7069;
      55103:data<=-16'd7227;
      55104:data<=-16'd6598;
      55105:data<=-16'd6763;
      55106:data<=-16'd6232;
      55107:data<=-16'd6137;
      55108:data<=-16'd6919;
      55109:data<=-16'd5607;
      55110:data<=-16'd4590;
      55111:data<=-16'd4281;
      55112:data<=-16'd3156;
      55113:data<=-16'd3501;
      55114:data<=-16'd3037;
      55115:data<=-16'd2707;
      55116:data<=-16'd3782;
      55117:data<=16'd3460;
      55118:data<=16'd14838;
      55119:data<=16'd16230;
      55120:data<=16'd13820;
      55121:data<=16'd13890;
      55122:data<=16'd12698;
      55123:data<=16'd15593;
      55124:data<=16'd21892;
      55125:data<=16'd22016;
      55126:data<=16'd19752;
      55127:data<=16'd19647;
      55128:data<=16'd17957;
      55129:data<=16'd16575;
      55130:data<=16'd16087;
      55131:data<=16'd14413;
      55132:data<=16'd14392;
      55133:data<=16'd14266;
      55134:data<=16'd13085;
      55135:data<=16'd14383;
      55136:data<=16'd14255;
      55137:data<=16'd12586;
      55138:data<=16'd13518;
      55139:data<=16'd12693;
      55140:data<=16'd10572;
      55141:data<=16'd10458;
      55142:data<=16'd9550;
      55143:data<=16'd9215;
      55144:data<=16'd9133;
      55145:data<=16'd7602;
      55146:data<=16'd8029;
      55147:data<=16'd8017;
      55148:data<=16'd7850;
      55149:data<=16'd10373;
      55150:data<=16'd5168;
      55151:data<=-16'd7659;
      55152:data<=-16'd12455;
      55153:data<=-16'd10786;
      55154:data<=-16'd11368;
      55155:data<=-16'd11226;
      55156:data<=-16'd10457;
      55157:data<=-16'd11411;
      55158:data<=-16'd10555;
      55159:data<=-16'd8927;
      55160:data<=-16'd9019;
      55161:data<=-16'd7853;
      55162:data<=-16'd7107;
      55163:data<=-16'd7893;
      55164:data<=-16'd6294;
      55165:data<=-16'd7679;
      55166:data<=-16'd14145;
      55167:data<=-16'd15864;
      55168:data<=-16'd14119;
      55169:data<=-16'd14481;
      55170:data<=-16'd14013;
      55171:data<=-16'd13568;
      55172:data<=-16'd12924;
      55173:data<=-16'd10557;
      55174:data<=-16'd10351;
      55175:data<=-16'd10608;
      55176:data<=-16'd9646;
      55177:data<=-16'd10169;
      55178:data<=-16'd9771;
      55179:data<=-16'd9335;
      55180:data<=-16'd10542;
      55181:data<=-16'd9608;
      55182:data<=-16'd9315;
      55183:data<=-16'd9379;
      55184:data<=-16'd1545;
      55185:data<=16'd8651;
      55186:data<=16'd10323;
      55187:data<=16'd7799;
      55188:data<=16'd7526;
      55189:data<=16'd7542;
      55190:data<=16'd7245;
      55191:data<=16'd7392;
      55192:data<=16'd6187;
      55193:data<=16'd4918;
      55194:data<=16'd4843;
      55195:data<=16'd4240;
      55196:data<=16'd4279;
      55197:data<=16'd3777;
      55198:data<=16'd1228;
      55199:data<=16'd1036;
      55200:data<=16'd1568;
      55201:data<=16'd315;
      55202:data<=16'd942;
      55203:data<=16'd804;
      55204:data<=-16'd79;
      55205:data<=16'd987;
      55206:data<=-16'd632;
      55207:data<=16'd429;
      55208:data<=16'd7189;
      55209:data<=16'd7996;
      55210:data<=16'd5172;
      55211:data<=16'd4808;
      55212:data<=16'd3410;
      55213:data<=16'd3912;
      55214:data<=16'd4055;
      55215:data<=16'd2452;
      55216:data<=16'd4831;
      55217:data<=16'd309;
      55218:data<=-16'd12783;
      55219:data<=-16'd16452;
      55220:data<=-16'd13670;
      55221:data<=-16'd13905;
      55222:data<=-16'd13873;
      55223:data<=-16'd14936;
      55224:data<=-16'd16134;
      55225:data<=-16'd14366;
      55226:data<=-16'd13461;
      55227:data<=-16'd13761;
      55228:data<=-16'd13341;
      55229:data<=-16'd12754;
      55230:data<=-16'd12339;
      55231:data<=-16'd12219;
      55232:data<=-16'd11417;
      55233:data<=-16'd10745;
      55234:data<=-16'd11254;
      55235:data<=-16'd11755;
      55236:data<=-16'd12363;
      55237:data<=-16'd12251;
      55238:data<=-16'd11556;
      55239:data<=-16'd11367;
      55240:data<=-16'd10266;
      55241:data<=-16'd10085;
      55242:data<=-16'd10449;
      55243:data<=-16'd8980;
      55244:data<=-16'd9232;
      55245:data<=-16'd9683;
      55246:data<=-16'd8997;
      55247:data<=-16'd10061;
      55248:data<=-16'd9326;
      55249:data<=-16'd11223;
      55250:data<=-16'd16374;
      55251:data<=-16'd9900;
      55252:data<=16'd819;
      55253:data<=16'd1127;
      55254:data<=-16'd32;
      55255:data<=16'd799;
      55256:data<=16'd194;
      55257:data<=16'd879;
      55258:data<=16'd916;
      55259:data<=-16'd82;
      55260:data<=-16'd717;
      55261:data<=-16'd2009;
      55262:data<=-16'd2105;
      55263:data<=-16'd1700;
      55264:data<=-16'd2206;
      55265:data<=-16'd2332;
      55266:data<=-16'd2094;
      55267:data<=-16'd1553;
      55268:data<=-16'd1760;
      55269:data<=-16'd2290;
      55270:data<=-16'd1811;
      55271:data<=-16'd1811;
      55272:data<=-16'd1844;
      55273:data<=-16'd2710;
      55274:data<=-16'd4303;
      55275:data<=-16'd3450;
      55276:data<=-16'd3215;
      55277:data<=-16'd3577;
      55278:data<=-16'd2496;
      55279:data<=-16'd3148;
      55280:data<=-16'd2261;
      55281:data<=-16'd1554;
      55282:data<=-16'd3278;
      55283:data<=-16'd365;
      55284:data<=-16'd4217;
      55285:data<=-16'd18845;
      55286:data<=-16'd23214;
      55287:data<=-16'd20227;
      55288:data<=-16'd20415;
      55289:data<=-16'd18859;
      55290:data<=-16'd19170;
      55291:data<=-16'd18104;
      55292:data<=-16'd10543;
      55293:data<=-16'd6807;
      55294:data<=-16'd7442;
      55295:data<=-16'd6987;
      55296:data<=-16'd6508;
      55297:data<=-16'd6115;
      55298:data<=-16'd7100;
      55299:data<=-16'd7579;
      55300:data<=-16'd6241;
      55301:data<=-16'd6199;
      55302:data<=-16'd5729;
      55303:data<=-16'd4664;
      55304:data<=-16'd4479;
      55305:data<=-16'd3695;
      55306:data<=-16'd3253;
      55307:data<=-16'd2875;
      55308:data<=-16'd2663;
      55309:data<=-16'd2983;
      55310:data<=-16'd2500;
      55311:data<=-16'd3660;
      55312:data<=-16'd4608;
      55313:data<=-16'd3395;
      55314:data<=-16'd3667;
      55315:data<=-16'd3228;
      55316:data<=-16'd3321;
      55317:data<=-16'd2708;
      55318:data<=16'd7571;
      55319:data<=16'd16888;
      55320:data<=16'd15887;
      55321:data<=16'd15255;
      55322:data<=16'd15051;
      55323:data<=16'd12455;
      55324:data<=16'd11761;
      55325:data<=16'd11250;
      55326:data<=16'd11024;
      55327:data<=16'd11056;
      55328:data<=16'd10241;
      55329:data<=16'd10840;
      55330:data<=16'd10313;
      55331:data<=16'd9409;
      55332:data<=16'd10698;
      55333:data<=16'd8657;
      55334:data<=16'd3380;
      55335:data<=-16'd99;
      55336:data<=-16'd1556;
      55337:data<=-16'd1927;
      55338:data<=-16'd2014;
      55339:data<=-16'd1438;
      55340:data<=-16'd773;
      55341:data<=-16'd787;
      55342:data<=-16'd397;
      55343:data<=-16'd684;
      55344:data<=-16'd540;
      55345:data<=16'd311;
      55346:data<=-16'd346;
      55347:data<=16'd135;
      55348:data<=-16'd805;
      55349:data<=-16'd3018;
      55350:data<=-16'd20;
      55351:data<=-16'd3603;
      55352:data<=-16'd16909;
      55353:data<=-16'd20498;
      55354:data<=-16'd16821;
      55355:data<=-16'd16800;
      55356:data<=-16'd15755;
      55357:data<=-16'd15038;
      55358:data<=-16'd15459;
      55359:data<=-16'd13302;
      55360:data<=-16'd12863;
      55361:data<=-16'd14424;
      55362:data<=-16'd13944;
      55363:data<=-16'd12910;
      55364:data<=-16'd12322;
      55365:data<=-16'd11397;
      55366:data<=-16'd10754;
      55367:data<=-16'd10596;
      55368:data<=-16'd9859;
      55369:data<=-16'd8583;
      55370:data<=-16'd7921;
      55371:data<=-16'd7418;
      55372:data<=-16'd6733;
      55373:data<=-16'd6981;
      55374:data<=-16'd7938;
      55375:data<=-16'd6087;
      55376:data<=-16'd211;
      55377:data<=16'd3021;
      55378:data<=16'd2199;
      55379:data<=16'd2981;
      55380:data<=16'd2907;
      55381:data<=16'd2215;
      55382:data<=16'd4088;
      55383:data<=16'd2870;
      55384:data<=16'd3903;
      55385:data<=16'd14324;
      55386:data<=16'd21561;
      55387:data<=16'd20973;
      55388:data<=16'd20557;
      55389:data<=16'd20418;
      55390:data<=16'd19552;
      55391:data<=16'd18850;
      55392:data<=16'd18390;
      55393:data<=16'd18351;
      55394:data<=16'd17452;
      55395:data<=16'd16660;
      55396:data<=16'd16358;
      55397:data<=16'd15506;
      55398:data<=16'd15793;
      55399:data<=16'd16486;
      55400:data<=16'd16322;
      55401:data<=16'd15985;
      55402:data<=16'd15057;
      55403:data<=16'd14439;
      55404:data<=16'd13973;
      55405:data<=16'd13435;
      55406:data<=16'd13870;
      55407:data<=16'd13204;
      55408:data<=16'd11958;
      55409:data<=16'd11690;
      55410:data<=16'd11767;
      55411:data<=16'd13631;
      55412:data<=16'd13957;
      55413:data<=16'd11855;
      55414:data<=16'd12287;
      55415:data<=16'd11600;
      55416:data<=16'd10968;
      55417:data<=16'd12372;
      55418:data<=16'd2441;
      55419:data<=-16'd13740;
      55420:data<=-16'd17194;
      55421:data<=-16'd14697;
      55422:data<=-16'd15270;
      55423:data<=-16'd13725;
      55424:data<=-16'd11546;
      55425:data<=-16'd11180;
      55426:data<=-16'd9979;
      55427:data<=-16'd8972;
      55428:data<=-16'd9444;
      55429:data<=-16'd9474;
      55430:data<=-16'd8575;
      55431:data<=-16'd7970;
      55432:data<=-16'd7504;
      55433:data<=-16'd7468;
      55434:data<=-16'd7689;
      55435:data<=-16'd5480;
      55436:data<=-16'd2168;
      55437:data<=-16'd1221;
      55438:data<=-16'd1351;
      55439:data<=-16'd1143;
      55440:data<=-16'd681;
      55441:data<=-16'd431;
      55442:data<=-16'd687;
      55443:data<=-16'd55;
      55444:data<=16'd326;
      55445:data<=16'd103;
      55446:data<=16'd588;
      55447:data<=-16'd475;
      55448:data<=-16'd99;
      55449:data<=16'd2870;
      55450:data<=16'd1710;
      55451:data<=16'd3378;
      55452:data<=16'd13820;
      55453:data<=16'd20236;
      55454:data<=16'd19726;
      55455:data<=16'd19337;
      55456:data<=16'd19099;
      55457:data<=16'd19049;
      55458:data<=16'd17725;
      55459:data<=16'd16607;
      55460:data<=16'd20644;
      55461:data<=16'd24209;
      55462:data<=16'd23450;
      55463:data<=16'd22703;
      55464:data<=16'd21649;
      55465:data<=16'd20289;
      55466:data<=16'd19708;
      55467:data<=16'd18906;
      55468:data<=16'd18624;
      55469:data<=16'd17866;
      55470:data<=16'd16539;
      55471:data<=16'd15923;
      55472:data<=16'd14963;
      55473:data<=16'd15283;
      55474:data<=16'd16345;
      55475:data<=16'd15414;
      55476:data<=16'd14624;
      55477:data<=16'd14038;
      55478:data<=16'd13247;
      55479:data<=16'd13086;
      55480:data<=16'd12049;
      55481:data<=16'd11773;
      55482:data<=16'd11248;
      55483:data<=16'd10179;
      55484:data<=16'd12151;
      55485:data<=16'd7394;
      55486:data<=-16'd5103;
      55487:data<=-16'd8061;
      55488:data<=-16'd5444;
      55489:data<=-16'd7109;
      55490:data<=-16'd6922;
      55491:data<=-16'd6437;
      55492:data<=-16'd7171;
      55493:data<=-16'd5799;
      55494:data<=-16'd5692;
      55495:data<=-16'd5797;
      55496:data<=-16'd5230;
      55497:data<=-16'd6090;
      55498:data<=-16'd5298;
      55499:data<=-16'd3936;
      55500:data<=-16'd3721;
      55501:data<=-16'd4120;
      55502:data<=-16'd7426;
      55503:data<=-16'd9821;
      55504:data<=-16'd8931;
      55505:data<=-16'd9180;
      55506:data<=-16'd9636;
      55507:data<=-16'd8960;
      55508:data<=-16'd8507;
      55509:data<=-16'd8014;
      55510:data<=-16'd7743;
      55511:data<=-16'd6819;
      55512:data<=-16'd5585;
      55513:data<=-16'd5799;
      55514:data<=-16'd6125;
      55515:data<=-16'd5312;
      55516:data<=-16'd4992;
      55517:data<=-16'd6757;
      55518:data<=-16'd4397;
      55519:data<=16'd6484;
      55520:data<=16'd13860;
      55521:data<=16'd12483;
      55522:data<=16'd11603;
      55523:data<=16'd12361;
      55524:data<=16'd13124;
      55525:data<=16'd13396;
      55526:data<=16'd11676;
      55527:data<=16'd11623;
      55528:data<=16'd11508;
      55529:data<=16'd9580;
      55530:data<=16'd9943;
      55531:data<=16'd9357;
      55532:data<=16'd7906;
      55533:data<=16'd8332;
      55534:data<=16'd7219;
      55535:data<=16'd7450;
      55536:data<=16'd8881;
      55537:data<=16'd7562;
      55538:data<=16'd7272;
      55539:data<=16'd7090;
      55540:data<=16'd6208;
      55541:data<=16'd6883;
      55542:data<=16'd5809;
      55543:data<=16'd5442;
      55544:data<=16'd8660;
      55545:data<=16'd11398;
      55546:data<=16'd11462;
      55547:data<=16'd9370;
      55548:data<=16'd9556;
      55549:data<=16'd10731;
      55550:data<=16'd9529;
      55551:data<=16'd11033;
      55552:data<=16'd6801;
      55553:data<=-16'd6931;
      55554:data<=-16'd11071;
      55555:data<=-16'd7956;
      55556:data<=-16'd9576;
      55557:data<=-16'd9300;
      55558:data<=-16'd8505;
      55559:data<=-16'd9800;
      55560:data<=-16'd8617;
      55561:data<=-16'd7347;
      55562:data<=-16'd6543;
      55563:data<=-16'd6273;
      55564:data<=-16'd7074;
      55565:data<=-16'd6216;
      55566:data<=-16'd6181;
      55567:data<=-16'd7051;
      55568:data<=-16'd6495;
      55569:data<=-16'd6481;
      55570:data<=-16'd5988;
      55571:data<=-16'd5607;
      55572:data<=-16'd6369;
      55573:data<=-16'd5476;
      55574:data<=-16'd4264;
      55575:data<=-16'd3583;
      55576:data<=-16'd2914;
      55577:data<=-16'd3635;
      55578:data<=-16'd4235;
      55579:data<=-16'd4035;
      55580:data<=-16'd3990;
      55581:data<=-16'd4285;
      55582:data<=-16'd4435;
      55583:data<=-16'd4232;
      55584:data<=-16'd5251;
      55585:data<=-16'd2457;
      55586:data<=16'd5568;
      55587:data<=16'd7809;
      55588:data<=16'd5927;
      55589:data<=16'd6587;
      55590:data<=16'd5850;
      55591:data<=16'd5715;
      55592:data<=16'd6115;
      55593:data<=16'd4625;
      55594:data<=16'd4978;
      55595:data<=16'd3905;
      55596:data<=16'd2340;
      55597:data<=16'd3709;
      55598:data<=16'd1932;
      55599:data<=-16'd112;
      55600:data<=16'd388;
      55601:data<=-16'd573;
      55602:data<=-16'd508;
      55603:data<=-16'd911;
      55604:data<=-16'd1912;
      55605:data<=-16'd837;
      55606:data<=-16'd1750;
      55607:data<=-16'd2000;
      55608:data<=-16'd652;
      55609:data<=-16'd1500;
      55610:data<=-16'd1434;
      55611:data<=-16'd2551;
      55612:data<=-16'd4349;
      55613:data<=-16'd3283;
      55614:data<=-16'd4076;
      55615:data<=-16'd4300;
      55616:data<=-16'd3915;
      55617:data<=-16'd5265;
      55618:data<=-16'd2563;
      55619:data<=-16'd6434;
      55620:data<=-16'd19969;
      55621:data<=-16'd23237;
      55622:data<=-16'd19418;
      55623:data<=-16'd20606;
      55624:data<=-16'd21667;
      55625:data<=-16'd21171;
      55626:data<=-16'd20961;
      55627:data<=-16'd20375;
      55628:data<=-16'd17350;
      55629:data<=-16'd12146;
      55630:data<=-16'd11151;
      55631:data<=-16'd12117;
      55632:data<=-16'd10827;
      55633:data<=-16'd10947;
      55634:data<=-16'd10517;
      55635:data<=-16'd9370;
      55636:data<=-16'd10389;
      55637:data<=-16'd10699;
      55638:data<=-16'd10593;
      55639:data<=-16'd10545;
      55640:data<=-16'd9586;
      55641:data<=-16'd9177;
      55642:data<=-16'd8731;
      55643:data<=-16'd8722;
      55644:data<=-16'd9021;
      55645:data<=-16'd8957;
      55646:data<=-16'd9091;
      55647:data<=-16'd7462;
      55648:data<=-16'd7509;
      55649:data<=-16'd9937;
      55650:data<=-16'd9586;
      55651:data<=-16'd10423;
      55652:data<=-16'd7699;
      55653:data<=16'd4340;
      55654:data<=16'd10548;
      55655:data<=16'd8804;
      55656:data<=16'd9138;
      55657:data<=16'd8874;
      55658:data<=16'd8229;
      55659:data<=16'd8408;
      55660:data<=16'd8014;
      55661:data<=16'd7779;
      55662:data<=16'd5403;
      55663:data<=16'd4308;
      55664:data<=16'd5254;
      55665:data<=16'd3603;
      55666:data<=16'd3767;
      55667:data<=16'd4087;
      55668:data<=16'd2696;
      55669:data<=16'd4561;
      55670:data<=16'd2071;
      55671:data<=-16'd3858;
      55672:data<=-16'd3374;
      55673:data<=-16'd3253;
      55674:data<=-16'd5474;
      55675:data<=-16'd5377;
      55676:data<=-16'd5247;
      55677:data<=-16'd4723;
      55678:data<=-16'd4525;
      55679:data<=-16'd4376;
      55680:data<=-16'd3412;
      55681:data<=-16'd4407;
      55682:data<=-16'd4012;
      55683:data<=-16'd3683;
      55684:data<=-16'd4863;
      55685:data<=-16'd1565;
      55686:data<=-16'd5934;
      55687:data<=-16'd21070;
      55688:data<=-16'd24950;
      55689:data<=-16'd20591;
      55690:data<=-16'd21181;
      55691:data<=-16'd20483;
      55692:data<=-16'd19167;
      55693:data<=-16'd19599;
      55694:data<=-16'd17925;
      55695:data<=-16'd17127;
      55696:data<=-16'd16982;
      55697:data<=-16'd15361;
      55698:data<=-16'd15282;
      55699:data<=-16'd16022;
      55700:data<=-16'd15784;
      55701:data<=-16'd15273;
      55702:data<=-16'd14377;
      55703:data<=-16'd13085;
      55704:data<=-16'd11969;
      55705:data<=-16'd11844;
      55706:data<=-16'd11685;
      55707:data<=-16'd10352;
      55708:data<=-16'd9597;
      55709:data<=-16'd9125;
      55710:data<=-16'd8580;
      55711:data<=-16'd9966;
      55712:data<=-16'd9562;
      55713:data<=-16'd4331;
      55714:data<=-16'd1504;
      55715:data<=-16'd3680;
      55716:data<=-16'd3363;
      55717:data<=-16'd1736;
      55718:data<=-16'd3601;
      55719:data<=16'd26;
      55720:data<=16'd11690;
      55721:data<=16'd17646;
      55722:data<=16'd16321;
      55723:data<=16'd15846;
      55724:data<=16'd14589;
      55725:data<=16'd12501;
      55726:data<=16'd12724;
      55727:data<=16'd12686;
      55728:data<=16'd11728;
      55729:data<=16'd11248;
      55730:data<=16'd10592;
      55731:data<=16'd10270;
      55732:data<=16'd10214;
      55733:data<=16'd9558;
      55734:data<=16'd8947;
      55735:data<=16'd8845;
      55736:data<=16'd8434;
      55737:data<=16'd6986;
      55738:data<=16'd5917;
      55739:data<=16'd5937;
      55740:data<=16'd5621;
      55741:data<=16'd5480;
      55742:data<=16'd5683;
      55743:data<=16'd5582;
      55744:data<=16'd5755;
      55745:data<=16'd5081;
      55746:data<=16'd4604;
      55747:data<=16'd5523;
      55748:data<=16'd4613;
      55749:data<=16'd3005;
      55750:data<=16'd2046;
      55751:data<=16'd1239;
      55752:data<=16'd3513;
      55753:data<=-16'd80;
      55754:data<=-16'd15145;
      55755:data<=-16'd23179;
      55756:data<=-16'd19839;
      55757:data<=-16'd19202;
      55758:data<=-16'd19713;
      55759:data<=-16'd18116;
      55760:data<=-16'd17396;
      55761:data<=-16'd16343;
      55762:data<=-16'd16688;
      55763:data<=-16'd17438;
      55764:data<=-16'd15726;
      55765:data<=-16'd15229;
      55766:data<=-16'd15164;
      55767:data<=-16'd13555;
      55768:data<=-16'd12919;
      55769:data<=-16'd12079;
      55770:data<=-16'd11044;
      55771:data<=-16'd10854;
      55772:data<=-16'd9448;
      55773:data<=-16'd8517;
      55774:data<=-16'd9227;
      55775:data<=-16'd9233;
      55776:data<=-16'd8883;
      55777:data<=-16'd8457;
      55778:data<=-16'd8050;
      55779:data<=-16'd8452;
      55780:data<=-16'd7339;
      55781:data<=-16'd5488;
      55782:data<=-16'd6243;
      55783:data<=-16'd5905;
      55784:data<=-16'd4162;
      55785:data<=-16'd5773;
      55786:data<=-16'd2325;
      55787:data<=16'd10334;
      55788:data<=16'd16436;
      55789:data<=16'd13581;
      55790:data<=16'd13820;
      55791:data<=16'd14715;
      55792:data<=16'd13157;
      55793:data<=16'd13508;
      55794:data<=16'd13314;
      55795:data<=16'd12031;
      55796:data<=16'd14126;
      55797:data<=16'd17593;
      55798:data<=16'd18333;
      55799:data<=16'd18052;
      55800:data<=16'd18930;
      55801:data<=16'd18747;
      55802:data<=16'd17681;
      55803:data<=16'd17823;
      55804:data<=16'd17321;
      55805:data<=16'd16669;
      55806:data<=16'd16556;
      55807:data<=16'd15262;
      55808:data<=16'd15188;
      55809:data<=16'd15396;
      55810:data<=16'd13958;
      55811:data<=16'd14628;
      55812:data<=16'd15829;
      55813:data<=16'd15285;
      55814:data<=16'd14454;
      55815:data<=16'd13450;
      55816:data<=16'd14107;
      55817:data<=16'd13564;
      55818:data<=16'd11906;
      55819:data<=16'd14023;
      55820:data<=16'd9097;
      55821:data<=-16'd3633;
      55822:data<=-16'd6689;
      55823:data<=-16'd4269;
      55824:data<=-16'd4672;
      55825:data<=-16'd3128;
      55826:data<=-16'd2811;
      55827:data<=-16'd3400;
      55828:data<=-16'd1606;
      55829:data<=-16'd1923;
      55830:data<=-16'd2458;
      55831:data<=-16'd1168;
      55832:data<=-16'd1454;
      55833:data<=-16'd1738;
      55834:data<=-16'd896;
      55835:data<=-16'd943;
      55836:data<=-16'd673;
      55837:data<=16'd1427;
      55838:data<=16'd1075;
      55839:data<=-16'd3247;
      55840:data<=-16'd4496;
      55841:data<=-16'd2919;
      55842:data<=-16'd3230;
      55843:data<=-16'd3031;
      55844:data<=-16'd3081;
      55845:data<=-16'd3683;
      55846:data<=-16'd2746;
      55847:data<=-16'd2755;
      55848:data<=-16'd2529;
      55849:data<=-16'd1651;
      55850:data<=-16'd905;
      55851:data<=16'd678;
      55852:data<=-16'd729;
      55853:data<=16'd2499;
      55854:data<=16'd14868;
      55855:data<=16'd19170;
      55856:data<=16'd16366;
      55857:data<=16'd17526;
      55858:data<=16'd16785;
      55859:data<=16'd15664;
      55860:data<=16'd15949;
      55861:data<=16'd14744;
      55862:data<=16'd16222;
      55863:data<=16'd16448;
      55864:data<=16'd14266;
      55865:data<=16'd14719;
      55866:data<=16'd14085;
      55867:data<=16'd13197;
      55868:data<=16'd13285;
      55869:data<=16'd12064;
      55870:data<=16'd12052;
      55871:data<=16'd11523;
      55872:data<=16'd10411;
      55873:data<=16'd10075;
      55874:data<=16'd9194;
      55875:data<=16'd11091;
      55876:data<=16'd11972;
      55877:data<=16'd10357;
      55878:data<=16'd11461;
      55879:data<=16'd10037;
      55880:data<=16'd10176;
      55881:data<=16'd15646;
      55882:data<=16'd15509;
      55883:data<=16'd14093;
      55884:data<=16'd14210;
      55885:data<=16'd12167;
      55886:data<=16'd14178;
      55887:data<=16'd10131;
      55888:data<=-16'd2138;
      55889:data<=-16'd4661;
      55890:data<=-16'd2811;
      55891:data<=-16'd4035;
      55892:data<=-16'd3638;
      55893:data<=-16'd4376;
      55894:data<=-16'd4178;
      55895:data<=-16'd2787;
      55896:data<=-16'd3242;
      55897:data<=-16'd2438;
      55898:data<=-16'd2670;
      55899:data<=-16'd2939;
      55900:data<=-16'd751;
      55901:data<=-16'd611;
      55902:data<=-16'd640;
      55903:data<=-16'd265;
      55904:data<=-16'd1189;
      55905:data<=-16'd464;
      55906:data<=-16'd115;
      55907:data<=-16'd517;
      55908:data<=-16'd347;
      55909:data<=-16'd1133;
      55910:data<=-16'd1113;
      55911:data<=-16'd951;
      55912:data<=-16'd405;
      55913:data<=16'd1001;
      55914:data<=16'd185;
      55915:data<=16'd281;
      55916:data<=16'd558;
      55917:data<=-16'd408;
      55918:data<=16'd910;
      55919:data<=-16'd936;
      55920:data<=16'd1485;
      55921:data<=16'd15138;
      55922:data<=16'd18023;
      55923:data<=16'd10134;
      55924:data<=16'd10428;
      55925:data<=16'd12037;
      55926:data<=16'd10810;
      55927:data<=16'd10991;
      55928:data<=16'd10090;
      55929:data<=16'd9765;
      55930:data<=16'd9157;
      55931:data<=16'd7741;
      55932:data<=16'd7767;
      55933:data<=16'd6705;
      55934:data<=16'd6135;
      55935:data<=16'd6267;
      55936:data<=16'd5215;
      55937:data<=16'd6159;
      55938:data<=16'd6862;
      55939:data<=16'd5820;
      55940:data<=16'd5614;
      55941:data<=16'd5127;
      55942:data<=16'd5324;
      55943:data<=16'd5372;
      55944:data<=16'd4202;
      55945:data<=16'd4572;
      55946:data<=16'd4396;
      55947:data<=16'd3368;
      55948:data<=16'd3207;
      55949:data<=16'd3253;
      55950:data<=16'd4739;
      55951:data<=16'd4259;
      55952:data<=16'd2955;
      55953:data<=16'd4567;
      55954:data<=-16'd1571;
      55955:data<=-16'd13359;
      55956:data<=-16'd15561;
      55957:data<=-16'd13253;
      55958:data<=-16'd13385;
      55959:data<=-16'd13117;
      55960:data<=-16'd13546;
      55961:data<=-16'd13118;
      55962:data<=-16'd11244;
      55963:data<=-16'd10745;
      55964:data<=-16'd8449;
      55965:data<=-16'd3736;
      55966:data<=-16'd2003;
      55967:data<=-16'd3192;
      55968:data<=-16'd2964;
      55969:data<=-16'd2055;
      55970:data<=-16'd2505;
      55971:data<=-16'd2390;
      55972:data<=-16'd2215;
      55973:data<=-16'd2892;
      55974:data<=-16'd2300;
      55975:data<=-16'd1193;
      55976:data<=-16'd526;
      55977:data<=-16'd682;
      55978:data<=-16'd1632;
      55979:data<=-16'd999;
      55980:data<=-16'd983;
      55981:data<=-16'd1680;
      55982:data<=-16'd346;
      55983:data<=-16'd1427;
      55984:data<=-16'd2432;
      55985:data<=-16'd732;
      55986:data<=-16'd2807;
      55987:data<=16'd150;
      55988:data<=16'd12301;
      55989:data<=16'd16795;
      55990:data<=16'd13907;
      55991:data<=16'd13832;
      55992:data<=16'd13471;
      55993:data<=16'd12390;
      55994:data<=16'd12160;
      55995:data<=16'd11160;
      55996:data<=16'd10298;
      55997:data<=16'd9723;
      55998:data<=16'd9212;
      55999:data<=16'd8153;
      56000:data<=16'd5985;
      56001:data<=16'd4954;
      56002:data<=16'd4936;
      56003:data<=16'd4187;
      56004:data<=16'd3656;
      56005:data<=16'd3756;
      56006:data<=16'd2256;
      56007:data<=-16'd1809;
      56008:data<=-16'd4475;
      56009:data<=-16'd4249;
      56010:data<=-16'd4329;
      56011:data<=-16'd4350;
      56012:data<=-16'd4752;
      56013:data<=-16'd6487;
      56014:data<=-16'd6461;
      56015:data<=-16'd5971;
      56016:data<=-16'd6385;
      56017:data<=-16'd6253;
      56018:data<=-16'd7404;
      56019:data<=-16'd7031;
      56020:data<=-16'd5829;
      56021:data<=-16'd13165;
      56022:data<=-16'd23375;
      56023:data<=-16'd24736;
      56024:data<=-16'd22736;
      56025:data<=-16'd23387;
      56026:data<=-16'd23278;
      56027:data<=-16'd22424;
      56028:data<=-16'd22457;
      56029:data<=-16'd21325;
      56030:data<=-16'd19831;
      56031:data<=-16'd19882;
      56032:data<=-16'd19033;
      56033:data<=-16'd17681;
      56034:data<=-16'd17779;
      56035:data<=-16'd16842;
      56036:data<=-16'd15617;
      56037:data<=-16'd16045;
      56038:data<=-16'd16260;
      56039:data<=-16'd16301;
      56040:data<=-16'd15954;
      56041:data<=-16'd15267;
      56042:data<=-16'd15148;
      56043:data<=-16'd13831;
      56044:data<=-16'd13162;
      56045:data<=-16'd13432;
      56046:data<=-16'd11909;
      56047:data<=-16'd12107;
      56048:data<=-16'd10994;
      56049:data<=-16'd5691;
      56050:data<=-16'd5103;
      56051:data<=-16'd6053;
      56052:data<=-16'd4278;
      56053:data<=-16'd6149;
      56054:data<=-16'd2099;
      56055:data<=16'd10727;
      56056:data<=16'd14919;
      56057:data<=16'd12104;
      56058:data<=16'd12458;
      56059:data<=16'd12537;
      56060:data<=16'd11999;
      56061:data<=16'd12035;
      56062:data<=16'd10516;
      56063:data<=16'd8904;
      56064:data<=16'd8208;
      56065:data<=16'd7702;
      56066:data<=16'd7200;
      56067:data<=16'd6677;
      56068:data<=16'd6285;
      56069:data<=16'd5918;
      56070:data<=16'd6024;
      56071:data<=16'd5893;
      56072:data<=16'd5184;
      56073:data<=16'd5515;
      56074:data<=16'd5147;
      56075:data<=16'd3259;
      56076:data<=16'd2507;
      56077:data<=16'd2367;
      56078:data<=16'd2312;
      56079:data<=16'd2467;
      56080:data<=16'd1950;
      56081:data<=16'd1833;
      56082:data<=16'd1779;
      56083:data<=16'd1903;
      56084:data<=16'd2284;
      56085:data<=16'd873;
      56086:data<=16'd1300;
      56087:data<=16'd917;
      56088:data<=-16'd9066;
      56089:data<=-16'd18806;
      56090:data<=-16'd20016;
      56091:data<=-16'd21963;
      56092:data<=-16'd24386;
      56093:data<=-16'd23056;
      56094:data<=-16'd22075;
      56095:data<=-16'd21217;
      56096:data<=-16'd19851;
      56097:data<=-16'd19305;
      56098:data<=-16'd18406;
      56099:data<=-16'd17750;
      56100:data<=-16'd17782;
      56101:data<=-16'd17907;
      56102:data<=-16'd17616;
      56103:data<=-16'd16650;
      56104:data<=-16'd16480;
      56105:data<=-16'd16051;
      56106:data<=-16'd14828;
      56107:data<=-16'd14650;
      56108:data<=-16'd13631;
      56109:data<=-16'd11938;
      56110:data<=-16'd11300;
      56111:data<=-16'd10572;
      56112:data<=-16'd11006;
      56113:data<=-16'd11984;
      56114:data<=-16'd12016;
      56115:data<=-16'd12072;
      56116:data<=-16'd11041;
      56117:data<=-16'd10443;
      56118:data<=-16'd9899;
      56119:data<=-16'd8311;
      56120:data<=-16'd9761;
      56121:data<=-16'd5392;
      56122:data<=16'd8193;
      56123:data<=16'd12477;
      56124:data<=16'd8851;
      56125:data<=16'd9279;
      56126:data<=16'd8205;
      56127:data<=16'd7103;
      56128:data<=16'd8178;
      56129:data<=16'd6946;
      56130:data<=16'd7254;
      56131:data<=16'd7518;
      56132:data<=16'd6742;
      56133:data<=16'd10652;
      56134:data<=16'd13480;
      56135:data<=16'd12289;
      56136:data<=16'd12155;
      56137:data<=16'd11370;
      56138:data<=16'd9529;
      56139:data<=16'd8457;
      56140:data<=16'd8328;
      56141:data<=16'd9197;
      56142:data<=16'd8719;
      56143:data<=16'd7870;
      56144:data<=16'd8298;
      56145:data<=16'd8191;
      56146:data<=16'd8287;
      56147:data<=16'd8182;
      56148:data<=16'd7192;
      56149:data<=16'd7077;
      56150:data<=16'd6614;
      56151:data<=16'd4798;
      56152:data<=16'd3198;
      56153:data<=16'd3850;
      56154:data<=16'd3817;
      56155:data<=-16'd3667;
      56156:data<=-16'd11899;
      56157:data<=-16'd11728;
      56158:data<=-16'd10000;
      56159:data<=-16'd10011;
      56160:data<=-16'd8919;
      56161:data<=-16'd9021;
      56162:data<=-16'd9468;
      56163:data<=-16'd9512;
      56164:data<=-16'd9947;
      56165:data<=-16'd9024;
      56166:data<=-16'd8388;
      56167:data<=-16'd8426;
      56168:data<=-16'd7473;
      56169:data<=-16'd7043;
      56170:data<=-16'd7024;
      56171:data<=-16'd7062;
      56172:data<=-16'd7191;
      56173:data<=-16'd6314;
      56174:data<=-16'd6646;
      56175:data<=-16'd9794;
      56176:data<=-16'd12906;
      56177:data<=-16'd13224;
      56178:data<=-16'd11953;
      56179:data<=-16'd11400;
      56180:data<=-16'd10483;
      56181:data<=-16'd9938;
      56182:data<=-16'd10378;
      56183:data<=-16'd8992;
      56184:data<=-16'd8088;
      56185:data<=-16'd8049;
      56186:data<=-16'd7380;
      56187:data<=-16'd8997;
      56188:data<=-16'd4622;
      56189:data<=16'd7733;
      56190:data<=16'd11353;
      56191:data<=16'd8241;
      56192:data<=16'd9297;
      56193:data<=16'd9591;
      56194:data<=16'd9037;
      56195:data<=16'd9423;
      56196:data<=16'd8361;
      56197:data<=16'd8778;
      56198:data<=16'd8981;
      56199:data<=16'd7345;
      56200:data<=16'd7971;
      56201:data<=16'd9071;
      56202:data<=16'd8868;
      56203:data<=16'd9210;
      56204:data<=16'd9364;
      56205:data<=16'd9021;
      56206:data<=16'd8795;
      56207:data<=16'd8821;
      56208:data<=16'd8942;
      56209:data<=16'd8690;
      56210:data<=16'd8241;
      56211:data<=16'd7832;
      56212:data<=16'd8329;
      56213:data<=16'd9770;
      56214:data<=16'd10466;
      56215:data<=16'd9797;
      56216:data<=16'd9274;
      56217:data<=16'd11988;
      56218:data<=16'd15211;
      56219:data<=16'd14176;
      56220:data<=16'd14057;
      56221:data<=16'd13612;
      56222:data<=16'd5092;
      56223:data<=-16'd2773;
      56224:data<=-16'd2948;
      56225:data<=-16'd1654;
      56226:data<=-16'd205;
      56227:data<=16'd1081;
      56228:data<=16'd813;
      56229:data<=16'd887;
      56230:data<=16'd943;
      56231:data<=16'd1154;
      56232:data<=16'd1618;
      56233:data<=16'd1395;
      56234:data<=16'd1568;
      56235:data<=16'd1356;
      56236:data<=16'd1095;
      56237:data<=16'd2129;
      56238:data<=16'd3046;
      56239:data<=16'd3792;
      56240:data<=16'd3641;
      56241:data<=16'd3039;
      56242:data<=16'd3864;
      56243:data<=16'd3883;
      56244:data<=16'd3706;
      56245:data<=16'd4035;
      56246:data<=16'd2968;
      56247:data<=16'd2933;
      56248:data<=16'd2637;
      56249:data<=16'd1727;
      56250:data<=16'd3709;
      56251:data<=16'd4664;
      56252:data<=16'd5271;
      56253:data<=16'd6238;
      56254:data<=16'd3350;
      56255:data<=16'd7201;
      56256:data<=16'd18399;
      56257:data<=16'd20754;
      56258:data<=16'd17890;
      56259:data<=16'd15896;
      56260:data<=16'd11212;
      56261:data<=16'd9373;
      56262:data<=16'd10736;
      56263:data<=16'd10702;
      56264:data<=16'd11383;
      56265:data<=16'd11561;
      56266:data<=16'd10336;
      56267:data<=16'd9938;
      56268:data<=16'd9580;
      56269:data<=16'd8880;
      56270:data<=16'd8522;
      56271:data<=16'd8674;
      56272:data<=16'd8434;
      56273:data<=16'd7377;
      56274:data<=16'd7262;
      56275:data<=16'd7973;
      56276:data<=16'd8757;
      56277:data<=16'd9279;
      56278:data<=16'd8705;
      56279:data<=16'd8437;
      56280:data<=16'd8247;
      56281:data<=16'd7727;
      56282:data<=16'd7832;
      56283:data<=16'd6560;
      56284:data<=16'd5783;
      56285:data<=16'd6370;
      56286:data<=16'd5065;
      56287:data<=16'd6035;
      56288:data<=16'd6583;
      56289:data<=-16'd1005;
      56290:data<=-16'd7691;
      56291:data<=-16'd7691;
      56292:data<=-16'd6913;
      56293:data<=-16'd6310;
      56294:data<=-16'd6469;
      56295:data<=-16'd7075;
      56296:data<=-16'd6595;
      56297:data<=-16'd6599;
      56298:data<=-16'd5764;
      56299:data<=-16'd5136;
      56300:data<=-16'd5380;
      56301:data<=-16'd1401;
      56302:data<=16'd3454;
      56303:data<=16'd3974;
      56304:data<=16'd3433;
      56305:data<=16'd3121;
      56306:data<=16'd2813;
      56307:data<=16'd2723;
      56308:data<=16'd2194;
      56309:data<=16'd2223;
      56310:data<=16'd2390;
      56311:data<=16'd2376;
      56312:data<=16'd2619;
      56313:data<=16'd2927;
      56314:data<=16'd4194;
      56315:data<=16'd4193;
      56316:data<=16'd2986;
      56317:data<=16'd3823;
      56318:data<=16'd3688;
      56319:data<=16'd3374;
      56320:data<=16'd3891;
      56321:data<=16'd1174;
      56322:data<=16'd4640;
      56323:data<=16'd16072;
      56324:data<=16'd18683;
      56325:data<=16'd15784;
      56326:data<=16'd17274;
      56327:data<=16'd16666;
      56328:data<=16'd15308;
      56329:data<=16'd16158;
      56330:data<=16'd14522;
      56331:data<=16'd13227;
      56332:data<=16'd13667;
      56333:data<=16'd12762;
      56334:data<=16'd11764;
      56335:data<=16'd10922;
      56336:data<=16'd10439;
      56337:data<=16'd10715;
      56338:data<=16'd10630;
      56339:data<=16'd11166;
      56340:data<=16'd10960;
      56341:data<=16'd9612;
      56342:data<=16'd9793;
      56343:data<=16'd7702;
      56344:data<=16'd2737;
      56345:data<=16'd1306;
      56346:data<=16'd1853;
      56347:data<=16'd1427;
      56348:data<=16'd1774;
      56349:data<=16'd1274;
      56350:data<=16'd464;
      56351:data<=16'd1833;
      56352:data<=16'd2021;
      56353:data<=16'd667;
      56354:data<=16'd1522;
      56355:data<=-16'd27;
      56356:data<=-16'd8558;
      56357:data<=-16'd15593;
      56358:data<=-16'd15215;
      56359:data<=-16'd13717;
      56360:data<=-16'd13582;
      56361:data<=-16'd12571;
      56362:data<=-16'd12119;
      56363:data<=-16'd11641;
      56364:data<=-16'd10129;
      56365:data<=-16'd9482;
      56366:data<=-16'd9495;
      56367:data<=-16'd9635;
      56368:data<=-16'd9615;
      56369:data<=-16'd8690;
      56370:data<=-16'd8176;
      56371:data<=-16'd8105;
      56372:data<=-16'd7735;
      56373:data<=-16'd7837;
      56374:data<=-16'd7732;
      56375:data<=-16'd7121;
      56376:data<=-16'd6329;
      56377:data<=-16'd5372;
      56378:data<=-16'd5509;
      56379:data<=-16'd5850;
      56380:data<=-16'd5256;
      56381:data<=-16'd5401;
      56382:data<=-16'd5759;
      56383:data<=-16'd5356;
      56384:data<=-16'd5315;
      56385:data<=-16'd3759;
      56386:data<=16'd866;
      56387:data<=16'd2517;
      56388:data<=-16'd649;
      56389:data<=16'd3287;
      56390:data<=16'd14730;
      56391:data<=16'd17411;
      56392:data<=16'd13494;
      56393:data<=16'd13902;
      56394:data<=16'd13396;
      56395:data<=16'd11570;
      56396:data<=16'd12263;
      56397:data<=16'd10978;
      56398:data<=16'd9943;
      56399:data<=16'd11203;
      56400:data<=16'd9946;
      56401:data<=16'd7686;
      56402:data<=16'd6376;
      56403:data<=16'd5327;
      56404:data<=16'd5362;
      56405:data<=16'd4893;
      56406:data<=16'd3929;
      56407:data<=16'd3686;
      56408:data<=16'd3350;
      56409:data<=16'd3441;
      56410:data<=16'd3136;
      56411:data<=16'd2184;
      56412:data<=16'd2434;
      56413:data<=16'd2017;
      56414:data<=16'd230;
      56415:data<=-16'd552;
      56416:data<=-16'd904;
      56417:data<=-16'd1177;
      56418:data<=-16'd831;
      56419:data<=-16'd1378;
      56420:data<=-16'd1905;
      56421:data<=-16'd805;
      56422:data<=-16'd3093;
      56423:data<=-16'd11623;
      56424:data<=-16'd18083;
      56425:data<=-16'd17723;
      56426:data<=-16'd16859;
      56427:data<=-16'd19296;
      56428:data<=-16'd22441;
      56429:data<=-16'd23258;
      56430:data<=-16'd22058;
      56431:data<=-16'd21365;
      56432:data<=-16'd20741;
      56433:data<=-16'd19933;
      56434:data<=-16'd19960;
      56435:data<=-16'd19139;
      56436:data<=-16'd17696;
      56437:data<=-16'd17111;
      56438:data<=-16'd17270;
      56439:data<=-16'd18239;
      56440:data<=-16'd18174;
      56441:data<=-16'd17214;
      56442:data<=-16'd17032;
      56443:data<=-16'd16299;
      56444:data<=-16'd15932;
      56445:data<=-16'd15800;
      56446:data<=-16'd14433;
      56447:data<=-16'd13967;
      56448:data<=-16'd13543;
      56449:data<=-16'd13006;
      56450:data<=-16'd13634;
      56451:data<=-16'd13420;
      56452:data<=-16'd13975;
      56453:data<=-16'd13769;
      56454:data<=-16'd12166;
      56455:data<=-16'd14084;
      56456:data<=-16'd9583;
      56457:data<=16'd3209;
      56458:data<=16'd5958;
      56459:data<=16'd2525;
      56460:data<=16'd3883;
      56461:data<=16'd3667;
      56462:data<=16'd2813;
      56463:data<=16'd3189;
      56464:data<=16'd986;
      56465:data<=-16'd83;
      56466:data<=16'd1436;
      56467:data<=16'd1851;
      56468:data<=16'd563;
      56469:data<=16'd1295;
      56470:data<=16'd5545;
      56471:data<=16'd7277;
      56472:data<=16'd6024;
      56473:data<=16'd6197;
      56474:data<=16'd6018;
      56475:data<=16'd5586;
      56476:data<=16'd5134;
      56477:data<=16'd3595;
      56478:data<=16'd3415;
      56479:data<=16'd3497;
      56480:data<=16'd3319;
      56481:data<=16'd3835;
      56482:data<=16'd3298;
      56483:data<=16'd3430;
      56484:data<=16'd3680;
      56485:data<=16'd2799;
      56486:data<=16'd3052;
      56487:data<=16'd2779;
      56488:data<=16'd2328;
      56489:data<=-16'd937;
      56490:data<=-16'd10796;
      56491:data<=-16'd16336;
      56492:data<=-16'd14718;
      56493:data<=-16'd14613;
      56494:data<=-16'd13934;
      56495:data<=-16'd12783;
      56496:data<=-16'd12968;
      56497:data<=-16'd11667;
      56498:data<=-16'd11025;
      56499:data<=-16'd10593;
      56500:data<=-16'd10151;
      56501:data<=-16'd11488;
      56502:data<=-16'd11376;
      56503:data<=-16'd10883;
      56504:data<=-16'd10569;
      56505:data<=-16'd9150;
      56506:data<=-16'd9464;
      56507:data<=-16'd9406;
      56508:data<=-16'd8989;
      56509:data<=-16'd8863;
      56510:data<=-16'd6414;
      56511:data<=-16'd8241;
      56512:data<=-16'd13083;
      56513:data<=-16'd13444;
      56514:data<=-16'd14216;
      56515:data<=-16'd14877;
      56516:data<=-16'd13972;
      56517:data<=-16'd14316;
      56518:data<=-16'd12543;
      56519:data<=-16'd11919;
      56520:data<=-16'd12075;
      56521:data<=-16'd10064;
      56522:data<=-16'd12011;
      56523:data<=-16'd7658;
      56524:data<=16'd5480;
      56525:data<=16'd7397;
      56526:data<=16'd3198;
      56527:data<=16'd4202;
      56528:data<=16'd3930;
      56529:data<=16'd3838;
      56530:data<=16'd4552;
      56531:data<=16'd3430;
      56532:data<=16'd3381;
      56533:data<=16'd3498;
      56534:data<=16'd3883;
      56535:data<=16'd4114;
      56536:data<=16'd2786;
      56537:data<=16'd3043;
      56538:data<=16'd3021;
      56539:data<=16'd1545;
      56540:data<=16'd1395;
      56541:data<=16'd1111;
      56542:data<=16'd1086;
      56543:data<=16'd1504;
      56544:data<=16'd1292;
      56545:data<=16'd1541;
      56546:data<=16'd1221;
      56547:data<=16'd1579;
      56548:data<=16'd2564;
      56549:data<=16'd2046;
      56550:data<=16'd2837;
      56551:data<=16'd2358;
      56552:data<=-16'd447;
      56553:data<=16'd1207;
      56554:data<=16'd5462;
      56555:data<=16'd7896;
      56556:data<=16'd5236;
      56557:data<=-16'd4220;
      56558:data<=-16'd9567;
      56559:data<=-16'd7542;
      56560:data<=-16'd7163;
      56561:data<=-16'd7615;
      56562:data<=-16'd6951;
      56563:data<=-16'd7051;
      56564:data<=-16'd7288;
      56565:data<=-16'd7644;
      56566:data<=-16'd6680;
      56567:data<=-16'd5529;
      56568:data<=-16'd6029;
      56569:data<=-16'd5401;
      56570:data<=-16'd4599;
      56571:data<=-16'd4607;
      56572:data<=-16'd3999;
      56573:data<=-16'd4053;
      56574:data<=-16'd3738;
      56575:data<=-16'd3078;
      56576:data<=-16'd3621;
      56577:data<=-16'd3944;
      56578:data<=-16'd4338;
      56579:data<=-16'd4109;
      56580:data<=-16'd3181;
      56581:data<=-16'd3424;
      56582:data<=-16'd2869;
      56583:data<=-16'd2676;
      56584:data<=-16'd3281;
      56585:data<=-16'd1814;
      56586:data<=-16'd1770;
      56587:data<=-16'd1762;
      56588:data<=-16'd462;
      56589:data<=-16'd2670;
      56590:data<=16'd1685;
      56591:data<=16'd14139;
      56592:data<=16'd16117;
      56593:data<=16'd12107;
      56594:data<=16'd14228;
      56595:data<=16'd13223;
      56596:data<=16'd7905;
      56597:data<=16'd6320;
      56598:data<=16'd6253;
      56599:data<=16'd5398;
      56600:data<=16'd4983;
      56601:data<=16'd5611;
      56602:data<=16'd7376;
      56603:data<=16'd7670;
      56604:data<=16'd6300;
      56605:data<=16'd6407;
      56606:data<=16'd7072;
      56607:data<=16'd6778;
      56608:data<=16'd6704;
      56609:data<=16'd6437;
      56610:data<=16'd6014;
      56611:data<=16'd6155;
      56612:data<=16'd5642;
      56613:data<=16'd5554;
      56614:data<=16'd7042;
      56615:data<=16'd7908;
      56616:data<=16'd8070;
      56617:data<=16'd7940;
      56618:data<=16'd7166;
      56619:data<=16'd7225;
      56620:data<=16'd7004;
      56621:data<=16'd6667;
      56622:data<=16'd7938;
      56623:data<=16'd4576;
      56624:data<=-16'd4924;
      56625:data<=-16'd10096;
      56626:data<=-16'd8428;
      56627:data<=-16'd6340;
      56628:data<=-16'd5485;
      56629:data<=-16'd5128;
      56630:data<=-16'd5316;
      56631:data<=-16'd5071;
      56632:data<=-16'd4463;
      56633:data<=-16'd4126;
      56634:data<=-16'd3122;
      56635:data<=-16'd2458;
      56636:data<=-16'd3418;
      56637:data<=-16'd1621;
      56638:data<=16'd3721;
      56639:data<=16'd6310;
      56640:data<=16'd6319;
      56641:data<=16'd6593;
      56642:data<=16'd5982;
      56643:data<=16'd6196;
      56644:data<=16'd6837;
      56645:data<=16'd5727;
      56646:data<=16'd5559;
      56647:data<=16'd5929;
      56648:data<=16'd5642;
      56649:data<=16'd6024;
      56650:data<=16'd5175;
      56651:data<=16'd5124;
      56652:data<=16'd7326;
      56653:data<=16'd7122;
      56654:data<=16'd7078;
      56655:data<=16'd7677;
      56656:data<=16'd5049;
      56657:data<=16'd8809;
      56658:data<=16'd19829;
      56659:data<=16'd22694;
      56660:data<=16'd19370;
      56661:data<=16'd19183;
      56662:data<=16'd18827;
      56663:data<=16'd18215;
      56664:data<=16'd19102;
      56665:data<=16'd18553;
      56666:data<=16'd17787;
      56667:data<=16'd17764;
      56668:data<=16'd16751;
      56669:data<=16'd15755;
      56670:data<=16'd14789;
      56671:data<=16'd13518;
      56672:data<=16'd13500;
      56673:data<=16'd13670;
      56674:data<=16'd12995;
      56675:data<=16'd12771;
      56676:data<=16'd12299;
      56677:data<=16'd12113;
      56678:data<=16'd13447;
      56679:data<=16'd11659;
      56680:data<=16'd6193;
      56681:data<=16'd4144;
      56682:data<=16'd4949;
      56683:data<=16'd4460;
      56684:data<=16'd4064;
      56685:data<=16'd3842;
      56686:data<=16'd3797;
      56687:data<=16'd3845;
      56688:data<=16'd3489;
      56689:data<=16'd5391;
      56690:data<=16'd3626;
      56691:data<=-16'd6267;
      56692:data<=-16'd11459;
      56693:data<=-16'd9464;
      56694:data<=-16'd9749;
      56695:data<=-16'd9914;
      56696:data<=-16'd8963;
      56697:data<=-16'd9336;
      56698:data<=-16'd8407;
      56699:data<=-16'd7864;
      56700:data<=-16'd7990;
      56701:data<=-16'd6490;
      56702:data<=-16'd5354;
      56703:data<=-16'd4584;
      56704:data<=-16'd3983;
      56705:data<=-16'd4076;
      56706:data<=-16'd3742;
      56707:data<=-16'd3638;
      56708:data<=-16'd3609;
      56709:data<=-16'd3874;
      56710:data<=-16'd4214;
      56711:data<=-16'd3062;
      56712:data<=-16'd3169;
      56713:data<=-16'd3651;
      56714:data<=-16'd2006;
      56715:data<=-16'd1595;
      56716:data<=-16'd1553;
      56717:data<=-16'd1359;
      56718:data<=-16'd1704;
      56719:data<=-16'd720;
      56720:data<=-16'd1897;
      56721:data<=-16'd919;
      56722:data<=16'd4617;
      56723:data<=16'd4188;
      56724:data<=16'd7118;
      56725:data<=16'd19041;
      56726:data<=16'd21722;
      56727:data<=16'd19114;
      56728:data<=16'd20551;
      56729:data<=16'd19036;
      56730:data<=16'd18199;
      56731:data<=16'd18251;
      56732:data<=16'd15385;
      56733:data<=16'd15171;
      56734:data<=16'd15262;
      56735:data<=16'd13976;
      56736:data<=16'd14102;
      56737:data<=16'd12646;
      56738:data<=16'd11489;
      56739:data<=16'd12390;
      56740:data<=16'd12674;
      56741:data<=16'd12333;
      56742:data<=16'd11320;
      56743:data<=16'd10978;
      56744:data<=16'd10951;
      56745:data<=16'd9990;
      56746:data<=16'd9758;
      56747:data<=16'd8598;
      56748:data<=16'd7679;
      56749:data<=16'd8581;
      56750:data<=16'd7934;
      56751:data<=16'd8108;
      56752:data<=16'd9139;
      56753:data<=16'd8320;
      56754:data<=16'd8069;
      56755:data<=16'd7512;
      56756:data<=16'd7483;
      56757:data<=16'd4614;
      56758:data<=-16'd5773;
      56759:data<=-16'd10608;
      56760:data<=-16'd8413;
      56761:data<=-16'd9984;
      56762:data<=-16'd9351;
      56763:data<=-16'd8692;
      56764:data<=-16'd12680;
      56765:data<=-16'd12668;
      56766:data<=-16'd11831;
      56767:data<=-16'd12627;
      56768:data<=-16'd11185;
      56769:data<=-16'd11608;
      56770:data<=-16'd11841;
      56771:data<=-16'd10310;
      56772:data<=-16'd10389;
      56773:data<=-16'd9655;
      56774:data<=-16'd8984;
      56775:data<=-16'd9210;
      56776:data<=-16'd8475;
      56777:data<=-16'd7641;
      56778:data<=-16'd6467;
      56779:data<=-16'd6683;
      56780:data<=-16'd7066;
      56781:data<=-16'd5629;
      56782:data<=-16'd6300;
      56783:data<=-16'd6584;
      56784:data<=-16'd5741;
      56785:data<=-16'd7048;
      56786:data<=-16'd6481;
      56787:data<=-16'd5682;
      56788:data<=-16'd5482;
      56789:data<=-16'd4250;
      56790:data<=-16'd6103;
      56791:data<=-16'd1579;
      56792:data<=16'd10044;
      56793:data<=16'd11189;
      56794:data<=16'd7837;
      56795:data<=16'd9081;
      56796:data<=16'd8263;
      56797:data<=16'd7774;
      56798:data<=16'd7700;
      56799:data<=16'd5871;
      56800:data<=16'd6297;
      56801:data<=16'd5961;
      56802:data<=16'd4332;
      56803:data<=16'd3817;
      56804:data<=16'd2106;
      56805:data<=16'd2397;
      56806:data<=16'd6290;
      56807:data<=16'd8560;
      56808:data<=16'd7818;
      56809:data<=16'd6948;
      56810:data<=16'd7068;
      56811:data<=16'd6493;
      56812:data<=16'd6175;
      56813:data<=16'd6504;
      56814:data<=16'd4798;
      56815:data<=16'd3243;
      56816:data<=16'd3031;
      56817:data<=16'd2551;
      56818:data<=16'd2705;
      56819:data<=16'd2302;
      56820:data<=16'd2015;
      56821:data<=16'd1932;
      56822:data<=16'd849;
      56823:data<=16'd2188;
      56824:data<=-16'd923;
      56825:data<=-16'd11897;
      56826:data<=-16'd16066;
      56827:data<=-16'd14195;
      56828:data<=-16'd15403;
      56829:data<=-16'd15314;
      56830:data<=-16'd14583;
      56831:data<=-16'd14671;
      56832:data<=-16'd13479;
      56833:data<=-16'd13444;
      56834:data<=-16'd12963;
      56835:data<=-16'd11785;
      56836:data<=-16'd12264;
      56837:data<=-16'd11955;
      56838:data<=-16'd11118;
      56839:data<=-16'd11386;
      56840:data<=-16'd12273;
      56841:data<=-16'd12449;
      56842:data<=-16'd11235;
      56843:data<=-16'd11253;
      56844:data<=-16'd11330;
      56845:data<=-16'd10285;
      56846:data<=-16'd10348;
      56847:data<=-16'd10128;
      56848:data<=-16'd12592;
      56849:data<=-16'd16836;
      56850:data<=-16'd15634;
      56851:data<=-16'd14919;
      56852:data<=-16'd16807;
      56853:data<=-16'd16087;
      56854:data<=-16'd16210;
      56855:data<=-16'd15003;
      56856:data<=-16'd13370;
      56857:data<=-16'd14794;
      56858:data<=-16'd8364;
      56859:data<=16'd2256;
      56860:data<=16'd3620;
      56861:data<=16'd1742;
      56862:data<=16'd1935;
      56863:data<=16'd2156;
      56864:data<=16'd1791;
      56865:data<=16'd96;
      56866:data<=-16'd255;
      56867:data<=16'd96;
      56868:data<=-16'd649;
      56869:data<=-16'd372;
      56870:data<=-16'd563;
      56871:data<=-16'd1166;
      56872:data<=-16'd1031;
      56873:data<=-16'd1201;
      56874:data<=-16'd779;
      56875:data<=-16'd1037;
      56876:data<=-16'd1707;
      56877:data<=-16'd1924;
      56878:data<=-16'd3289;
      56879:data<=-16'd2855;
      56880:data<=-16'd2009;
      56881:data<=-16'd3016;
      56882:data<=-16'd2144;
      56883:data<=-16'd2102;
      56884:data<=-16'd2460;
      56885:data<=-16'd1184;
      56886:data<=-16'd2479;
      56887:data<=-16'd1994;
      56888:data<=-16'd1011;
      56889:data<=-16'd2887;
      56890:data<=16'd967;
      56891:data<=16'd875;
      56892:data<=-16'd10111;
      56893:data<=-16'd14169;
      56894:data<=-16'd11823;
      56895:data<=-16'd12179;
      56896:data<=-16'd11317;
      56897:data<=-16'd10869;
      56898:data<=-16'd10762;
      56899:data<=-16'd9439;
      56900:data<=-16'd9418;
      56901:data<=-16'd8624;
      56902:data<=-16'd8526;
      56903:data<=-16'd9912;
      56904:data<=-16'd9324;
      56905:data<=-16'd9013;
      56906:data<=-16'd8856;
      56907:data<=-16'd7624;
      56908:data<=-16'd7427;
      56909:data<=-16'd6951;
      56910:data<=-16'd6238;
      56911:data<=-16'd5937;
      56912:data<=-16'd5195;
      56913:data<=-16'd4901;
      56914:data<=-16'd4993;
      56915:data<=-16'd6416;
      56916:data<=-16'd7618;
      56917:data<=-16'd6231;
      56918:data<=-16'd6266;
      56919:data<=-16'd6745;
      56920:data<=-16'd5539;
      56921:data<=-16'd5718;
      56922:data<=-16'd4622;
      56923:data<=-16'd4087;
      56924:data<=-16'd5601;
      56925:data<=16'd1130;
      56926:data<=16'd11215;
      56927:data<=16'd11482;
      56928:data<=16'd8179;
      56929:data<=16'd8152;
      56930:data<=16'd8748;
      56931:data<=16'd8525;
      56932:data<=16'd5785;
      56933:data<=16'd1750;
      56934:data<=16'd626;
      56935:data<=16'd1459;
      56936:data<=16'd1353;
      56937:data<=16'd995;
      56938:data<=16'd876;
      56939:data<=-16'd2;
      56940:data<=-16'd798;
      56941:data<=-16'd1051;
      56942:data<=-16'd1148;
      56943:data<=-16'd757;
      56944:data<=-16'd1133;
      56945:data<=-16'd1300;
      56946:data<=-16'd56;
      56947:data<=-16'd325;
      56948:data<=-16'd591;
      56949:data<=16'd288;
      56950:data<=-16'd227;
      56951:data<=16'd523;
      56952:data<=16'd594;
      56953:data<=-16'd2093;
      56954:data<=-16'd1448;
      56955:data<=-16'd986;
      56956:data<=-16'd1983;
      56957:data<=16'd1295;
      56958:data<=-16'd1986;
      56959:data<=-16'd13421;
      56960:data<=-16'd16557;
      56961:data<=-16'd14245;
      56962:data<=-16'd14698;
      56963:data<=-16'd13887;
      56964:data<=-16'd13270;
      56965:data<=-16'd14155;
      56966:data<=-16'd13535;
      56967:data<=-16'd12583;
      56968:data<=-16'd11714;
      56969:data<=-16'd10951;
      56970:data<=-16'd10596;
      56971:data<=-16'd9018;
      56972:data<=-16'd8258;
      56973:data<=-16'd9051;
      56974:data<=-16'd6288;
      56975:data<=-16'd949;
      56976:data<=16'd447;
      56977:data<=-16'd1321;
      56978:data<=-16'd2036;
      56979:data<=-16'd1856;
      56980:data<=-16'd1304;
      56981:data<=-16'd842;
      56982:data<=-16'd1356;
      56983:data<=-16'd1037;
      56984:data<=-16'd281;
      56985:data<=-16'd819;
      56986:data<=-16'd487;
      56987:data<=-16'd39;
      56988:data<=-16'd560;
      56989:data<=16'd535;
      56990:data<=16'd328;
      56991:data<=-16'd349;
      56992:data<=16'd6678;
      56993:data<=16'd15590;
      56994:data<=16'd16252;
      56995:data<=16'd14377;
      56996:data<=16'd15208;
      56997:data<=16'd15430;
      56998:data<=16'd14660;
      56999:data<=16'd13937;
      57000:data<=16'd12837;
      57001:data<=16'd11941;
      57002:data<=16'd11981;
      57003:data<=16'd13032;
      57004:data<=16'd13664;
      57005:data<=16'd12869;
      57006:data<=16'd12184;
      57007:data<=16'd11878;
      57008:data<=16'd11377;
      57009:data<=16'd11646;
      57010:data<=16'd11520;
      57011:data<=16'd10243;
      57012:data<=16'd10120;
      57013:data<=16'd10055;
      57014:data<=16'd9309;
      57015:data<=16'd10739;
      57016:data<=16'd10251;
      57017:data<=16'd5225;
      57018:data<=16'd3697;
      57019:data<=16'd5285;
      57020:data<=16'd4285;
      57021:data<=16'd4185;
      57022:data<=16'd3820;
      57023:data<=16'd2658;
      57024:data<=16'd5529;
      57025:data<=16'd2259;
      57026:data<=-16'd9784;
      57027:data<=-16'd12753;
      57028:data<=-16'd8228;
      57029:data<=-16'd8370;
      57030:data<=-16'd8540;
      57031:data<=-16'd7127;
      57032:data<=-16'd7222;
      57033:data<=-16'd6552;
      57034:data<=-16'd5812;
      57035:data<=-16'd5421;
      57036:data<=-16'd4701;
      57037:data<=-16'd4877;
      57038:data<=-16'd4687;
      57039:data<=-16'd4026;
      57040:data<=-16'd3371;
      57041:data<=-16'd1689;
      57042:data<=-16'd1019;
      57043:data<=-16'd1706;
      57044:data<=-16'd1471;
      57045:data<=-16'd1137;
      57046:data<=-16'd1316;
      57047:data<=-16'd1133;
      57048:data<=-16'd616;
      57049:data<=-16'd5;
      57050:data<=16'd58;
      57051:data<=-16'd549;
      57052:data<=16'd82;
      57053:data<=16'd1959;
      57054:data<=16'd1905;
      57055:data<=16'd1671;
      57056:data<=16'd3212;
      57057:data<=16'd1428;
      57058:data<=16'd2276;
      57059:data<=16'd14744;
      57060:data<=16'd24577;
      57061:data<=16'd22650;
      57062:data<=16'd20747;
      57063:data<=16'd21215;
      57064:data<=16'd20624;
      57065:data<=16'd20979;
      57066:data<=16'd20639;
      57067:data<=16'd19391;
      57068:data<=16'd18619;
      57069:data<=16'd17697;
      57070:data<=16'd17443;
      57071:data<=16'd17041;
      57072:data<=16'd15884;
      57073:data<=16'd14889;
      57074:data<=16'd13919;
      57075:data<=16'd13474;
      57076:data<=16'd13098;
      57077:data<=16'd13080;
      57078:data<=16'd13744;
      57079:data<=16'd13191;
      57080:data<=16'd12747;
      57081:data<=16'd12554;
      57082:data<=16'd11220;
      57083:data<=16'd10851;
      57084:data<=16'd10605;
      57085:data<=16'd10404;
      57086:data<=16'd10793;
      57087:data<=16'd9388;
      57088:data<=16'd8799;
      57089:data<=16'd8363;
      57090:data<=16'd7870;
      57091:data<=16'd11532;
      57092:data<=16'd7981;
      57093:data<=-16'd4440;
      57094:data<=-16'd7517;
      57095:data<=-16'd4889;
      57096:data<=-16'd6041;
      57097:data<=-16'd6419;
      57098:data<=-16'd6484;
      57099:data<=-16'd5600;
      57100:data<=-16'd6038;
      57101:data<=-16'd11239;
      57102:data<=-16'd11875;
      57103:data<=-16'd8573;
      57104:data<=-16'd8528;
      57105:data<=-16'd7846;
      57106:data<=-16'd7241;
      57107:data<=-16'd7971;
      57108:data<=-16'd7269;
      57109:data<=-16'd6824;
      57110:data<=-16'd6783;
      57111:data<=-16'd7186;
      57112:data<=-16'd7565;
      57113:data<=-16'd6670;
      57114:data<=-16'd6699;
      57115:data<=-16'd5651;
      57116:data<=-16'd3324;
      57117:data<=-16'd3327;
      57118:data<=-16'd3266;
      57119:data<=-16'd3146;
      57120:data<=-16'd3714;
      57121:data<=-16'd3348;
      57122:data<=-16'd3645;
      57123:data<=-16'd3189;
      57124:data<=-16'd3039;
      57125:data<=-16'd2725;
      57126:data<=16'd5053;
      57127:data<=16'd13060;
      57128:data<=16'd13400;
      57129:data<=16'd13150;
      57130:data<=16'd12892;
      57131:data<=16'd11996;
      57132:data<=16'd12524;
      57133:data<=16'd11277;
      57134:data<=16'd10102;
      57135:data<=16'd9758;
      57136:data<=16'd8510;
      57137:data<=16'd8807;
      57138:data<=16'd8479;
      57139:data<=16'd7656;
      57140:data<=16'd8558;
      57141:data<=16'd8122;
      57142:data<=16'd9596;
      57143:data<=16'd14302;
      57144:data<=16'd15262;
      57145:data<=16'd13015;
      57146:data<=16'd12336;
      57147:data<=16'd12704;
      57148:data<=16'd11699;
      57149:data<=16'd10548;
      57150:data<=16'd10813;
      57151:data<=16'd9912;
      57152:data<=16'd9647;
      57153:data<=16'd11215;
      57154:data<=16'd10542;
      57155:data<=16'd10096;
      57156:data<=16'd9624;
      57157:data<=16'd7888;
      57158:data<=16'd9454;
      57159:data<=16'd5248;
      57160:data<=-16'd6681;
      57161:data<=-16'd9544;
      57162:data<=-16'd6672;
      57163:data<=-16'd8025;
      57164:data<=-16'd7999;
      57165:data<=-16'd6458;
      57166:data<=-16'd5512;
      57167:data<=-16'd4363;
      57168:data<=-16'd4640;
      57169:data<=-16'd4554;
      57170:data<=-16'd4099;
      57171:data<=-16'd4417;
      57172:data<=-16'd3955;
      57173:data<=-16'd4090;
      57174:data<=-16'd4491;
      57175:data<=-16'd4185;
      57176:data<=-16'd4666;
      57177:data<=-16'd4447;
      57178:data<=-16'd3287;
      57179:data<=-16'd2693;
      57180:data<=-16'd2428;
      57181:data<=-16'd2911;
      57182:data<=-16'd2983;
      57183:data<=-16'd2223;
      57184:data<=-16'd4021;
      57185:data<=-16'd8464;
      57186:data<=-16'd10440;
      57187:data<=-16'd8821;
      57188:data<=-16'd8628;
      57189:data<=-16'd9216;
      57190:data<=-16'd7808;
      57191:data<=-16'd8693;
      57192:data<=-16'd7850;
      57193:data<=16'd986;
      57194:data<=16'd7649;
      57195:data<=16'd6996;
      57196:data<=16'd5906;
      57197:data<=16'd5366;
      57198:data<=16'd5297;
      57199:data<=16'd6075;
      57200:data<=16'd5230;
      57201:data<=16'd3997;
      57202:data<=16'd3416;
      57203:data<=16'd2097;
      57204:data<=16'd978;
      57205:data<=16'd876;
      57206:data<=16'd544;
      57207:data<=-16'd288;
      57208:data<=-16'd215;
      57209:data<=16'd176;
      57210:data<=16'd77;
      57211:data<=16'd502;
      57212:data<=-16'd6;
      57213:data<=-16'd839;
      57214:data<=-16'd20;
      57215:data<=-16'd1030;
      57216:data<=-16'd3060;
      57217:data<=-16'd2766;
      57218:data<=-16'd2664;
      57219:data<=-16'd2453;
      57220:data<=-16'd1994;
      57221:data<=-16'd2936;
      57222:data<=-16'd2717;
      57223:data<=-16'd2472;
      57224:data<=-16'd2611;
      57225:data<=-16'd1359;
      57226:data<=-16'd4686;
      57227:data<=-16'd11417;
      57228:data<=-16'd13038;
      57229:data<=-16'd12411;
      57230:data<=-16'd12994;
      57231:data<=-16'd12466;
      57232:data<=-16'd11919;
      57233:data<=-16'd11700;
      57234:data<=-16'd10837;
      57235:data<=-16'd10349;
      57236:data<=-16'd10032;
      57237:data<=-16'd9505;
      57238:data<=-16'd9113;
      57239:data<=-16'd8419;
      57240:data<=-16'd8443;
      57241:data<=-16'd10234;
      57242:data<=-16'd11069;
      57243:data<=-16'd10132;
      57244:data<=-16'd10249;
      57245:data<=-16'd10255;
      57246:data<=-16'd9312;
      57247:data<=-16'd9297;
      57248:data<=-16'd8272;
      57249:data<=-16'd7228;
      57250:data<=-16'd8276;
      57251:data<=-16'd7653;
      57252:data<=-16'd6833;
      57253:data<=-16'd8429;
      57254:data<=-16'd8995;
      57255:data<=-16'd9150;
      57256:data<=-16'd8887;
      57257:data<=-16'd7326;
      57258:data<=-16'd8085;
      57259:data<=-16'd6498;
      57260:data<=16'd2171;
      57261:data<=16'd8828;
      57262:data<=16'd8376;
      57263:data<=16'd6948;
      57264:data<=16'd7430;
      57265:data<=16'd6449;
      57266:data<=16'd4325;
      57267:data<=16'd4426;
      57268:data<=16'd2773;
      57269:data<=-16'd2355;
      57270:data<=-16'd4059;
      57271:data<=-16'd2998;
      57272:data<=-16'd3263;
      57273:data<=-16'd3087;
      57274:data<=-16'd3248;
      57275:data<=-16'd3915;
      57276:data<=-16'd2977;
      57277:data<=-16'd1891;
      57278:data<=-16'd2359;
      57279:data<=-16'd4385;
      57280:data<=-16'd5190;
      57281:data<=-16'd3603;
      57282:data<=-16'd3389;
      57283:data<=-16'd3571;
      57284:data<=-16'd2805;
      57285:data<=-16'd3256;
      57286:data<=-16'd2460;
      57287:data<=-16'd1659;
      57288:data<=-16'd2604;
      57289:data<=-16'd1629;
      57290:data<=-16'd2908;
      57291:data<=-16'd5485;
      57292:data<=-16'd3127;
      57293:data<=-16'd7077;
      57294:data<=-16'd18550;
      57295:data<=-16'd20811;
      57296:data<=-16'd17259;
      57297:data<=-16'd17643;
      57298:data<=-16'd17315;
      57299:data<=-16'd15987;
      57300:data<=-16'd15970;
      57301:data<=-16'd14630;
      57302:data<=-16'd13016;
      57303:data<=-16'd13297;
      57304:data<=-16'd13884;
      57305:data<=-16'd13464;
      57306:data<=-16'd12652;
      57307:data<=-16'd11461;
      57308:data<=-16'd10519;
      57309:data<=-16'd11015;
      57310:data<=-16'd9376;
      57311:data<=-16'd4557;
      57312:data<=-16'd2657;
      57313:data<=-16'd3213;
      57314:data<=-16'd2284;
      57315:data<=-16'd2259;
      57316:data<=-16'd3416;
      57317:data<=-16'd3776;
      57318:data<=-16'd3802;
      57319:data<=-16'd3477;
      57320:data<=-16'd2831;
      57321:data<=-16'd2458;
      57322:data<=-16'd3024;
      57323:data<=-16'd2914;
      57324:data<=-16'd1389;
      57325:data<=-16'd2622;
      57326:data<=-16'd1566;
      57327:data<=16'd8223;
      57328:data<=16'd14325;
      57329:data<=16'd11532;
      57330:data<=16'd10425;
      57331:data<=16'd10816;
      57332:data<=16'd10281;
      57333:data<=16'd10801;
      57334:data<=16'd9805;
      57335:data<=16'd8696;
      57336:data<=16'd9006;
      57337:data<=16'd8023;
      57338:data<=16'd7219;
      57339:data<=16'd7550;
      57340:data<=16'd7247;
      57341:data<=16'd5894;
      57342:data<=16'd4585;
      57343:data<=16'd4981;
      57344:data<=16'd5683;
      57345:data<=16'd5635;
      57346:data<=16'd5482;
      57347:data<=16'd4707;
      57348:data<=16'd4916;
      57349:data<=16'd5009;
      57350:data<=16'd3550;
      57351:data<=16'd4117;
      57352:data<=16'd3380;
      57353:data<=-16'd1478;
      57354:data<=-16'd4232;
      57355:data<=-16'd4002;
      57356:data<=-16'd3559;
      57357:data<=-16'd4170;
      57358:data<=-16'd4387;
      57359:data<=-16'd1882;
      57360:data<=-16'd5903;
      57361:data<=-16'd16986;
      57362:data<=-16'd19387;
      57363:data<=-16'd16231;
      57364:data<=-16'd16521;
      57365:data<=-16'd15634;
      57366:data<=-16'd15338;
      57367:data<=-16'd16120;
      57368:data<=-16'd14157;
      57369:data<=-16'd13353;
      57370:data<=-16'd13323;
      57371:data<=-16'd11752;
      57372:data<=-16'd10860;
      57373:data<=-16'd9909;
      57374:data<=-16'd9247;
      57375:data<=-16'd9517;
      57376:data<=-16'd9095;
      57377:data<=-16'd8722;
      57378:data<=-16'd9034;
      57379:data<=-16'd9582;
      57380:data<=-16'd9532;
      57381:data<=-16'd8639;
      57382:data<=-16'd8214;
      57383:data<=-16'd7750;
      57384:data<=-16'd7171;
      57385:data<=-16'd6880;
      57386:data<=-16'd5893;
      57387:data<=-16'd5304;
      57388:data<=-16'd5244;
      57389:data<=-16'd5060;
      57390:data<=-16'd4411;
      57391:data<=-16'd2701;
      57392:data<=-16'd3419;
      57393:data<=-16'd2181;
      57394:data<=16'd9000;
      57395:data<=16'd19027;
      57396:data<=16'd19717;
      57397:data<=16'd19042;
      57398:data<=16'd18363;
      57399:data<=16'd17048;
      57400:data<=16'd17095;
      57401:data<=16'd16389;
      57402:data<=16'd15614;
      57403:data<=16'd15728;
      57404:data<=16'd15964;
      57405:data<=16'd16190;
      57406:data<=16'd15277;
      57407:data<=16'd14932;
      57408:data<=16'd14918;
      57409:data<=16'd13467;
      57410:data<=16'd13644;
      57411:data<=16'd14396;
      57412:data<=16'd13385;
      57413:data<=16'd12654;
      57414:data<=16'd12170;
      57415:data<=16'd12511;
      57416:data<=16'd13514;
      57417:data<=16'd13488;
      57418:data<=16'd13450;
      57419:data<=16'd12889;
      57420:data<=16'd12231;
      57421:data<=16'd12003;
      57422:data<=16'd11154;
      57423:data<=16'd11489;
      57424:data<=16'd10554;
      57425:data<=16'd9371;
      57426:data<=16'd11963;
      57427:data<=16'd7025;
      57428:data<=-16'd4332;
      57429:data<=-16'd5062;
      57430:data<=-16'd2005;
      57431:data<=-16'd3626;
      57432:data<=-16'd2877;
      57433:data<=-16'd2502;
      57434:data<=-16'd3507;
      57435:data<=-16'd1665;
      57436:data<=-16'd2529;
      57437:data<=-16'd6995;
      57438:data<=-16'd8668;
      57439:data<=-16'd7652;
      57440:data<=-16'd7027;
      57441:data<=-16'd6134;
      57442:data<=-16'd4373;
      57443:data<=-16'd3974;
      57444:data<=-16'd4491;
      57445:data<=-16'd4199;
      57446:data<=-16'd4162;
      57447:data<=-16'd3947;
      57448:data<=-16'd3582;
      57449:data<=-16'd3667;
      57450:data<=-16'd2746;
      57451:data<=-16'd2206;
      57452:data<=-16'd2705;
      57453:data<=-16'd1976;
      57454:data<=-16'd156;
      57455:data<=16'd951;
      57456:data<=16'd267;
      57457:data<=16'd667;
      57458:data<=16'd1770;
      57459:data<=-16'd675;
      57460:data<=16'd1780;
      57461:data<=16'd12091;
      57462:data<=16'd16283;
      57463:data<=16'd14821;
      57464:data<=16'd14945;
      57465:data<=16'd13703;
      57466:data<=16'd13496;
      57467:data<=16'd14865;
      57468:data<=16'd14041;
      57469:data<=16'd13612;
      57470:data<=16'd13280;
      57471:data<=16'd12005;
      57472:data<=16'd11866;
      57473:data<=16'd11674;
      57474:data<=16'd11239;
      57475:data<=16'd11182;
      57476:data<=16'd10636;
      57477:data<=16'd9917;
      57478:data<=16'd11166;
      57479:data<=16'd15676;
      57480:data<=16'd18098;
      57481:data<=16'd16431;
      57482:data<=16'd16219;
      57483:data<=16'd15725;
      57484:data<=16'd13863;
      57485:data<=16'd13969;
      57486:data<=16'd13100;
      57487:data<=16'd11953;
      57488:data<=16'd12316;
      57489:data<=16'd11549;
      57490:data<=16'd11177;
      57491:data<=16'd10660;
      57492:data<=16'd11201;
      57493:data<=16'd13932;
      57494:data<=16'd8176;
      57495:data<=-16'd3348;
      57496:data<=-16'd5894;
      57497:data<=-16'd4018;
      57498:data<=-16'd4607;
      57499:data<=-16'd4491;
      57500:data<=-16'd4309;
      57501:data<=-16'd4323;
      57502:data<=-16'd3764;
      57503:data<=-16'd3506;
      57504:data<=-16'd2749;
      57505:data<=-16'd1833;
      57506:data<=-16'd1296;
      57507:data<=-16'd974;
      57508:data<=-16'd1378;
      57509:data<=-16'd1782;
      57510:data<=-16'd1528;
      57511:data<=-16'd1431;
      57512:data<=-16'd2161;
      57513:data<=-16'd2393;
      57514:data<=-16'd1807;
      57515:data<=-16'd2413;
      57516:data<=-16'd1999;
      57517:data<=16'd59;
      57518:data<=-16'd171;
      57519:data<=-16'd352;
      57520:data<=-16'd49;
      57521:data<=-16'd2631;
      57522:data<=-16'd4570;
      57523:data<=-16'd4890;
      57524:data<=-16'd4491;
      57525:data<=-16'd3254;
      57526:data<=-16'd4875;
      57527:data<=-16'd2766;
      57528:data<=16'd7718;
      57529:data<=16'd13614;
      57530:data<=16'd12686;
      57531:data<=16'd12516;
      57532:data<=16'd11535;
      57533:data<=16'd10252;
      57534:data<=16'd9993;
      57535:data<=16'd9389;
      57536:data<=16'd9210;
      57537:data<=16'd8210;
      57538:data<=16'd7520;
      57539:data<=16'd8270;
      57540:data<=16'd7514;
      57541:data<=16'd7401;
      57542:data<=16'd8728;
      57543:data<=16'd8345;
      57544:data<=16'd8020;
      57545:data<=16'd8202;
      57546:data<=16'd7453;
      57547:data<=16'd6886;
      57548:data<=16'd6731;
      57549:data<=16'd6623;
      57550:data<=16'd5824;
      57551:data<=16'd5054;
      57552:data<=16'd4984;
      57553:data<=16'd4143;
      57554:data<=16'd4708;
      57555:data<=16'd6031;
      57556:data<=16'd5230;
      57557:data<=16'd5864;
      57558:data<=16'd5702;
      57559:data<=16'd4044;
      57560:data<=16'd6205;
      57561:data<=16'd1680;
      57562:data<=-16'd10249;
      57563:data<=-16'd10574;
      57564:data<=-16'd4948;
      57565:data<=-16'd6026;
      57566:data<=-16'd5826;
      57567:data<=-16'd3750;
      57568:data<=-16'd4074;
      57569:data<=-16'd3559;
      57570:data<=-16'd3318;
      57571:data<=-16'd3868;
      57572:data<=-16'd3621;
      57573:data<=-16'd3836;
      57574:data<=-16'd3883;
      57575:data<=-16'd3747;
      57576:data<=-16'd4065;
      57577:data<=-16'd4015;
      57578:data<=-16'd4050;
      57579:data<=-16'd3377;
      57580:data<=-16'd1967;
      57581:data<=-16'd2235;
      57582:data<=-16'd2969;
      57583:data<=-16'd2264;
      57584:data<=-16'd1859;
      57585:data<=-16'd2284;
      57586:data<=-16'd2420;
      57587:data<=-16'd2587;
      57588:data<=-16'd2399;
      57589:data<=-16'd1848;
      57590:data<=-16'd2769;
      57591:data<=-16'd3136;
      57592:data<=-16'd2490;
      57593:data<=-16'd4285;
      57594:data<=-16'd1453;
      57595:data<=16'd8900;
      57596:data<=16'd12863;
      57597:data<=16'd10211;
      57598:data<=16'd10616;
      57599:data<=16'd10019;
      57600:data<=16'd7909;
      57601:data<=16'd7934;
      57602:data<=16'd7084;
      57603:data<=16'd6290;
      57604:data<=16'd5304;
      57605:data<=16'd1513;
      57606:data<=-16'd1274;
      57607:data<=-16'd1450;
      57608:data<=-16'd1077;
      57609:data<=-16'd1004;
      57610:data<=-16'd1568;
      57611:data<=-16'd1466;
      57612:data<=-16'd989;
      57613:data<=-16'd1186;
      57614:data<=-16'd1383;
      57615:data<=-16'd1707;
      57616:data<=-16'd2261;
      57617:data<=-16'd3704;
      57618:data<=-16'd4901;
      57619:data<=-16'd4147;
      57620:data<=-16'd4285;
      57621:data<=-16'd4642;
      57622:data<=-16'd3899;
      57623:data<=-16'd4598;
      57624:data<=-16'd4338;
      57625:data<=-16'd4173;
      57626:data<=-16'd5010;
      57627:data<=-16'd2726;
      57628:data<=-16'd6993;
      57629:data<=-16'd19376;
      57630:data<=-16'd22732;
      57631:data<=-16'd19478;
      57632:data<=-16'd19220;
      57633:data<=-16'd18305;
      57634:data<=-16'd17758;
      57635:data<=-16'd17635;
      57636:data<=-16'd15752;
      57637:data<=-16'd15305;
      57638:data<=-16'd15239;
      57639:data<=-16'd14542;
      57640:data<=-16'd14324;
      57641:data<=-16'd13799;
      57642:data<=-16'd14675;
      57643:data<=-16'd15540;
      57644:data<=-16'd14346;
      57645:data<=-16'd14322;
      57646:data<=-16'd14431;
      57647:data<=-16'd11775;
      57648:data<=-16'd9009;
      57649:data<=-16'd8170;
      57650:data<=-16'd7368;
      57651:data<=-16'd6305;
      57652:data<=-16'd6649;
      57653:data<=-16'd6855;
      57654:data<=-16'd6916;
      57655:data<=-16'd8228;
      57656:data<=-16'd8182;
      57657:data<=-16'd7891;
      57658:data<=-16'd7744;
      57659:data<=-16'd6219;
      57660:data<=-16'd7650;
      57661:data<=-16'd5228;
      57662:data<=16'd5961;
      57663:data<=16'd10229;
      57664:data<=16'd7482;
      57665:data<=16'd8449;
      57666:data<=16'd7470;
      57667:data<=16'd4576;
      57668:data<=16'd4009;
      57669:data<=16'd3448;
      57670:data<=16'd3674;
      57671:data<=16'd3330;
      57672:data<=16'd2833;
      57673:data<=16'd3909;
      57674:data<=16'd3347;
      57675:data<=16'd3289;
      57676:data<=16'd3941;
      57677:data<=16'd2863;
      57678:data<=16'd3415;
      57679:data<=16'd3221;
      57680:data<=16'd999;
      57681:data<=16'd681;
      57682:data<=16'd569;
      57683:data<=16'd305;
      57684:data<=16'd152;
      57685:data<=-16'd206;
      57686:data<=16'd485;
      57687:data<=16'd17;
      57688:data<=-16'd9;
      57689:data<=-16'd91;
      57690:data<=-16'd3612;
      57691:data<=-16'd4705;
      57692:data<=-16'd5009;
      57693:data<=-16'd6586;
      57694:data<=-16'd4055;
      57695:data<=-16'd8357;
      57696:data<=-16'd19635;
      57697:data<=-16'd20909;
      57698:data<=-16'd18117;
      57699:data<=-16'd18219;
      57700:data<=-16'd16290;
      57701:data<=-16'd15869;
      57702:data<=-16'd16172;
      57703:data<=-16'd14462;
      57704:data<=-16'd13976;
      57705:data<=-16'd14410;
      57706:data<=-16'd15139;
      57707:data<=-16'd14833;
      57708:data<=-16'd13142;
      57709:data<=-16'd12624;
      57710:data<=-16'd12122;
      57711:data<=-16'd11952;
      57712:data<=-16'd12384;
      57713:data<=-16'd11176;
      57714:data<=-16'd10117;
      57715:data<=-16'd9755;
      57716:data<=-16'd9397;
      57717:data<=-16'd9398;
      57718:data<=-16'd8928;
      57719:data<=-16'd8924;
      57720:data<=-16'd8640;
      57721:data<=-16'd8062;
      57722:data<=-16'd8308;
      57723:data<=-16'd7295;
      57724:data<=-16'd7166;
      57725:data<=-16'd6846;
      57726:data<=-16'd5125;
      57727:data<=-16'd7556;
      57728:data<=-16'd3985;
      57729:data<=16'd8032;
      57730:data<=16'd9573;
      57731:data<=16'd7147;
      57732:data<=16'd11794;
      57733:data<=16'd12540;
      57734:data<=16'd10681;
      57735:data<=16'd10813;
      57736:data<=16'd9982;
      57737:data<=16'd10144;
      57738:data<=16'd9611;
      57739:data<=16'd8745;
      57740:data<=16'd9409;
      57741:data<=16'd8649;
      57742:data<=16'd8034;
      57743:data<=16'd7083;
      57744:data<=16'd5644;
      57745:data<=16'd6596;
      57746:data<=16'd6401;
      57747:data<=16'd5776;
      57748:data<=16'd6385;
      57749:data<=16'd5457;
      57750:data<=16'd5363;
      57751:data<=16'd5039;
      57752:data<=16'd4338;
      57753:data<=16'd5827;
      57754:data<=16'd4655;
      57755:data<=16'd2822;
      57756:data<=16'd3256;
      57757:data<=16'd2499;
      57758:data<=16'd3068;
      57759:data<=16'd2846;
      57760:data<=16'd2093;
      57761:data<=16'd4525;
      57762:data<=-16'd970;
      57763:data<=-16'd11712;
      57764:data<=-16'd12634;
      57765:data<=-16'd10157;
      57766:data<=-16'd10596;
      57767:data<=-16'd11004;
      57768:data<=-16'd11740;
      57769:data<=-16'd10933;
      57770:data<=-16'd10052;
      57771:data<=-16'd10075;
      57772:data<=-16'd8569;
      57773:data<=-16'd9418;
      57774:data<=-16'd12192;
      57775:data<=-16'd12188;
      57776:data<=-16'd11063;
      57777:data<=-16'd10304;
      57778:data<=-16'd9970;
      57779:data<=-16'd10386;
      57780:data<=-16'd10822;
      57781:data<=-16'd10624;
      57782:data<=-16'd9832;
      57783:data<=-16'd9467;
      57784:data<=-16'd8326;
      57785:data<=-16'd6763;
      57786:data<=-16'd7131;
      57787:data<=-16'd6754;
      57788:data<=-16'd6052;
      57789:data<=-16'd6408;
      57790:data<=-16'd5248;
      57791:data<=-16'd5432;
      57792:data<=-16'd5189;
      57793:data<=-16'd2854;
      57794:data<=-16'd4628;
      57795:data<=-16'd1486;
      57796:data<=16'd10096;
      57797:data<=16'd13429;
      57798:data<=16'd10813;
      57799:data<=16'd11750;
      57800:data<=16'd11386;
      57801:data<=16'd10696;
      57802:data<=16'd10971;
      57803:data<=16'd9993;
      57804:data<=16'd10354;
      57805:data<=16'd11233;
      57806:data<=16'd11286;
      57807:data<=16'd11259;
      57808:data<=16'd11062;
      57809:data<=16'd11600;
      57810:data<=16'd10909;
      57811:data<=16'd9439;
      57812:data<=16'd10487;
      57813:data<=16'd10972;
      57814:data<=16'd9964;
      57815:data<=16'd11054;
      57816:data<=16'd13312;
      57817:data<=16'd14198;
      57818:data<=16'd14145;
      57819:data<=16'd14612;
      57820:data<=16'd14131;
      57821:data<=16'd12605;
      57822:data<=16'd13117;
      57823:data<=16'd13127;
      57824:data<=16'd11694;
      57825:data<=16'd12164;
      57826:data<=16'd11715;
      57827:data<=16'd11268;
      57828:data<=16'd12132;
      57829:data<=16'd6308;
      57830:data<=-16'd2408;
      57831:data<=-16'd3527;
      57832:data<=-16'd1809;
      57833:data<=-16'd2100;
      57834:data<=-16'd1798;
      57835:data<=-16'd1745;
      57836:data<=-16'd2231;
      57837:data<=-16'd1377;
      57838:data<=-16'd546;
      57839:data<=-16'd870;
      57840:data<=-16'd919;
      57841:data<=-16'd722;
      57842:data<=-16'd159;
      57843:data<=16'd1601;
      57844:data<=16'd2177;
      57845:data<=16'd1202;
      57846:data<=16'd992;
      57847:data<=16'd854;
      57848:data<=16'd1318;
      57849:data<=16'd2050;
      57850:data<=16'd1289;
      57851:data<=16'd1776;
      57852:data<=16'd2491;
      57853:data<=16'd1416;
      57854:data<=16'd1932;
      57855:data<=16'd2986;
      57856:data<=16'd3777;
      57857:data<=16'd3469;
      57858:data<=-16'd1107;
      57859:data<=-16'd2346;
      57860:data<=-16'd62;
      57861:data<=-16'd2687;
      57862:data<=16'd980;
      57863:data<=16'd12751;
      57864:data<=16'd15540;
      57865:data<=16'd12886;
      57866:data<=16'd13248;
      57867:data<=16'd12935;
      57868:data<=16'd13444;
      57869:data<=16'd14149;
      57870:data<=16'd12490;
      57871:data<=16'd11699;
      57872:data<=16'd11317;
      57873:data<=16'd10314;
      57874:data<=16'd10128;
      57875:data<=16'd10188;
      57876:data<=16'd10073;
      57877:data<=16'd9242;
      57878:data<=16'd8589;
      57879:data<=16'd9482;
      57880:data<=16'd10369;
      57881:data<=16'd10763;
      57882:data<=16'd10393;
      57883:data<=16'd8959;
      57884:data<=16'd8097;
      57885:data<=16'd7582;
      57886:data<=16'd7391;
      57887:data<=16'd7518;
      57888:data<=16'd6604;
      57889:data<=16'd6234;
      57890:data<=16'd6144;
      57891:data<=16'd5403;
      57892:data<=16'd6399;
      57893:data<=16'd7553;
      57894:data<=16'd8081;
      57895:data<=16'd7758;
      57896:data<=16'd995;
      57897:data<=-16'd8131;
      57898:data<=-16'd10147;
      57899:data<=-16'd7382;
      57900:data<=-16'd4316;
      57901:data<=-16'd2591;
      57902:data<=-16'd3260;
      57903:data<=-16'd3659;
      57904:data<=-16'd2802;
      57905:data<=-16'd1550;
      57906:data<=-16'd240;
      57907:data<=-16'd578;
      57908:data<=-16'd1604;
      57909:data<=-16'd1582;
      57910:data<=-16'd1415;
      57911:data<=-16'd1330;
      57912:data<=-16'd1477;
      57913:data<=-16'd1967;
      57914:data<=-16'd2105;
      57915:data<=-16'd1830;
      57916:data<=-16'd1727;
      57917:data<=-16'd1503;
      57918:data<=16'd288;
      57919:data<=16'd1378;
      57920:data<=16'd59;
      57921:data<=16'd171;
      57922:data<=16'd194;
      57923:data<=-16'd1234;
      57924:data<=-16'd347;
      57925:data<=-16'd582;
      57926:data<=-16'd1234;
      57927:data<=16'd284;
      57928:data<=-16'd1733;
      57929:data<=16'd1280;
      57930:data<=16'd13476;
      57931:data<=16'd17367;
      57932:data<=16'd14319;
      57933:data<=16'd14807;
      57934:data<=16'd13629;
      57935:data<=16'd11624;
      57936:data<=16'd11394;
      57937:data<=16'd10657;
      57938:data<=16'd10446;
      57939:data<=16'd9690;
      57940:data<=16'd9329;
      57941:data<=16'd8690;
      57942:data<=16'd5413;
      57943:data<=16'd5301;
      57944:data<=16'd6660;
      57945:data<=16'd4922;
      57946:data<=16'd5212;
      57947:data<=16'd5655;
      57948:data<=16'd4316;
      57949:data<=16'd4596;
      57950:data<=16'd3803;
      57951:data<=16'd2608;
      57952:data<=16'd2705;
      57953:data<=16'd2067;
      57954:data<=16'd2268;
      57955:data<=16'd3010;
      57956:data<=16'd3533;
      57957:data<=16'd3993;
      57958:data<=16'd3245;
      57959:data<=16'd2972;
      57960:data<=16'd2187;
      57961:data<=16'd1821;
      57962:data<=16'd2651;
      57963:data<=-16'd4147;
      57964:data<=-16'd13590;
      57965:data<=-16'd13863;
      57966:data<=-16'd12463;
      57967:data<=-16'd12427;
      57968:data<=-16'd9567;
      57969:data<=-16'd8573;
      57970:data<=-16'd9159;
      57971:data<=-16'd8543;
      57972:data<=-16'd8181;
      57973:data<=-16'd8094;
      57974:data<=-16'd8777;
      57975:data<=-16'd9051;
      57976:data<=-16'd8279;
      57977:data<=-16'd7846;
      57978:data<=-16'd7263;
      57979:data<=-16'd7350;
      57980:data<=-16'd6801;
      57981:data<=-16'd4931;
      57982:data<=-16'd5187;
      57983:data<=-16'd4613;
      57984:data<=-16'd1216;
      57985:data<=16'd312;
      57986:data<=-16'd287;
      57987:data<=-16'd798;
      57988:data<=-16'd738;
      57989:data<=-16'd1215;
      57990:data<=-16'd1753;
      57991:data<=-16'd719;
      57992:data<=-16'd1545;
      57993:data<=-16'd2176;
      57994:data<=-16'd681;
      57995:data<=-16'd3253;
      57996:data<=-16'd563;
      57997:data<=16'd11309;
      57998:data<=16'd14213;
      57999:data<=16'd10916;
      58000:data<=16'd12172;
      58001:data<=16'd11282;
      58002:data<=16'd9559;
      58003:data<=16'd9676;
      58004:data<=16'd8379;
      58005:data<=16'd7594;
      58006:data<=16'd6213;
      58007:data<=16'd4693;
      58008:data<=16'd5087;
      58009:data<=16'd4746;
      58010:data<=16'd4532;
      58011:data<=16'd4153;
      58012:data<=16'd3310;
      58013:data<=16'd4118;
      58014:data<=16'd3300;
      58015:data<=16'd2055;
      58016:data<=16'd2981;
      58017:data<=16'd1942;
      58018:data<=16'd2;
      58019:data<=-16'd772;
      58020:data<=-16'd1213;
      58021:data<=-16'd819;
      58022:data<=-16'd1309;
      58023:data<=-16'd1630;
      58024:data<=-16'd860;
      58025:data<=-16'd2055;
      58026:data<=-16'd4552;
      58027:data<=-16'd6428;
      58028:data<=-16'd5457;
      58029:data<=-16'd4781;
      58030:data<=-16'd12677;
      58031:data<=-16'd21611;
      58032:data<=-16'd21996;
      58033:data<=-16'd20641;
      58034:data<=-16'd20034;
      58035:data<=-16'd18171;
      58036:data<=-16'd17688;
      58037:data<=-16'd17471;
      58038:data<=-16'd16311;
      58039:data<=-16'd15415;
      58040:data<=-16'd15097;
      58041:data<=-16'd15317;
      58042:data<=-16'd15314;
      58043:data<=-16'd15579;
      58044:data<=-16'd15828;
      58045:data<=-16'd15218;
      58046:data<=-16'd14847;
      58047:data<=-16'd14078;
      58048:data<=-16'd13103;
      58049:data<=-16'd12750;
      58050:data<=-16'd12178;
      58051:data<=-16'd12108;
      58052:data<=-16'd11309;
      58053:data<=-16'd9817;
      58054:data<=-16'd10009;
      58055:data<=-16'd10160;
      58056:data<=-16'd10945;
      58057:data<=-16'd11768;
      58058:data<=-16'd10020;
      58059:data<=-16'd9967;
      58060:data<=-16'd9696;
      58061:data<=-16'd7932;
      58062:data<=-16'd10141;
      58063:data<=-16'd6376;
      58064:data<=16'd5395;
      58065:data<=16'd8439;
      58066:data<=16'd5882;
      58067:data<=16'd7509;
      58068:data<=16'd8381;
      58069:data<=16'd7756;
      58070:data<=16'd7658;
      58071:data<=16'd7004;
      58072:data<=16'd6692;
      58073:data<=16'd6925;
      58074:data<=16'd7151;
      58075:data<=16'd6986;
      58076:data<=16'd6687;
      58077:data<=16'd6267;
      58078:data<=16'd5439;
      58079:data<=16'd5627;
      58080:data<=16'd5131;
      58081:data<=16'd3024;
      58082:data<=16'd2773;
      58083:data<=16'd3353;
      58084:data<=16'd3242;
      58085:data<=16'd3018;
      58086:data<=16'd2111;
      58087:data<=16'd2347;
      58088:data<=16'd2497;
      58089:data<=16'd1604;
      58090:data<=16'd2523;
      58091:data<=16'd2607;
      58092:data<=16'd1720;
      58093:data<=16'd1278;
      58094:data<=-16'd1158;
      58095:data<=-16'd805;
      58096:data<=-16'd155;
      58097:data<=-16'd7920;
      58098:data<=-16'd14895;
      58099:data<=-16'd14624;
      58100:data<=-16'd13869;
      58101:data<=-16'd13201;
      58102:data<=-16'd11838;
      58103:data<=-16'd11086;
      58104:data<=-16'd10705;
      58105:data<=-16'd11135;
      58106:data<=-16'd11524;
      58107:data<=-16'd11708;
      58108:data<=-16'd11552;
      58109:data<=-16'd11447;
      58110:data<=-16'd13200;
      58111:data<=-16'd13820;
      58112:data<=-16'd12825;
      58113:data<=-16'd13083;
      58114:data<=-16'd12292;
      58115:data<=-16'd11003;
      58116:data<=-16'd10595;
      58117:data<=-16'd10135;
      58118:data<=-16'd11192;
      58119:data<=-16'd11141;
      58120:data<=-16'd9814;
      58121:data<=-16'd10278;
      58122:data<=-16'd9054;
      58123:data<=-16'd7988;
      58124:data<=-16'd8774;
      58125:data<=-16'd7309;
      58126:data<=-16'd7048;
      58127:data<=-16'd6880;
      58128:data<=-16'd5221;
      58129:data<=-16'd7529;
      58130:data<=-16'd4349;
      58131:data<=16'd6587;
      58132:data<=16'd8994;
      58133:data<=16'd6401;
      58134:data<=16'd7877;
      58135:data<=16'd7574;
      58136:data<=16'd6476;
      58137:data<=16'd7063;
      58138:data<=16'd6196;
      58139:data<=16'd5759;
      58140:data<=16'd6617;
      58141:data<=16'd6617;
      58142:data<=16'd5905;
      58143:data<=16'd4830;
      58144:data<=16'd3676;
      58145:data<=16'd3339;
      58146:data<=16'd3832;
      58147:data<=16'd3911;
      58148:data<=16'd3706;
      58149:data<=16'd4052;
      58150:data<=16'd3886;
      58151:data<=16'd4194;
      58152:data<=16'd6105;
      58153:data<=16'd7491;
      58154:data<=16'd7932;
      58155:data<=16'd7101;
      58156:data<=16'd5156;
      58157:data<=16'd4636;
      58158:data<=16'd4563;
      58159:data<=16'd4655;
      58160:data<=16'd5371;
      58161:data<=16'd4405;
      58162:data<=16'd4702;
      58163:data<=16'd4328;
      58164:data<=-16'd3886;
      58165:data<=-16'd11030;
      58166:data<=-16'd10031;
      58167:data<=-16'd9561;
      58168:data<=-16'd10742;
      58169:data<=-16'd10134;
      58170:data<=-16'd9859;
      58171:data<=-16'd9423;
      58172:data<=-16'd8622;
      58173:data<=-16'd8184;
      58174:data<=-16'd7316;
      58175:data<=-16'd7019;
      58176:data<=-16'd7018;
      58177:data<=-16'd6398;
      58178:data<=-16'd5791;
      58179:data<=-16'd5269;
      58180:data<=-16'd5623;
      58181:data<=-16'd6508;
      58182:data<=-16'd6422;
      58183:data<=-16'd5924;
      58184:data<=-16'd5497;
      58185:data<=-16'd5009;
      58186:data<=-16'd4262;
      58187:data<=-16'd3653;
      58188:data<=-16'd3820;
      58189:data<=-16'd3353;
      58190:data<=-16'd2987;
      58191:data<=-16'd3354;
      58192:data<=-16'd2353;
      58193:data<=-16'd2717;
      58194:data<=-16'd4531;
      58195:data<=-16'd5056;
      58196:data<=-16'd6813;
      58197:data<=-16'd3110;
      58198:data<=16'd8601;
      58199:data<=16'd12477;
      58200:data<=16'd9171;
      58201:data<=16'd10107;
      58202:data<=16'd10255;
      58203:data<=16'd8789;
      58204:data<=16'd9229;
      58205:data<=16'd8581;
      58206:data<=16'd9188;
      58207:data<=16'd10728;
      58208:data<=16'd9661;
      58209:data<=16'd9200;
      58210:data<=16'd9549;
      58211:data<=16'd9353;
      58212:data<=16'd9700;
      58213:data<=16'd9075;
      58214:data<=16'd8461;
      58215:data<=16'd9198;
      58216:data<=16'd9048;
      58217:data<=16'd8331;
      58218:data<=16'd8399;
      58219:data<=16'd8765;
      58220:data<=16'd9016;
      58221:data<=16'd8930;
      58222:data<=16'd8598;
      58223:data<=16'd8355;
      58224:data<=16'd8390;
      58225:data<=16'd8257;
      58226:data<=16'd7911;
      58227:data<=16'd7482;
      58228:data<=16'd6586;
      58229:data<=16'd6881;
      58230:data<=16'd5959;
      58231:data<=-16'd1163;
      58232:data<=-16'd7338;
      58233:data<=-16'd6602;
      58234:data<=-16'd6026;
      58235:data<=-16'd6231;
      58236:data<=-16'd3166;
      58237:data<=-16'd435;
      58238:data<=-16'd70;
      58239:data<=-16'd5;
      58240:data<=16'd635;
      58241:data<=16'd746;
      58242:data<=16'd23;
      58243:data<=16'd775;
      58244:data<=16'd2132;
      58245:data<=16'd2235;
      58246:data<=16'd2557;
      58247:data<=16'd2532;
      58248:data<=16'd2029;
      58249:data<=16'd2353;
      58250:data<=16'd2514;
      58251:data<=16'd2502;
      58252:data<=16'd2731;
      58253:data<=16'd2937;
      58254:data<=16'd2930;
      58255:data<=16'd2948;
      58256:data<=16'd4228;
      58257:data<=16'd4516;
      58258:data<=16'd3647;
      58259:data<=16'd4755;
      58260:data<=16'd4698;
      58261:data<=16'd4593;
      58262:data<=16'd5900;
      58263:data<=16'd3207;
      58264:data<=16'd6128;
      58265:data<=16'd18254;
      58266:data<=16'd21039;
      58267:data<=16'd16797;
      58268:data<=16'd18315;
      58269:data<=16'd19052;
      58270:data<=16'd17443;
      58271:data<=16'd17271;
      58272:data<=16'd15922;
      58273:data<=16'd14715;
      58274:data<=16'd14697;
      58275:data<=16'd14134;
      58276:data<=16'd13532;
      58277:data<=16'd13019;
      58278:data<=16'd11359;
      58279:data<=16'd8402;
      58280:data<=16'd7401;
      58281:data<=16'd8668;
      58282:data<=16'd8492;
      58283:data<=16'd8146;
      58284:data<=16'd8317;
      58285:data<=16'd7136;
      58286:data<=16'd6449;
      58287:data<=16'd6546;
      58288:data<=16'd6288;
      58289:data<=16'd6031;
      58290:data<=16'd6040;
      58291:data<=16'd6099;
      58292:data<=16'd5048;
      58293:data<=16'd5389;
      58294:data<=16'd7279;
      58295:data<=16'd6484;
      58296:data<=16'd6531;
      58297:data<=16'd4958;
      58298:data<=-16'd4704;
      58299:data<=-16'd11145;
      58300:data<=-16'd9693;
      58301:data<=-16'd9474;
      58302:data<=-16'd9564;
      58303:data<=-16'd8681;
      58304:data<=-16'd8645;
      58305:data<=-16'd7821;
      58306:data<=-16'd6640;
      58307:data<=-16'd5098;
      58308:data<=-16'd4678;
      58309:data<=-16'd5650;
      58310:data<=-16'd5131;
      58311:data<=-16'd5365;
      58312:data<=-16'd5606;
      58313:data<=-16'd4320;
      58314:data<=-16'd4814;
      58315:data<=-16'd4690;
      58316:data<=-16'd4100;
      58317:data<=-16'd4842;
      58318:data<=-16'd3571;
      58319:data<=-16'd2529;
      58320:data<=-16'd896;
      58321:data<=16'd2667;
      58322:data<=16'd2552;
      58323:data<=16'd1867;
      58324:data<=16'd2193;
      58325:data<=16'd1131;
      58326:data<=16'd2190;
      58327:data<=16'd2080;
      58328:data<=16'd1480;
      58329:data<=16'd2637;
      58330:data<=-16'd126;
      58331:data<=16'd4053;
      58332:data<=16'd17082;
      58333:data<=16'd19179;
      58334:data<=16'd15470;
      58335:data<=16'd16469;
      58336:data<=16'd15091;
      58337:data<=16'd13668;
      58338:data<=16'd14178;
      58339:data<=16'd12619;
      58340:data<=16'd11602;
      58341:data<=16'd11314;
      58342:data<=16'd10469;
      58343:data<=16'd10325;
      58344:data<=16'd10906;
      58345:data<=16'd11307;
      58346:data<=16'd10449;
      58347:data<=16'd9761;
      58348:data<=16'd9268;
      58349:data<=16'd7999;
      58350:data<=16'd8134;
      58351:data<=16'd8011;
      58352:data<=16'd6490;
      58353:data<=16'd5847;
      58354:data<=16'd5150;
      58355:data<=16'd5034;
      58356:data<=16'd5583;
      58357:data<=16'd5730;
      58358:data<=16'd6338;
      58359:data<=16'd5338;
      58360:data<=16'd4854;
      58361:data<=16'd5629;
      58362:data<=16'd2449;
      58363:data<=16'd117;
      58364:data<=-16'd2080;
      58365:data<=-16'd11371;
      58366:data<=-16'd17520;
      58367:data<=-16'd16145;
      58368:data<=-16'd15317;
      58369:data<=-16'd13944;
      58370:data<=-16'd12377;
      58371:data<=-16'd12565;
      58372:data<=-16'd12217;
      58373:data<=-16'd12028;
      58374:data<=-16'd11509;
      58375:data<=-16'd10924;
      58376:data<=-16'd11279;
      58377:data<=-16'd10837;
      58378:data<=-16'd10721;
      58379:data<=-16'd10666;
      58380:data<=-16'd9964;
      58381:data<=-16'd9717;
      58382:data<=-16'd8012;
      58383:data<=-16'd6828;
      58384:data<=-16'd7441;
      58385:data<=-16'd6869;
      58386:data<=-16'd7050;
      58387:data<=-16'd7269;
      58388:data<=-16'd6346;
      58389:data<=-16'd6799;
      58390:data<=-16'd6282;
      58391:data<=-16'd5967;
      58392:data<=-16'd6828;
      58393:data<=-16'd5538;
      58394:data<=-16'd5745;
      58395:data<=-16'd5956;
      58396:data<=-16'd4766;
      58397:data<=-16'd7286;
      58398:data<=-16'd3046;
      58399:data<=16'd8953;
      58400:data<=16'd10771;
      58401:data<=16'd7694;
      58402:data<=16'd9069;
      58403:data<=16'd7548;
      58404:data<=16'd7235;
      58405:data<=16'd11057;
      58406:data<=16'd10210;
      58407:data<=16'd7356;
      58408:data<=16'd7585;
      58409:data<=16'd7139;
      58410:data<=16'd6173;
      58411:data<=16'd6284;
      58412:data<=16'd5292;
      58413:data<=16'd4391;
      58414:data<=16'd4817;
      58415:data<=16'd4017;
      58416:data<=16'd3057;
      58417:data<=16'd3615;
      58418:data<=16'd3074;
      58419:data<=16'd1066;
      58420:data<=-16'd631;
      58421:data<=-16'd936;
      58422:data<=-16'd47;
      58423:data<=-16'd318;
      58424:data<=-16'd785;
      58425:data<=-16'd411;
      58426:data<=-16'd1068;
      58427:data<=-16'd863;
      58428:data<=-16'd872;
      58429:data<=-16'd2085;
      58430:data<=-16'd140;
      58431:data<=-16'd2834;
      58432:data<=-16'd14628;
      58433:data<=-16'd20266;
      58434:data<=-16'd17954;
      58435:data<=-16'd17860;
      58436:data<=-16'd17411;
      58437:data<=-16'd15869;
      58438:data<=-16'd15861;
      58439:data<=-16'd14904;
      58440:data<=-16'd14357;
      58441:data<=-16'd14606;
      58442:data<=-16'd13436;
      58443:data<=-16'd13444;
      58444:data<=-16'd14615;
      58445:data<=-16'd14233;
      58446:data<=-16'd14791;
      58447:data<=-16'd17441;
      58448:data<=-16'd17961;
      58449:data<=-16'd16157;
      58450:data<=-16'd15782;
      58451:data<=-16'd15459;
      58452:data<=-16'd14013;
      58453:data<=-16'd13844;
      58454:data<=-16'd13256;
      58455:data<=-16'd12102;
      58456:data<=-16'd12944;
      58457:data<=-16'd13330;
      58458:data<=-16'd12883;
      58459:data<=-16'd12689;
      58460:data<=-16'd11523;
      58461:data<=-16'd11265;
      58462:data<=-16'd10449;
      58463:data<=-16'd9091;
      58464:data<=-16'd11042;
      58465:data<=-16'd6877;
      58466:data<=16'd5103;
      58467:data<=16'd8237;
      58468:data<=16'd4678;
      58469:data<=16'd4792;
      58470:data<=16'd3980;
      58471:data<=16'd3159;
      58472:data<=16'd4208;
      58473:data<=16'd3002;
      58474:data<=16'd2655;
      58475:data<=16'd3307;
      58476:data<=16'd2341;
      58477:data<=16'd2828;
      58478:data<=16'd3068;
      58479:data<=16'd2190;
      58480:data<=16'd2996;
      58481:data<=16'd2376;
      58482:data<=16'd564;
      58483:data<=16'd675;
      58484:data<=16'd347;
      58485:data<=16'd229;
      58486:data<=16'd893;
      58487:data<=-16'd329;
      58488:data<=16'd555;
      58489:data<=16'd4667;
      58490:data<=16'd5398;
      58491:data<=16'd4203;
      58492:data<=16'd4663;
      58493:data<=16'd3794;
      58494:data<=16'd2508;
      58495:data<=16'd1765;
      58496:data<=16'd916;
      58497:data<=16'd2582;
      58498:data<=16'd317;
      58499:data<=-16'd9791;
      58500:data<=-16'd14973;
      58501:data<=-16'd13101;
      58502:data<=-16'd12757;
      58503:data<=-16'd12345;
      58504:data<=-16'd11371;
      58505:data<=-16'd11127;
      58506:data<=-16'd10237;
      58507:data<=-16'd11030;
      58508:data<=-16'd11808;
      58509:data<=-16'd10546;
      58510:data<=-16'd10194;
      58511:data<=-16'd9740;
      58512:data<=-16'd9074;
      58513:data<=-16'd9127;
      58514:data<=-16'd8129;
      58515:data<=-16'd7611;
      58516:data<=-16'd7542;
      58517:data<=-16'd6384;
      58518:data<=-16'd5653;
      58519:data<=-16'd5808;
      58520:data<=-16'd6787;
      58521:data<=-16'd7071;
      58522:data<=-16'd6273;
      58523:data<=-16'd6166;
      58524:data<=-16'd5142;
      58525:data<=-16'd4831;
      58526:data<=-16'd5627;
      58527:data<=-16'd4208;
      58528:data<=-16'd4162;
      58529:data<=-16'd3550;
      58530:data<=-16'd2504;
      58531:data<=-16'd8246;
      58532:data<=-16'd6623;
      58533:data<=16'd6106;
      58534:data<=16'd8525;
      58535:data<=16'd5653;
      58536:data<=16'd7794;
      58537:data<=16'd6734;
      58538:data<=16'd6162;
      58539:data<=16'd7674;
      58540:data<=16'd6311;
      58541:data<=16'd6156;
      58542:data<=16'd6566;
      58543:data<=16'd6310;
      58544:data<=16'd6341;
      58545:data<=16'd4482;
      58546:data<=16'd4093;
      58547:data<=16'd5016;
      58548:data<=16'd3883;
      58549:data<=16'd3686;
      58550:data<=16'd3839;
      58551:data<=16'd3233;
      58552:data<=16'd3647;
      58553:data<=16'd3465;
      58554:data<=16'd2951;
      58555:data<=16'd3559;
      58556:data<=16'd3454;
      58557:data<=16'd1707;
      58558:data<=16'd958;
      58559:data<=16'd1798;
      58560:data<=16'd1231;
      58561:data<=16'd1158;
      58562:data<=16'd1701;
      58563:data<=16'd520;
      58564:data<=16'd2143;
      58565:data<=16'd196;
      58566:data<=-16'd10477;
      58567:data<=-16'd14442;
      58568:data<=-16'd11926;
      58569:data<=-16'd13221;
      58570:data<=-16'd13211;
      58571:data<=-16'd12812;
      58572:data<=-16'd12075;
      58573:data<=-16'd7524;
      58574:data<=-16'd6068;
      58575:data<=-16'd6088;
      58576:data<=-16'd4388;
      58577:data<=-16'd4936;
      58578:data<=-16'd4901;
      58579:data<=-16'd4425;
      58580:data<=-16'd4457;
      58581:data<=-16'd3833;
      58582:data<=-16'd5586;
      58583:data<=-16'd6059;
      58584:data<=-16'd4291;
      58585:data<=-16'd4196;
      58586:data<=-16'd3286;
      58587:data<=-16'd3245;
      58588:data<=-16'd3870;
      58589:data<=-16'd2543;
      58590:data<=-16'd2364;
      58591:data<=-16'd1303;
      58592:data<=-16'd707;
      58593:data<=-16'd2117;
      58594:data<=-16'd711;
      58595:data<=-16'd673;
      58596:data<=-16'd505;
      58597:data<=16'd1383;
      58598:data<=-16'd1691;
      58599:data<=16'd3021;
      58600:data<=16'd15976;
      58601:data<=16'd17303;
      58602:data<=16'd14575;
      58603:data<=16'd15719;
      58604:data<=16'd14287;
      58605:data<=16'd14364;
      58606:data<=16'd14794;
      58607:data<=16'd13838;
      58608:data<=16'd14868;
      58609:data<=16'd14428;
      58610:data<=16'd13741;
      58611:data<=16'd13570;
      58612:data<=16'd12389;
      58613:data<=16'd13374;
      58614:data<=16'd12407;
      58615:data<=16'd8548;
      58616:data<=16'd7764;
      58617:data<=16'd7641;
      58618:data<=16'd6473;
      58619:data<=16'd6878;
      58620:data<=16'd8487;
      58621:data<=16'd8931;
      58622:data<=16'd7874;
      58623:data<=16'd8003;
      58624:data<=16'd7706;
      58625:data<=16'd6772;
      58626:data<=16'd7632;
      58627:data<=16'd6869;
      58628:data<=16'd6736;
      58629:data<=16'd7653;
      58630:data<=16'd5463;
      58631:data<=16'd6884;
      58632:data<=16'd6058;
      58633:data<=-16'd4407;
      58634:data<=-16'd8519;
      58635:data<=-16'd6109;
      58636:data<=-16'd7274;
      58637:data<=-16'd6849;
      58638:data<=-16'd6197;
      58639:data<=-16'd6278;
      58640:data<=-16'd4918;
      58641:data<=-16'd5497;
      58642:data<=-16'd4907;
      58643:data<=-16'd4055;
      58644:data<=-16'd4651;
      58645:data<=-16'd2214;
      58646:data<=-16'd1472;
      58647:data<=-16'd2531;
      58648:data<=-16'd1306;
      58649:data<=-16'd1936;
      58650:data<=-16'd2087;
      58651:data<=-16'd776;
      58652:data<=-16'd910;
      58653:data<=16'd182;
      58654:data<=16'd227;
      58655:data<=-16'd917;
      58656:data<=16'd957;
      58657:data<=16'd4572;
      58658:data<=16'd7464;
      58659:data<=16'd6675;
      58660:data<=16'd5685;
      58661:data<=16'd7321;
      58662:data<=16'd5667;
      58663:data<=16'd5541;
      58664:data<=16'd7251;
      58665:data<=16'd3997;
      58666:data<=16'd8768;
      58667:data<=16'd20219;
      58668:data<=16'd20894;
      58669:data<=16'd18841;
      58670:data<=16'd20409;
      58671:data<=16'd19079;
      58672:data<=16'd18360;
      58673:data<=16'd18615;
      58674:data<=16'd17136;
      58675:data<=16'd16468;
      58676:data<=16'd16169;
      58677:data<=16'd15336;
      58678:data<=16'd14528;
      58679:data<=16'd14016;
      58680:data<=16'd13823;
      58681:data<=16'd13455;
      58682:data<=16'd13712;
      58683:data<=16'd14079;
      58684:data<=16'd13515;
      58685:data<=16'd12656;
      58686:data<=16'd11776;
      58687:data<=16'd11417;
      58688:data<=16'd10869;
      58689:data<=16'd9994;
      58690:data<=16'd9585;
      58691:data<=16'd8617;
      58692:data<=16'd8680;
      58693:data<=16'd8819;
      58694:data<=16'd7480;
      58695:data<=16'd9030;
      58696:data<=16'd9667;
      58697:data<=16'd7633;
      58698:data<=16'd8470;
      58699:data<=16'd2764;
      58700:data<=-16'd9644;
      58701:data<=-16'd13007;
      58702:data<=-16'd11761;
      58703:data<=-16'd12913;
      58704:data<=-16'd11870;
      58705:data<=-16'd10959;
      58706:data<=-16'd10856;
      58707:data<=-16'd9294;
      58708:data<=-16'd7952;
      58709:data<=-16'd7219;
      58710:data<=-16'd7451;
      58711:data<=-16'd7535;
      58712:data<=-16'd6927;
      58713:data<=-16'd7100;
      58714:data<=-16'd6946;
      58715:data<=-16'd7060;
      58716:data<=-16'd7128;
      58717:data<=-16'd6276;
      58718:data<=-16'd6828;
      58719:data<=-16'd5993;
      58720:data<=-16'd3483;
      58721:data<=-16'd3360;
      58722:data<=-16'd3265;
      58723:data<=-16'd3198;
      58724:data<=-16'd3357;
      58725:data<=-16'd2246;
      58726:data<=-16'd3463;
      58727:data<=-16'd4094;
      58728:data<=-16'd2710;
      58729:data<=-16'd3718;
      58730:data<=-16'd2846;
      58731:data<=-16'd2287;
      58732:data<=-16'd3751;
      58733:data<=16'd4109;
      58734:data<=16'd14566;
      58735:data<=16'd14850;
      58736:data<=16'd12815;
      58737:data<=16'd12989;
      58738:data<=16'd12252;
      58739:data<=16'd11576;
      58740:data<=16'd11671;
      58741:data<=16'd13273;
      58742:data<=16'd14371;
      58743:data<=16'd13135;
      58744:data<=16'd12901;
      58745:data<=16'd13621;
      58746:data<=16'd13165;
      58747:data<=16'd12706;
      58748:data<=16'd12609;
      58749:data<=16'd11809;
      58750:data<=16'd10308;
      58751:data<=16'd9592;
      58752:data<=16'd9298;
      58753:data<=16'd8266;
      58754:data<=16'd7806;
      58755:data<=16'd7163;
      58756:data<=16'd6097;
      58757:data<=16'd6570;
      58758:data<=16'd6855;
      58759:data<=16'd6799;
      58760:data<=16'd7109;
      58761:data<=16'd6108;
      58762:data<=16'd5658;
      58763:data<=16'd5042;
      58764:data<=16'd3791;
      58765:data<=16'd5303;
      58766:data<=16'd2005;
      58767:data<=-16'd8733;
      58768:data<=-16'd13170;
      58769:data<=-16'd10830;
      58770:data<=-16'd10278;
      58771:data<=-16'd9643;
      58772:data<=-16'd8786;
      58773:data<=-16'd9028;
      58774:data<=-16'd8354;
      58775:data<=-16'd8046;
      58776:data<=-16'd8434;
      58777:data<=-16'd8320;
      58778:data<=-16'd8160;
      58779:data<=-16'd7771;
      58780:data<=-16'd7881;
      58781:data<=-16'd8408;
      58782:data<=-16'd8296;
      58783:data<=-16'd8901;
      58784:data<=-16'd9908;
      58785:data<=-16'd9746;
      58786:data<=-16'd9338;
      58787:data<=-16'd8983;
      58788:data<=-16'd8366;
      58789:data<=-16'd8354;
      58790:data<=-16'd8784;
      58791:data<=-16'd8072;
      58792:data<=-16'd6919;
      58793:data<=-16'd7520;
      58794:data<=-16'd7905;
      58795:data<=-16'd6984;
      58796:data<=-16'd7006;
      58797:data<=-16'd6294;
      58798:data<=-16'd5974;
      58799:data<=-16'd6975;
      58800:data<=-16'd808;
      58801:data<=16'd8752;
      58802:data<=16'd9373;
      58803:data<=16'd7174;
      58804:data<=16'd7718;
      58805:data<=16'd6449;
      58806:data<=16'd5932;
      58807:data<=16'd6125;
      58808:data<=16'd4035;
      58809:data<=16'd3075;
      58810:data<=16'd2978;
      58811:data<=16'd2325;
      58812:data<=16'd2315;
      58813:data<=16'd1542;
      58814:data<=16'd1166;
      58815:data<=16'd2264;
      58816:data<=16'd2053;
      58817:data<=16'd987;
      58818:data<=16'd728;
      58819:data<=16'd318;
      58820:data<=-16'd757;
      58821:data<=-16'd1657;
      58822:data<=-16'd2008;
      58823:data<=-16'd2532;
      58824:data<=-16'd2296;
      58825:data<=-16'd161;
      58826:data<=16'd1651;
      58827:data<=16'd1603;
      58828:data<=16'd1168;
      58829:data<=16'd931;
      58830:data<=-16'd356;
      58831:data<=-16'd793;
      58832:data<=16'd658;
      58833:data<=-16'd4200;
      58834:data<=-16'd15235;
      58835:data<=-16'd18803;
      58836:data<=-16'd16372;
      58837:data<=-16'd16835;
      58838:data<=-16'd16659;
      58839:data<=-16'd15558;
      58840:data<=-16'd15508;
      58841:data<=-16'd14327;
      58842:data<=-16'd14023;
      58843:data<=-16'd13999;
      58844:data<=-16'd12860;
      58845:data<=-16'd13359;
      58846:data<=-16'd13943;
      58847:data<=-16'd13640;
      58848:data<=-16'd13838;
      58849:data<=-16'd13462;
      58850:data<=-16'd12892;
      58851:data<=-16'd12336;
      58852:data<=-16'd11597;
      58853:data<=-16'd11210;
      58854:data<=-16'd10622;
      58855:data<=-16'd10278;
      58856:data<=-16'd9661;
      58857:data<=-16'd9320;
      58858:data<=-16'd10552;
      58859:data<=-16'd10213;
      58860:data<=-16'd9274;
      58861:data<=-16'd9966;
      58862:data<=-16'd9377;
      58863:data<=-16'd8619;
      58864:data<=-16'd7973;
      58865:data<=-16'd7171;
      58866:data<=-16'd7758;
      58867:data<=-16'd3412;
      58868:data<=16'd3971;
      58869:data<=16'd4481;
      58870:data<=16'd2491;
      58871:data<=16'd1920;
      58872:data<=16'd896;
      58873:data<=16'd1456;
      58874:data<=16'd1703;
      58875:data<=16'd1386;
      58876:data<=16'd2038;
      58877:data<=16'd1400;
      58878:data<=16'd1218;
      58879:data<=16'd1348;
      58880:data<=16'd575;
      58881:data<=16'd1694;
      58882:data<=16'd1994;
      58883:data<=16'd50;
      58884:data<=-16'd688;
      58885:data<=-16'd781;
      58886:data<=-16'd1031;
      58887:data<=-16'd1262;
      58888:data<=-16'd1149;
      58889:data<=-16'd785;
      58890:data<=-16'd1424;
      58891:data<=-16'd1400;
      58892:data<=-16'd1312;
      58893:data<=-16'd2080;
      58894:data<=-16'd1221;
      58895:data<=-16'd1709;
      58896:data<=-16'd3776;
      58897:data<=-16'd3803;
      58898:data<=-16'd3497;
      58899:data<=-16'd2350;
      58900:data<=-16'd4690;
      58901:data<=-16'd13863;
      58902:data<=-16'd17429;
      58903:data<=-16'd14187;
      58904:data<=-16'd14246;
      58905:data<=-16'd14396;
      58906:data<=-16'd12869;
      58907:data<=-16'd13100;
      58908:data<=-16'd13330;
      58909:data<=-16'd11721;
      58910:data<=-16'd8505;
      58911:data<=-16'd7127;
      58912:data<=-16'd7803;
      58913:data<=-16'd6757;
      58914:data<=-16'd6514;
      58915:data<=-16'd7289;
      58916:data<=-16'd6141;
      58917:data<=-16'd5823;
      58918:data<=-16'd6162;
      58919:data<=-16'd5265;
      58920:data<=-16'd5197;
      58921:data<=-16'd6260;
      58922:data<=-16'd6435;
      58923:data<=-16'd5277;
      58924:data<=-16'd4972;
      58925:data<=-16'd4836;
      58926:data<=-16'd3342;
      58927:data<=-16'd3383;
      58928:data<=-16'd3372;
      58929:data<=-16'd2120;
      58930:data<=-16'd2494;
      58931:data<=-16'd1770;
      58932:data<=-16'd2059;
      58933:data<=-16'd3817;
      58934:data<=16'd2349;
      58935:data<=16'd10386;
      58936:data<=16'd10628;
      58937:data<=16'd9643;
      58938:data<=16'd9805;
      58939:data<=16'd9124;
      58940:data<=16'd9080;
      58941:data<=16'd9206;
      58942:data<=16'd9230;
      58943:data<=16'd8728;
      58944:data<=16'd8634;
      58945:data<=16'd8458;
      58946:data<=16'd6028;
      58947:data<=16'd5641;
      58948:data<=16'd6816;
      58949:data<=16'd5902;
      58950:data<=16'd6152;
      58951:data<=16'd4752;
      58952:data<=16'd1239;
      58953:data<=16'd1257;
      58954:data<=16'd1492;
      58955:data<=16'd1318;
      58956:data<=16'd2114;
      58957:data<=16'd811;
      58958:data<=-16'd209;
      58959:data<=-16'd801;
      58960:data<=-16'd1404;
      58961:data<=-16'd232;
      58962:data<=-16'd476;
      58963:data<=-16'd229;
      58964:data<=16'd705;
      58965:data<=-16'd332;
      58966:data<=16'd1343;
      58967:data<=-16'd1051;
      58968:data<=-16'd10646;
      58969:data<=-16'd12848;
      58970:data<=-16'd10681;
      58971:data<=-16'd12690;
      58972:data<=-16'd12696;
      58973:data<=-16'd11482;
      58974:data<=-16'd11306;
      58975:data<=-16'd10293;
      58976:data<=-16'd9970;
      58977:data<=-16'd9277;
      58978:data<=-16'd8414;
      58979:data<=-16'd8241;
      58980:data<=-16'd7342;
      58981:data<=-16'd7342;
      58982:data<=-16'd7830;
      58983:data<=-16'd7832;
      58984:data<=-16'd8287;
      58985:data<=-16'd7921;
      58986:data<=-16'd7282;
      58987:data<=-16'd6590;
      58988:data<=-16'd5418;
      58989:data<=-16'd5127;
      58990:data<=-16'd4250;
      58991:data<=-16'd3448;
      58992:data<=-16'd3468;
      58993:data<=-16'd779;
      58994:data<=16'd2457;
      58995:data<=16'd2955;
      58996:data<=16'd2475;
      58997:data<=16'd2516;
      58998:data<=16'd3342;
      58999:data<=16'd2601;
      59000:data<=16'd3212;
      59001:data<=16'd10803;
      59002:data<=16'd17244;
      59003:data<=16'd16628;
      59004:data<=16'd15797;
      59005:data<=16'd15893;
      59006:data<=16'd14956;
      59007:data<=16'd14915;
      59008:data<=16'd15802;
      59009:data<=16'd16468;
      59010:data<=16'd16064;
      59011:data<=16'd15429;
      59012:data<=16'd15352;
      59013:data<=16'd14919;
      59014:data<=16'd14960;
      59015:data<=16'd14968;
      59016:data<=16'd14176;
      59017:data<=16'd14176;
      59018:data<=16'd13808;
      59019:data<=16'd12989;
      59020:data<=16'd13443;
      59021:data<=16'd13835;
      59022:data<=16'd13796;
      59023:data<=16'd13361;
      59024:data<=16'd12612;
      59025:data<=16'd12605;
      59026:data<=16'd11969;
      59027:data<=16'd11257;
      59028:data<=16'd11458;
      59029:data<=16'd10919;
      59030:data<=16'd10921;
      59031:data<=16'd10560;
      59032:data<=16'd9442;
      59033:data<=16'd11415;
      59034:data<=16'd9492;
      59035:data<=-16'd1193;
      59036:data<=-16'd7632;
      59037:data<=-16'd5958;
      59038:data<=-16'd5553;
      59039:data<=-16'd6243;
      59040:data<=-16'd5319;
      59041:data<=-16'd5166;
      59042:data<=-16'd5069;
      59043:data<=-16'd4470;
      59044:data<=-16'd4687;
      59045:data<=-16'd3958;
      59046:data<=-16'd1918;
      59047:data<=-16'd1190;
      59048:data<=-16'd1721;
      59049:data<=-16'd2099;
      59050:data<=-16'd2005;
      59051:data<=-16'd1738;
      59052:data<=-16'd2030;
      59053:data<=-16'd1873;
      59054:data<=-16'd860;
      59055:data<=-16'd617;
      59056:data<=-16'd466;
      59057:data<=16'd5;
      59058:data<=16'd437;
      59059:data<=16'd1973;
      59060:data<=16'd2740;
      59061:data<=16'd2080;
      59062:data<=16'd2309;
      59063:data<=16'd2000;
      59064:data<=16'd1720;
      59065:data<=16'd2490;
      59066:data<=16'd1275;
      59067:data<=16'd2487;
      59068:data<=16'd9893;
      59069:data<=16'd15026;
      59070:data<=16'd14939;
      59071:data<=16'd15303;
      59072:data<=16'd15864;
      59073:data<=16'd14869;
      59074:data<=16'd14543;
      59075:data<=16'd14533;
      59076:data<=16'd13223;
      59077:data<=16'd13628;
      59078:data<=16'd16381;
      59079:data<=16'd16753;
      59080:data<=16'd15571;
      59081:data<=16'd15625;
      59082:data<=16'd14792;
      59083:data<=16'd14534;
      59084:data<=16'd15857;
      59085:data<=16'd15227;
      59086:data<=16'd14122;
      59087:data<=16'd13808;
      59088:data<=16'd12272;
      59089:data<=16'd11253;
      59090:data<=16'd10925;
      59091:data<=16'd9975;
      59092:data<=16'd9647;
      59093:data<=16'd9333;
      59094:data<=16'd8837;
      59095:data<=16'd9168;
      59096:data<=16'd10100;
      59097:data<=16'd11062;
      59098:data<=16'd9806;
      59099:data<=16'd8572;
      59100:data<=16'd10202;
      59101:data<=16'd6150;
      59102:data<=-16'd4053;
      59103:data<=-16'd7336;
      59104:data<=-16'd5066;
      59105:data<=-16'd5277;
      59106:data<=-16'd5480;
      59107:data<=-16'd5177;
      59108:data<=-16'd4952;
      59109:data<=-16'd2811;
      59110:data<=-16'd1927;
      59111:data<=-16'd3234;
      59112:data<=-16'd3380;
      59113:data<=-16'd3069;
      59114:data<=-16'd3090;
      59115:data<=-16'd3084;
      59116:data<=-16'd4079;
      59117:data<=-16'd4391;
      59118:data<=-16'd3521;
      59119:data<=-16'd5109;
      59120:data<=-16'd7612;
      59121:data<=-16'd6579;
      59122:data<=-16'd4567;
      59123:data<=-16'd4379;
      59124:data<=-16'd4305;
      59125:data<=-16'd4317;
      59126:data<=-16'd4375;
      59127:data<=-16'd3855;
      59128:data<=-16'd4099;
      59129:data<=-16'd4608;
      59130:data<=-16'd4502;
      59131:data<=-16'd4299;
      59132:data<=-16'd4147;
      59133:data<=-16'd4299;
      59134:data<=-16'd1071;
      59135:data<=16'd6962;
      59136:data<=16'd11785;
      59137:data<=16'd11157;
      59138:data<=16'd10323;
      59139:data<=16'd9600;
      59140:data<=16'd8965;
      59141:data<=16'd9021;
      59142:data<=16'd8393;
      59143:data<=16'd7370;
      59144:data<=16'd6293;
      59145:data<=16'd6313;
      59146:data<=16'd7805;
      59147:data<=16'd8147;
      59148:data<=16'd7583;
      59149:data<=16'd7191;
      59150:data<=16'd6724;
      59151:data<=16'd6657;
      59152:data<=16'd6075;
      59153:data<=16'd5526;
      59154:data<=16'd5325;
      59155:data<=16'd4149;
      59156:data<=16'd3427;
      59157:data<=16'd2749;
      59158:data<=16'd2546;
      59159:data<=16'd3965;
      59160:data<=16'd3398;
      59161:data<=16'd4159;
      59162:data<=16'd7949;
      59163:data<=16'd7612;
      59164:data<=16'd6437;
      59165:data<=16'd6398;
      59166:data<=16'd4676;
      59167:data<=16'd5987;
      59168:data<=16'd2834;
      59169:data<=-16'd7973;
      59170:data<=-16'd10343;
      59171:data<=-16'd6601;
      59172:data<=-16'd6799;
      59173:data<=-16'd6752;
      59174:data<=-16'd6819;
      59175:data<=-16'd7329;
      59176:data<=-16'd6357;
      59177:data<=-16'd6302;
      59178:data<=-16'd6276;
      59179:data<=-16'd6772;
      59180:data<=-16'd7480;
      59181:data<=-16'd6432;
      59182:data<=-16'd7081;
      59183:data<=-16'd7492;
      59184:data<=-16'd5462;
      59185:data<=-16'd5339;
      59186:data<=-16'd5595;
      59187:data<=-16'd4998;
      59188:data<=-16'd5200;
      59189:data<=-16'd4746;
      59190:data<=-16'd4443;
      59191:data<=-16'd4420;
      59192:data<=-16'd4167;
      59193:data<=-16'd4219;
      59194:data<=-16'd3442;
      59195:data<=-16'd3626;
      59196:data<=-16'd4666;
      59197:data<=-16'd4325;
      59198:data<=-16'd4091;
      59199:data<=-16'd3814;
      59200:data<=-16'd4664;
      59201:data<=-16'd3941;
      59202:data<=16'd4073;
      59203:data<=16'd8716;
      59204:data<=16'd4405;
      59205:data<=16'd2801;
      59206:data<=16'd3541;
      59207:data<=16'd2370;
      59208:data<=16'd2120;
      59209:data<=16'd1061;
      59210:data<=-16'd183;
      59211:data<=-16'd385;
      59212:data<=-16'd1005;
      59213:data<=-16'd537;
      59214:data<=-16'd443;
      59215:data<=-16'd1210;
      59216:data<=-16'd729;
      59217:data<=-16'd649;
      59218:data<=-16'd600;
      59219:data<=-16'd214;
      59220:data<=-16'd1257;
      59221:data<=-16'd2786;
      59222:data<=-16'd4026;
      59223:data<=-16'd4309;
      59224:data<=-16'd4217;
      59225:data<=-16'd5025;
      59226:data<=-16'd5289;
      59227:data<=-16'd5589;
      59228:data<=-16'd5495;
      59229:data<=-16'd4222;
      59230:data<=-16'd4572;
      59231:data<=-16'd4692;
      59232:data<=-16'd4581;
      59233:data<=-16'd6097;
      59234:data<=-16'd5641;
      59235:data<=-16'd9295;
      59236:data<=-16'd19077;
      59237:data<=-16'd21460;
      59238:data<=-16'd18512;
      59239:data<=-16'd18936;
      59240:data<=-16'd18553;
      59241:data<=-16'd17699;
      59242:data<=-16'd17523;
      59243:data<=-16'd16095;
      59244:data<=-16'd15694;
      59245:data<=-16'd14222;
      59246:data<=-16'd11459;
      59247:data<=-16'd11658;
      59248:data<=-16'd11884;
      59249:data<=-16'd10963;
      59250:data<=-16'd11715;
      59251:data<=-16'd12060;
      59252:data<=-16'd11421;
      59253:data<=-16'd11220;
      59254:data<=-16'd10413;
      59255:data<=-16'd9661;
      59256:data<=-16'd9424;
      59257:data<=-16'd8475;
      59258:data<=-16'd8501;
      59259:data<=-16'd9861;
      59260:data<=-16'd9709;
      59261:data<=-16'd8974;
      59262:data<=-16'd9042;
      59263:data<=-16'd8810;
      59264:data<=-16'd8863;
      59265:data<=-16'd8040;
      59266:data<=-16'd6834;
      59267:data<=-16'd8219;
      59268:data<=-16'd5981;
      59269:data<=16'd2823;
      59270:data<=16'd7837;
      59271:data<=16'd6241;
      59272:data<=16'd4306;
      59273:data<=16'd3786;
      59274:data<=16'd3829;
      59275:data<=16'd3607;
      59276:data<=16'd3432;
      59277:data<=16'd3500;
      59278:data<=16'd2843;
      59279:data<=16'd2552;
      59280:data<=16'd2502;
      59281:data<=16'd2149;
      59282:data<=16'd2825;
      59283:data<=16'd2808;
      59284:data<=16'd1339;
      59285:data<=16'd823;
      59286:data<=16'd1231;
      59287:data<=16'd97;
      59288:data<=-16'd3654;
      59289:data<=-16'd5422;
      59290:data<=-16'd3623;
      59291:data<=-16'd3824;
      59292:data<=-16'd4451;
      59293:data<=-16'd3568;
      59294:data<=-16'd4262;
      59295:data<=-16'd3512;
      59296:data<=-16'd3315;
      59297:data<=-16'd6378;
      59298:data<=-16'd6096;
      59299:data<=-16'd5369;
      59300:data<=-16'd6134;
      59301:data<=-16'd3594;
      59302:data<=-16'd6940;
      59303:data<=-16'd16471;
      59304:data<=-16'd18346;
      59305:data<=-16'd16049;
      59306:data<=-16'd16264;
      59307:data<=-16'd15646;
      59308:data<=-16'd14998;
      59309:data<=-16'd15223;
      59310:data<=-16'd14947;
      59311:data<=-16'd14505;
      59312:data<=-16'd13890;
      59313:data<=-16'd13530;
      59314:data<=-16'd12839;
      59315:data<=-16'd11650;
      59316:data<=-16'd11621;
      59317:data<=-16'd11787;
      59318:data<=-16'd11141;
      59319:data<=-16'd10351;
      59320:data<=-16'd9471;
      59321:data<=-16'd9495;
      59322:data<=-16'd10241;
      59323:data<=-16'd9831;
      59324:data<=-16'd8898;
      59325:data<=-16'd8781;
      59326:data<=-16'd8358;
      59327:data<=-16'd7407;
      59328:data<=-16'd7322;
      59329:data<=-16'd6005;
      59330:data<=-16'd2643;
      59331:data<=-16'd1322;
      59332:data<=-16'd798;
      59333:data<=16'd56;
      59334:data<=-16'd2481;
      59335:data<=-16'd1362;
      59336:data<=16'd7741;
      59337:data<=16'd12499;
      59338:data<=16'd10837;
      59339:data<=16'd11095;
      59340:data<=16'd11426;
      59341:data<=16'd10199;
      59342:data<=16'd9961;
      59343:data<=16'd9993;
      59344:data<=16'd10276;
      59345:data<=16'd10369;
      59346:data<=16'd8974;
      59347:data<=16'd7533;
      59348:data<=16'd7133;
      59349:data<=16'd7415;
      59350:data<=16'd7761;
      59351:data<=16'd7682;
      59352:data<=16'd7747;
      59353:data<=16'd8025;
      59354:data<=16'd7658;
      59355:data<=16'd6693;
      59356:data<=16'd6443;
      59357:data<=16'd6869;
      59358:data<=16'd6152;
      59359:data<=16'd5095;
      59360:data<=16'd4672;
      59361:data<=16'd3896;
      59362:data<=16'd4071;
      59363:data<=16'd4408;
      59364:data<=16'd3425;
      59365:data<=16'd3683;
      59366:data<=16'd3689;
      59367:data<=16'd3445;
      59368:data<=16'd5321;
      59369:data<=16'd1688;
      59370:data<=-16'd7415;
      59371:data<=-16'd11414;
      59372:data<=-16'd12956;
      59373:data<=-16'd15120;
      59374:data<=-16'd14093;
      59375:data<=-16'd13077;
      59376:data<=-16'd12707;
      59377:data<=-16'd11060;
      59378:data<=-16'd10543;
      59379:data<=-16'd10037;
      59380:data<=-16'd9132;
      59381:data<=-16'd8828;
      59382:data<=-16'd7814;
      59383:data<=-16'd7961;
      59384:data<=-16'd9125;
      59385:data<=-16'd9003;
      59386:data<=-16'd8843;
      59387:data<=-16'd8282;
      59388:data<=-16'd7289;
      59389:data<=-16'd6805;
      59390:data<=-16'd5579;
      59391:data<=-16'd4869;
      59392:data<=-16'd5095;
      59393:data<=-16'd4281;
      59394:data<=-16'd3648;
      59395:data<=-16'd3761;
      59396:data<=-16'd3096;
      59397:data<=-16'd2308;
      59398:data<=-16'd2455;
      59399:data<=-16'd1818;
      59400:data<=-16'd623;
      59401:data<=-16'd1701;
      59402:data<=16'd848;
      59403:data<=16'd10366;
      59404:data<=16'd14751;
      59405:data<=16'd12449;
      59406:data<=16'd12801;
      59407:data<=16'd13124;
      59408:data<=16'd12158;
      59409:data<=16'd13080;
      59410:data<=16'd13655;
      59411:data<=16'd13620;
      59412:data<=16'd12742;
      59413:data<=16'd12508;
      59414:data<=16'd15479;
      59415:data<=16'd16897;
      59416:data<=16'd16267;
      59417:data<=16'd16393;
      59418:data<=16'd15458;
      59419:data<=16'd15282;
      59420:data<=16'd15719;
      59421:data<=16'd15226;
      59422:data<=16'd16004;
      59423:data<=16'd16075;
      59424:data<=16'd15406;
      59425:data<=16'd15420;
      59426:data<=16'd14258;
      59427:data<=16'd13850;
      59428:data<=16'd13673;
      59429:data<=16'd12689;
      59430:data<=16'd12886;
      59431:data<=16'd12193;
      59432:data<=16'd11796;
      59433:data<=16'd11803;
      59434:data<=16'd11162;
      59435:data<=16'd13696;
      59436:data<=16'd10439;
      59437:data<=-16'd557;
      59438:data<=-16'd2707;
      59439:data<=-16'd92;
      59440:data<=-16'd1324;
      59441:data<=-16'd414;
      59442:data<=-16'd358;
      59443:data<=-16'd1104;
      59444:data<=16'd540;
      59445:data<=16'd2;
      59446:data<=16'd253;
      59447:data<=16'd2102;
      59448:data<=16'd2093;
      59449:data<=16'd2587;
      59450:data<=16'd2196;
      59451:data<=16'd1612;
      59452:data<=16'd2264;
      59453:data<=16'd1283;
      59454:data<=16'd1744;
      59455:data<=16'd2061;
      59456:data<=-16'd1272;
      59457:data<=-16'd2513;
      59458:data<=-16'd1883;
      59459:data<=-16'd1486;
      59460:data<=16'd684;
      59461:data<=16'd1569;
      59462:data<=16'd943;
      59463:data<=16'd1309;
      59464:data<=16'd1289;
      59465:data<=16'd860;
      59466:data<=16'd1392;
      59467:data<=16'd1905;
      59468:data<=16'd898;
      59469:data<=16'd3447;
      59470:data<=16'd11979;
      59471:data<=16'd16211;
      59472:data<=16'd14935;
      59473:data<=16'd15659;
      59474:data<=16'd15388;
      59475:data<=16'd13749;
      59476:data<=16'd13743;
      59477:data<=16'd13347;
      59478:data<=16'd13230;
      59479:data<=16'd12581;
      59480:data<=16'd11115;
      59481:data<=16'd11414;
      59482:data<=16'd11086;
      59483:data<=16'd10170;
      59484:data<=16'd10830;
      59485:data<=16'd11740;
      59486:data<=16'd12640;
      59487:data<=16'd12457;
      59488:data<=16'd11449;
      59489:data<=16'd10749;
      59490:data<=16'd9491;
      59491:data<=16'd9289;
      59492:data<=16'd9050;
      59493:data<=16'd7823;
      59494:data<=16'd7917;
      59495:data<=16'd6872;
      59496:data<=16'd6325;
      59497:data<=16'd9006;
      59498:data<=16'd11051;
      59499:data<=16'd12657;
      59500:data<=16'd12380;
      59501:data<=16'd10807;
      59502:data<=16'd12325;
      59503:data<=16'd7787;
      59504:data<=-16'd2593;
      59505:data<=-16'd4614;
      59506:data<=-16'd2519;
      59507:data<=-16'd3136;
      59508:data<=-16'd3148;
      59509:data<=-16'd2737;
      59510:data<=-16'd1554;
      59511:data<=-16'd663;
      59512:data<=-16'd1060;
      59513:data<=-16'd628;
      59514:data<=-16'd945;
      59515:data<=-16'd1095;
      59516:data<=-16'd375;
      59517:data<=-16'd1474;
      59518:data<=-16'd2159;
      59519:data<=-16'd2326;
      59520:data<=-16'd3116;
      59521:data<=-16'd2276;
      59522:data<=-16'd996;
      59523:data<=-16'd138;
      59524:data<=16'd358;
      59525:data<=16'd229;
      59526:data<=16'd591;
      59527:data<=16'd102;
      59528:data<=-16'd306;
      59529:data<=16'd268;
      59530:data<=-16'd86;
      59531:data<=16'd265;
      59532:data<=-16'd179;
      59533:data<=-16'd1277;
      59534:data<=16'd218;
      59535:data<=16'd400;
      59536:data<=16'd3401;
      59537:data<=16'd12398;
      59538:data<=16'd15376;
      59539:data<=16'd12595;
      59540:data<=16'd10777;
      59541:data<=16'd8132;
      59542:data<=16'd7247;
      59543:data<=16'd7292;
      59544:data<=16'd6018;
      59545:data<=16'd5915;
      59546:data<=16'd5095;
      59547:data<=16'd5134;
      59548:data<=16'd6799;
      59549:data<=16'd6131;
      59550:data<=16'd5830;
      59551:data<=16'd6006;
      59552:data<=16'd5197;
      59553:data<=16'd5747;
      59554:data<=16'd5447;
      59555:data<=16'd4587;
      59556:data<=16'd4269;
      59557:data<=16'd2890;
      59558:data<=16'd2607;
      59559:data<=16'd2670;
      59560:data<=16'd3068;
      59561:data<=16'd4552;
      59562:data<=16'd3248;
      59563:data<=16'd2322;
      59564:data<=16'd3046;
      59565:data<=16'd1721;
      59566:data<=16'd1839;
      59567:data<=16'd1791;
      59568:data<=16'd889;
      59569:data<=16'd2399;
      59570:data<=-16'd2094;
      59571:data<=-16'd10460;
      59572:data<=-16'd10684;
      59573:data<=-16'd8147;
      59574:data<=-16'd8395;
      59575:data<=-16'd8207;
      59576:data<=-16'd7908;
      59577:data<=-16'd8056;
      59578:data<=-16'd8184;
      59579:data<=-16'd7671;
      59580:data<=-16'd7271;
      59581:data<=-16'd7773;
      59582:data<=-16'd6657;
      59583:data<=-16'd5225;
      59584:data<=-16'd5106;
      59585:data<=-16'd4131;
      59586:data<=-16'd3657;
      59587:data<=-16'd4065;
      59588:data<=-16'd3923;
      59589:data<=-16'd3861;
      59590:data<=-16'd3668;
      59591:data<=-16'd3862;
      59592:data<=-16'd3732;
      59593:data<=-16'd3057;
      59594:data<=-16'd3838;
      59595:data<=-16'd4027;
      59596:data<=-16'd3723;
      59597:data<=-16'd4096;
      59598:data<=-16'd3101;
      59599:data<=-16'd3391;
      59600:data<=-16'd4085;
      59601:data<=-16'd3444;
      59602:data<=-16'd5110;
      59603:data<=-16'd1958;
      59604:data<=16'd7480;
      59605:data<=16'd10157;
      59606:data<=16'd7899;
      59607:data<=16'd7946;
      59608:data<=16'd7697;
      59609:data<=16'd6557;
      59610:data<=16'd4716;
      59611:data<=16'd3591;
      59612:data<=16'd4026;
      59613:data<=16'd3013;
      59614:data<=16'd2344;
      59615:data<=16'd2604;
      59616:data<=16'd1674;
      59617:data<=16'd1774;
      59618:data<=16'd2064;
      59619:data<=16'd1525;
      59620:data<=16'd1733;
      59621:data<=16'd1397;
      59622:data<=16'd646;
      59623:data<=-16'd820;
      59624:data<=-16'd3485;
      59625:data<=-16'd4899;
      59626:data<=-16'd5342;
      59627:data<=-16'd4915;
      59628:data<=-16'd4364;
      59629:data<=-16'd5686;
      59630:data<=-16'd5447;
      59631:data<=-16'd4496;
      59632:data<=-16'd5626;
      59633:data<=-16'd5213;
      59634:data<=-16'd5598;
      59635:data<=-16'd7353;
      59636:data<=-16'd6722;
      59637:data<=-16'd11044;
      59638:data<=-16'd19634;
      59639:data<=-16'd20983;
      59640:data<=-16'd18726;
      59641:data<=-16'd18941;
      59642:data<=-16'd18272;
      59643:data<=-16'd17400;
      59644:data<=-16'd17575;
      59645:data<=-16'd16586;
      59646:data<=-16'd15437;
      59647:data<=-16'd16099;
      59648:data<=-16'd17371;
      59649:data<=-16'd17262;
      59650:data<=-16'd16368;
      59651:data<=-16'd15993;
      59652:data<=-16'd15716;
      59653:data<=-16'd15488;
      59654:data<=-16'd15400;
      59655:data<=-16'd14775;
      59656:data<=-16'd13951;
      59657:data<=-16'd13268;
      59658:data<=-16'd12308;
      59659:data<=-16'd11750;
      59660:data<=-16'd12417;
      59661:data<=-16'd13071;
      59662:data<=-16'd12842;
      59663:data<=-16'd12604;
      59664:data<=-16'd11896;
      59665:data<=-16'd10922;
      59666:data<=-16'd10505;
      59667:data<=-16'd8493;
      59668:data<=-16'd7262;
      59669:data<=-16'd9226;
      59670:data<=-16'd5256;
      59671:data<=16'd4672;
      59672:data<=16'd6830;
      59673:data<=16'd3318;
      59674:data<=16'd3538;
      59675:data<=16'd3941;
      59676:data<=16'd2898;
      59677:data<=16'd3121;
      59678:data<=16'd2863;
      59679:data<=16'd2203;
      59680:data<=16'd2256;
      59681:data<=16'd2105;
      59682:data<=16'd2235;
      59683:data<=16'd2751;
      59684:data<=16'd2519;
      59685:data<=16'd1368;
      59686:data<=16'd459;
      59687:data<=16'd567;
      59688:data<=16'd635;
      59689:data<=16'd452;
      59690:data<=16'd470;
      59691:data<=16'd111;
      59692:data<=-16'd187;
      59693:data<=-16'd321;
      59694:data<=-16'd525;
      59695:data<=-16'd79;
      59696:data<=16'd32;
      59697:data<=-16'd957;
      59698:data<=-16'd2391;
      59699:data<=-16'd3345;
      59700:data<=-16'd2831;
      59701:data<=-16'd2748;
      59702:data<=-16'd2911;
      59703:data<=-16'd2009;
      59704:data<=-16'd6197;
      59705:data<=-16'd14211;
      59706:data<=-16'd15618;
      59707:data<=-16'd13292;
      59708:data<=-16'd13837;
      59709:data<=-16'd14871;
      59710:data<=-16'd15788;
      59711:data<=-16'd16201;
      59712:data<=-16'd14959;
      59713:data<=-16'd14207;
      59714:data<=-16'd14004;
      59715:data<=-16'd13594;
      59716:data<=-16'd13317;
      59717:data<=-16'd12425;
      59718:data<=-16'd11609;
      59719:data<=-16'd11447;
      59720:data<=-16'd10736;
      59721:data<=-16'd9747;
      59722:data<=-16'd10138;
      59723:data<=-16'd11420;
      59724:data<=-16'd11183;
      59725:data<=-16'd9964;
      59726:data<=-16'd9468;
      59727:data<=-16'd8998;
      59728:data<=-16'd8575;
      59729:data<=-16'd8313;
      59730:data<=-16'd7838;
      59731:data<=-16'd7077;
      59732:data<=-16'd5739;
      59733:data<=-16'd5385;
      59734:data<=-16'd5280;
      59735:data<=-16'd5150;
      59736:data<=-16'd7398;
      59737:data<=-16'd4244;
      59738:data<=16'd5909;
      59739:data<=16'd8802;
      59740:data<=16'd6593;
      59741:data<=16'd8041;
      59742:data<=16'd7700;
      59743:data<=16'd6666;
      59744:data<=16'd7847;
      59745:data<=16'd7764;
      59746:data<=16'd7501;
      59747:data<=16'd6335;
      59748:data<=16'd4370;
      59749:data<=16'd4581;
      59750:data<=16'd5365;
      59751:data<=16'd6836;
      59752:data<=16'd7850;
      59753:data<=16'd6857;
      59754:data<=16'd7459;
      59755:data<=16'd8120;
      59756:data<=16'd7426;
      59757:data<=16'd7718;
      59758:data<=16'd7350;
      59759:data<=16'd6728;
      59760:data<=16'd5830;
      59761:data<=16'd4240;
      59762:data<=16'd4828;
      59763:data<=16'd5025;
      59764:data<=16'd4270;
      59765:data<=16'd4786;
      59766:data<=16'd3982;
      59767:data<=16'd3862;
      59768:data<=16'd4752;
      59769:data<=16'd4402;
      59770:data<=16'd4576;
      59771:data<=-16'd177;
      59772:data<=-16'd8742;
      59773:data<=-16'd10516;
      59774:data<=-16'd9219;
      59775:data<=-16'd9292;
      59776:data<=-16'd8099;
      59777:data<=-16'd7712;
      59778:data<=-16'd7559;
      59779:data<=-16'd6598;
      59780:data<=-16'd5964;
      59781:data<=-16'd5048;
      59782:data<=-16'd5034;
      59783:data<=-16'd4764;
      59784:data<=-16'd3987;
      59785:data<=-16'd5298;
      59786:data<=-16'd6211;
      59787:data<=-16'd5788;
      59788:data<=-16'd5507;
      59789:data<=-16'd5095;
      59790:data<=-16'd4978;
      59791:data<=-16'd3751;
      59792:data<=-16'd3074;
      59793:data<=-16'd4817;
      59794:data<=-16'd4924;
      59795:data<=-16'd4115;
      59796:data<=-16'd4206;
      59797:data<=-16'd3557;
      59798:data<=-16'd3046;
      59799:data<=-16'd2372;
      59800:data<=-16'd2173;
      59801:data<=-16'd1858;
      59802:data<=-16'd635;
      59803:data<=-16'd2223;
      59804:data<=16'd989;
      59805:data<=16'd11626;
      59806:data<=16'd14137;
      59807:data<=16'd11365;
      59808:data<=16'd12853;
      59809:data<=16'd12427;
      59810:data<=16'd12269;
      59811:data<=16'd14290;
      59812:data<=16'd13503;
      59813:data<=16'd12928;
      59814:data<=16'd12760;
      59815:data<=16'd11861;
      59816:data<=16'd12201;
      59817:data<=16'd11988;
      59818:data<=16'd11861;
      59819:data<=16'd11994;
      59820:data<=16'd11241;
      59821:data<=16'd11447;
      59822:data<=16'd11884;
      59823:data<=16'd12631;
      59824:data<=16'd13327;
      59825:data<=16'd12110;
      59826:data<=16'd11715;
      59827:data<=16'd11826;
      59828:data<=16'd11253;
      59829:data<=16'd11635;
      59830:data<=16'd10977;
      59831:data<=16'd10354;
      59832:data<=16'd10683;
      59833:data<=16'd9624;
      59834:data<=16'd9796;
      59835:data<=16'd11505;
      59836:data<=16'd13274;
      59837:data<=16'd13341;
      59838:data<=16'd6684;
      59839:data<=-16'd641;
      59840:data<=-16'd1115;
      59841:data<=-16'd246;
      59842:data<=-16'd414;
      59843:data<=-16'd115;
      59844:data<=-16'd68;
      59845:data<=16'd138;
      59846:data<=16'd86;
      59847:data<=16'd992;
      59848:data<=16'd2605;
      59849:data<=16'd2731;
      59850:data<=16'd3071;
      59851:data<=16'd3289;
      59852:data<=16'd2798;
      59853:data<=16'd2772;
      59854:data<=16'd2293;
      59855:data<=16'd2667;
      59856:data<=16'd3096;
      59857:data<=16'd2406;
      59858:data<=16'd3106;
      59859:data<=16'd2964;
      59860:data<=16'd2726;
      59861:data<=16'd4915;
      59862:data<=16'd5184;
      59863:data<=16'd4504;
      59864:data<=16'd4663;
      59865:data<=16'd4322;
      59866:data<=16'd5066;
      59867:data<=16'd4552;
      59868:data<=16'd4366;
      59869:data<=16'd5551;
      59870:data<=16'd2795;
      59871:data<=16'd5457;
      59872:data<=16'd16169;
      59873:data<=16'd19132;
      59874:data<=16'd17054;
      59875:data<=16'd18001;
      59876:data<=16'd16883;
      59877:data<=16'd14551;
      59878:data<=16'd13591;
      59879:data<=16'd13168;
      59880:data<=16'd12775;
      59881:data<=16'd11527;
      59882:data<=16'd11348;
      59883:data<=16'd11079;
      59884:data<=16'd9624;
      59885:data<=16'd10419;
      59886:data<=16'd11618;
      59887:data<=16'd11505;
      59888:data<=16'd11312;
      59889:data<=16'd10433;
      59890:data<=16'd10154;
      59891:data<=16'd9734;
      59892:data<=16'd8504;
      59893:data<=16'd8378;
      59894:data<=16'd7905;
      59895:data<=16'd7467;
      59896:data<=16'd7357;
      59897:data<=16'd6590;
      59898:data<=16'd7765;
      59899:data<=16'd8728;
      59900:data<=16'd7952;
      59901:data<=16'd8069;
      59902:data<=16'd7112;
      59903:data<=16'd6831;
      59904:data<=16'd6570;
      59905:data<=-16'd185;
      59906:data<=-16'd6951;
      59907:data<=-16'd7351;
      59908:data<=-16'd6916;
      59909:data<=-16'd6981;
      59910:data<=-16'd5883;
      59911:data<=-16'd4469;
      59912:data<=-16'd3768;
      59913:data<=-16'd3950;
      59914:data<=-16'd3548;
      59915:data<=-16'd3327;
      59916:data<=-16'd3601;
      59917:data<=-16'd3277;
      59918:data<=-16'd3130;
      59919:data<=-16'd2002;
      59920:data<=-16'd1186;
      59921:data<=-16'd2370;
      59922:data<=-16'd1800;
      59923:data<=-16'd403;
      59924:data<=16'd118;
      59925:data<=16'd1113;
      59926:data<=16'd431;
      59927:data<=-16'd246;
      59928:data<=16'd438;
      59929:data<=16'd187;
      59930:data<=16'd531;
      59931:data<=16'd36;
      59932:data<=-16'd843;
      59933:data<=16'd373;
      59934:data<=-16'd466;
      59935:data<=-16'd211;
      59936:data<=16'd2206;
      59937:data<=16'd343;
      59938:data<=16'd3272;
      59939:data<=16'd12871;
      59940:data<=16'd14640;
      59941:data<=16'd11964;
      59942:data<=16'd12557;
      59943:data<=16'd12038;
      59944:data<=16'd10768;
      59945:data<=16'd10654;
      59946:data<=16'd10164;
      59947:data<=16'd9370;
      59948:data<=16'd9216;
      59949:data<=16'd9903;
      59950:data<=16'd9565;
      59951:data<=16'd8520;
      59952:data<=16'd8414;
      59953:data<=16'd7865;
      59954:data<=16'd7462;
      59955:data<=16'd7385;
      59956:data<=16'd6331;
      59957:data<=16'd6015;
      59958:data<=16'd5733;
      59959:data<=16'd4560;
      59960:data<=16'd4385;
      59961:data<=16'd4262;
      59962:data<=16'd3742;
      59963:data<=16'd3424;
      59964:data<=16'd2752;
      59965:data<=16'd2388;
      59966:data<=16'd2020;
      59967:data<=16'd1686;
      59968:data<=16'd1372;
      59969:data<=16'd277;
      59970:data<=16'd817;
      59971:data<=-16'd144;
      59972:data<=-16'd7347;
      59973:data<=-16'd12404;
      59974:data<=-16'd10889;
      59975:data<=-16'd10072;
      59976:data<=-16'd10621;
      59977:data<=-16'd10091;
      59978:data<=-16'd10013;
      59979:data<=-16'd9867;
      59980:data<=-16'd9192;
      59981:data<=-16'd8937;
      59982:data<=-16'd8748;
      59983:data<=-16'd8683;
      59984:data<=-16'd9174;
      59985:data<=-16'd8843;
      59986:data<=-16'd7131;
      59987:data<=-16'd6579;
      59988:data<=-16'd7288;
      59989:data<=-16'd6913;
      59990:data<=-16'd6560;
      59991:data<=-16'd6664;
      59992:data<=-16'd6285;
      59993:data<=-16'd6405;
      59994:data<=-16'd6144;
      59995:data<=-16'd5433;
      59996:data<=-16'd5624;
      59997:data<=-16'd5758;
      59998:data<=-16'd6314;
      59999:data<=-16'd6307;
      60000:data<=-16'd4954;
      60001:data<=-16'd5673;
      60002:data<=-16'd5418;
      60003:data<=-16'd3193;
      60004:data<=-16'd4349;
      60005:data<=-16'd1278;
      60006:data<=16'd8216;
      60007:data<=16'd10326;
      60008:data<=16'd7541;
      60009:data<=16'd8536;
      60010:data<=16'd7727;
      60011:data<=16'd4971;
      60012:data<=16'd4505;
      60013:data<=16'd4193;
      60014:data<=16'd3538;
      60015:data<=16'd2954;
      60016:data<=16'd2317;
      60017:data<=16'd2209;
      60018:data<=16'd1821;
      60019:data<=16'd1659;
      60020:data<=16'd1941;
      60021:data<=16'd1653;
      60022:data<=16'd1462;
      60023:data<=16'd640;
      60024:data<=-16'd1080;
      60025:data<=-16'd1541;
      60026:data<=-16'd1575;
      60027:data<=-16'd2522;
      60028:data<=-16'd2766;
      60029:data<=-16'd2320;
      60030:data<=-16'd2648;
      60031:data<=-16'd3008;
      60032:data<=-16'd2954;
      60033:data<=-16'd3240;
      60034:data<=-16'd3116;
      60035:data<=-16'd3644;
      60036:data<=-16'd5724;
      60037:data<=-16'd5782;
      60038:data<=-16'd6731;
      60039:data<=-16'd13671;
      60040:data<=-16'd18809;
      60041:data<=-16'd17798;
      60042:data<=-16'd17121;
      60043:data<=-16'd17212;
      60044:data<=-16'd16716;
      60045:data<=-16'd17500;
      60046:data<=-16'd17796;
      60047:data<=-16'd16724;
      60048:data<=-16'd16398;
      60049:data<=-16'd17249;
      60050:data<=-16'd17693;
      60051:data<=-16'd17145;
      60052:data<=-16'd16763;
      60053:data<=-16'd15902;
      60054:data<=-16'd15106;
      60055:data<=-16'd15858;
      60056:data<=-16'd15391;
      60057:data<=-16'd14087;
      60058:data<=-16'd13964;
      60059:data<=-16'd12953;
      60060:data<=-16'd12643;
      60061:data<=-16'd13693;
      60062:data<=-16'd13597;
      60063:data<=-16'd13485;
      60064:data<=-16'd13030;
      60065:data<=-16'd12387;
      60066:data<=-16'd12192;
      60067:data<=-16'd10872;
      60068:data<=-16'd10941;
      60069:data<=-16'd10850;
      60070:data<=-16'd9395;
      60071:data<=-16'd11047;
      60072:data<=-16'd7262;
      60073:data<=16'd2880;
      60074:data<=16'd3753;
      60075:data<=16'd705;
      60076:data<=16'd2532;
      60077:data<=16'd2111;
      60078:data<=16'd1340;
      60079:data<=16'd2200;
      60080:data<=16'd1313;
      60081:data<=16'd1319;
      60082:data<=16'd1234;
      60083:data<=16'd634;
      60084:data<=16'd1522;
      60085:data<=16'd1039;
      60086:data<=16'd253;
      60087:data<=16'd1004;
      60088:data<=16'd1389;
      60089:data<=16'd1553;
      60090:data<=16'd1216;
      60091:data<=16'd963;
      60092:data<=16'd1518;
      60093:data<=16'd1325;
      60094:data<=16'd981;
      60095:data<=16'd660;
      60096:data<=16'd341;
      60097:data<=16'd999;
      60098:data<=16'd535;
      60099:data<=-16'd1422;
      60100:data<=-16'd2332;
      60101:data<=-16'd1829;
      60102:data<=-16'd1697;
      60103:data<=-16'd2247;
      60104:data<=-16'd998;
      60105:data<=-16'd1968;
      60106:data<=-16'd9561;
      60107:data<=-16'd14677;
      60108:data<=-16'd13600;
      60109:data<=-16'd13164;
      60110:data<=-16'd12901;
      60111:data<=-16'd12483;
      60112:data<=-16'd13508;
      60113:data<=-16'd13000;
      60114:data<=-16'd11688;
      60115:data<=-16'd11241;
      60116:data<=-16'd10624;
      60117:data<=-16'd10225;
      60118:data<=-16'd10017;
      60119:data<=-16'd9811;
      60120:data<=-16'd9371;
      60121:data<=-16'd8878;
      60122:data<=-16'd8939;
      60123:data<=-16'd8677;
      60124:data<=-16'd9034;
      60125:data<=-16'd9644;
      60126:data<=-16'd8675;
      60127:data<=-16'd8191;
      60128:data<=-16'd7970;
      60129:data<=-16'd7732;
      60130:data<=-16'd8787;
      60131:data<=-16'd8366;
      60132:data<=-16'd7774;
      60133:data<=-16'd8061;
      60134:data<=-16'd6717;
      60135:data<=-16'd6975;
      60136:data<=-16'd7468;
      60137:data<=-16'd7045;
      60138:data<=-16'd9139;
      60139:data<=-16'd4880;
      60140:data<=16'd5418;
      60141:data<=16'd7729;
      60142:data<=16'd6170;
      60143:data<=16'd7095;
      60144:data<=16'd6396;
      60145:data<=16'd5648;
      60146:data<=16'd5832;
      60147:data<=16'd5644;
      60148:data<=16'd5181;
      60149:data<=16'd3771;
      60150:data<=16'd3501;
      60151:data<=16'd4034;
      60152:data<=16'd3556;
      60153:data<=16'd3755;
      60154:data<=16'd4058;
      60155:data<=16'd4114;
      60156:data<=16'd4308;
      60157:data<=16'd3776;
      60158:data<=16'd3805;
      60159:data<=16'd3991;
      60160:data<=16'd3468;
      60161:data<=16'd2638;
      60162:data<=16'd1101;
      60163:data<=16'd1058;
      60164:data<=16'd2132;
      60165:data<=16'd1979;
      60166:data<=16'd2102;
      60167:data<=16'd1997;
      60168:data<=16'd1983;
      60169:data<=16'd2403;
      60170:data<=16'd1900;
      60171:data<=16'd4037;
      60172:data<=16'd4056;
      60173:data<=-16'd4507;
      60174:data<=-16'd10604;
      60175:data<=-16'd9882;
      60176:data<=-16'd9521;
      60177:data<=-16'd8687;
      60178:data<=-16'd7588;
      60179:data<=-16'd7600;
      60180:data<=-16'd6766;
      60181:data<=-16'd6070;
      60182:data<=-16'd5339;
      60183:data<=-16'd4696;
      60184:data<=-16'd4836;
      60185:data<=-16'd4270;
      60186:data<=-16'd4670;
      60187:data<=-16'd5773;
      60188:data<=-16'd5342;
      60189:data<=-16'd4952;
      60190:data<=-16'd4605;
      60191:data<=-16'd4390;
      60192:data<=-16'd4516;
      60193:data<=-16'd3325;
      60194:data<=-16'd2317;
      60195:data<=-16'd1964;
      60196:data<=-16'd1524;
      60197:data<=-16'd1597;
      60198:data<=-16'd1155;
      60199:data<=-16'd1318;
      60200:data<=-16'd1465;
      60201:data<=-16'd140;
      60202:data<=-16'd570;
      60203:data<=-16'd124;
      60204:data<=16'd1275;
      60205:data<=-16'd911;
      60206:data<=16'd2740;
      60207:data<=16'd12912;
      60208:data<=16'd15150;
      60209:data<=16'd12610;
      60210:data<=16'd12901;
      60211:data<=16'd12975;
      60212:data<=16'd13455;
      60213:data<=16'd13494;
      60214:data<=16'd11543;
      60215:data<=16'd11068;
      60216:data<=16'd11306;
      60217:data<=16'd10854;
      60218:data<=16'd11050;
      60219:data<=16'd10859;
      60220:data<=16'd10222;
      60221:data<=16'd10163;
      60222:data<=16'd10154;
      60223:data<=16'd10126;
      60224:data<=16'd10695;
      60225:data<=16'd11662;
      60226:data<=16'd11815;
      60227:data<=16'd11101;
      60228:data<=16'd10439;
      60229:data<=16'd9859;
      60230:data<=16'd9676;
      60231:data<=16'd9894;
      60232:data<=16'd10075;
      60233:data<=16'd10099;
      60234:data<=16'd9492;
      60235:data<=16'd9147;
      60236:data<=16'd9639;
      60237:data<=16'd10593;
      60238:data<=16'd11958;
      60239:data<=16'd9270;
      60240:data<=16'd1378;
      60241:data<=-16'd3107;
      60242:data<=-16'd2400;
      60243:data<=-16'd2071;
      60244:data<=-16'd1891;
      60245:data<=-16'd1119;
      60246:data<=-16'd1022;
      60247:data<=-16'd1039;
      60248:data<=-16'd432;
      60249:data<=16'd1110;
      60250:data<=16'd2056;
      60251:data<=16'd1694;
      60252:data<=16'd1879;
      60253:data<=16'd1865;
      60254:data<=16'd1460;
      60255:data<=16'd2570;
      60256:data<=16'd3874;
      60257:data<=16'd4187;
      60258:data<=16'd4185;
      60259:data<=16'd3850;
      60260:data<=16'd3748;
      60261:data<=16'd4836;
      60262:data<=16'd6758;
      60263:data<=16'd7257;
      60264:data<=16'd6302;
      60265:data<=16'd6322;
      60266:data<=16'd5776;
      60267:data<=16'd4851;
      60268:data<=16'd5658;
      60269:data<=16'd5156;
      60270:data<=16'd4845;
      60271:data<=16'd5526;
      60272:data<=16'd3134;
      60273:data<=16'd6593;
      60274:data<=16'd17638;
      60275:data<=16'd20274;
      60276:data<=16'd17165;
      60277:data<=16'd18133;
      60278:data<=16'd17352;
      60279:data<=16'd15388;
      60280:data<=16'd15699;
      60281:data<=16'd14687;
      60282:data<=16'd13960;
      60283:data<=16'd14380;
      60284:data<=16'd13537;
      60285:data<=16'd12681;
      60286:data<=16'd12718;
      60287:data<=16'd13661;
      60288:data<=16'd14170;
      60289:data<=16'd12794;
      60290:data<=16'd11734;
      60291:data<=16'd11364;
      60292:data<=16'd10809;
      60293:data<=16'd10853;
      60294:data<=16'd10081;
      60295:data<=16'd8660;
      60296:data<=16'd8429;
      60297:data<=16'd7530;
      60298:data<=16'd5876;
      60299:data<=16'd6584;
      60300:data<=16'd8085;
      60301:data<=16'd7515;
      60302:data<=16'd7263;
      60303:data<=16'd7530;
      60304:data<=16'd6448;
      60305:data<=16'd6599;
      60306:data<=16'd4552;
      60307:data<=-16'd3442;
      60308:data<=-16'd7844;
      60309:data<=-16'd6608;
      60310:data<=-16'd7178;
      60311:data<=-16'd6575;
      60312:data<=-16'd3853;
      60313:data<=-16'd3600;
      60314:data<=-16'd3962;
      60315:data<=-16'd3821;
      60316:data<=-16'd3680;
      60317:data<=-16'd3306;
      60318:data<=-16'd3812;
      60319:data<=-16'd3991;
      60320:data<=-16'd3609;
      60321:data<=-16'd3550;
      60322:data<=-16'd3131;
      60323:data<=-16'd3130;
      60324:data<=-16'd2669;
      60325:data<=-16'd1475;
      60326:data<=-16'd1445;
      60327:data<=-16'd1219;
      60328:data<=-16'd745;
      60329:data<=-16'd911;
      60330:data<=-16'd943;
      60331:data<=-16'd1425;
      60332:data<=-16'd1300;
      60333:data<=-16'd963;
      60334:data<=-16'd1610;
      60335:data<=-16'd1322;
      60336:data<=-16'd913;
      60337:data<=16'd356;
      60338:data<=16'd1480;
      60339:data<=-16'd587;
      60340:data<=16'd4015;
      60341:data<=16'd14627;
      60342:data<=16'd15317;
      60343:data<=16'd11879;
      60344:data<=16'd12901;
      60345:data<=16'd11906;
      60346:data<=16'd11033;
      60347:data<=16'd11720;
      60348:data<=16'd10266;
      60349:data<=16'd9911;
      60350:data<=16'd10862;
      60351:data<=16'd10815;
      60352:data<=16'd10240;
      60353:data<=16'd9330;
      60354:data<=16'd9037;
      60355:data<=16'd8611;
      60356:data<=16'd7752;
      60357:data<=16'd7420;
      60358:data<=16'd6831;
      60359:data<=16'd6633;
      60360:data<=16'd6355;
      60361:data<=16'd5565;
      60362:data<=16'd5899;
      60363:data<=16'd5882;
      60364:data<=16'd5377;
      60365:data<=16'd5315;
      60366:data<=16'd4752;
      60367:data<=16'd4494;
      60368:data<=16'd3883;
      60369:data<=16'd3506;
      60370:data<=16'd3883;
      60371:data<=16'd3025;
      60372:data<=16'd3624;
      60373:data<=16'd1472;
      60374:data<=-16'd7125;
      60375:data<=-16'd9861;
      60376:data<=-16'd7354;
      60377:data<=-16'd8652;
      60378:data<=-16'd8367;
      60379:data<=-16'd7225;
      60380:data<=-16'd8070;
      60381:data<=-16'd8156;
      60382:data<=-16'd9787;
      60383:data<=-16'd9949;
      60384:data<=-16'd8381;
      60385:data<=-16'd9937;
      60386:data<=-16'd9527;
      60387:data<=-16'd7206;
      60388:data<=-16'd7081;
      60389:data<=-16'd6822;
      60390:data<=-16'd7181;
      60391:data<=-16'd7298;
      60392:data<=-16'd6648;
      60393:data<=-16'd7133;
      60394:data<=-16'd6237;
      60395:data<=-16'd5611;
      60396:data<=-16'd6194;
      60397:data<=-16'd5624;
      60398:data<=-16'd6024;
      60399:data<=-16'd5867;
      60400:data<=-16'd5291;
      60401:data<=-16'd6131;
      60402:data<=-16'd5359;
      60403:data<=-16'd5806;
      60404:data<=-16'd6375;
      60405:data<=-16'd5030;
      60406:data<=-16'd7359;
      60407:data<=-16'd4361;
      60408:data<=16'd5970;
      60409:data<=16'd7392;
      60410:data<=16'd4541;
      60411:data<=16'd5371;
      60412:data<=16'd3574;
      60413:data<=16'd1955;
      60414:data<=16'd2370;
      60415:data<=16'd1536;
      60416:data<=16'd1180;
      60417:data<=16'd1424;
      60418:data<=16'd1641;
      60419:data<=16'd1060;
      60420:data<=16'd14;
      60421:data<=16'd258;
      60422:data<=-16'd91;
      60423:data<=16'd220;
      60424:data<=16'd1500;
      60425:data<=16'd15;
      60426:data<=-16'd1152;
      60427:data<=-16'd914;
      60428:data<=-16'd1938;
      60429:data<=-16'd2290;
      60430:data<=-16'd2188;
      60431:data<=-16'd2106;
      60432:data<=-16'd1739;
      60433:data<=-16'd2234;
      60434:data<=-16'd2262;
      60435:data<=-16'd2218;
      60436:data<=-16'd2528;
      60437:data<=-16'd3251;
      60438:data<=-16'd4955;
      60439:data<=-16'd4009;
      60440:data<=-16'd5615;
      60441:data<=-16'd14340;
      60442:data<=-16'd17870;
      60443:data<=-16'd15822;
      60444:data<=-16'd16680;
      60445:data<=-16'd15857;
      60446:data<=-16'd14308;
      60447:data<=-16'd14871;
      60448:data<=-16'd13958;
      60449:data<=-16'd14072;
      60450:data<=-16'd15112;
      60451:data<=-16'd14612;
      60452:data<=-16'd14663;
      60453:data<=-16'd14289;
      60454:data<=-16'd13080;
      60455:data<=-16'd12363;
      60456:data<=-16'd11987;
      60457:data<=-16'd12217;
      60458:data<=-16'd11975;
      60459:data<=-16'd11486;
      60460:data<=-16'd11036;
      60461:data<=-16'd10081;
      60462:data<=-16'd10721;
      60463:data<=-16'd11512;
      60464:data<=-16'd11062;
      60465:data<=-16'd11650;
      60466:data<=-16'd12040;
      60467:data<=-16'd12273;
      60468:data<=-16'd12499;
      60469:data<=-16'd11307;
      60470:data<=-16'd11106;
      60471:data<=-16'd10492;
      60472:data<=-16'd9703;
      60473:data<=-16'd11418;
      60474:data<=-16'd7511;
      60475:data<=16'd1121;
      60476:data<=16'd2572;
      60477:data<=16'd740;
      60478:data<=16'd1826;
      60479:data<=16'd2153;
      60480:data<=16'd1680;
      60481:data<=16'd1839;
      60482:data<=16'd1814;
      60483:data<=16'd1648;
      60484:data<=16'd1792;
      60485:data<=16'd2144;
      60486:data<=16'd1569;
      60487:data<=16'd509;
      60488:data<=-16'd11;
      60489:data<=-16'd362;
      60490:data<=-16'd276;
      60491:data<=-16'd121;
      60492:data<=-16'd194;
      60493:data<=-16'd285;
      60494:data<=-16'd588;
      60495:data<=-16'd340;
      60496:data<=-16'd593;
      60497:data<=-16'd1034;
      60498:data<=16'd168;
      60499:data<=-16'd384;
      60500:data<=-16'd2241;
      60501:data<=-16'd1850;
      60502:data<=-16'd1635;
      60503:data<=-16'd1413;
      60504:data<=-16'd1315;
      60505:data<=-16'd2328;
      60506:data<=-16'd781;
      60507:data<=-16'd2093;
      60508:data<=-16'd9394;
      60509:data<=-16'd12007;
      60510:data<=-16'd10343;
      60511:data<=-16'd10827;
      60512:data<=-16'd10916;
      60513:data<=-16'd11028;
      60514:data<=-16'd11570;
      60515:data<=-16'd10648;
      60516:data<=-16'd9928;
      60517:data<=-16'd9464;
      60518:data<=-16'd9078;
      60519:data<=-16'd8872;
      60520:data<=-16'd8062;
      60521:data<=-16'd8126;
      60522:data<=-16'd7965;
      60523:data<=-16'd6643;
      60524:data<=-16'd7077;
      60525:data<=-16'd8492;
      60526:data<=-16'd8636;
      60527:data<=-16'd7689;
      60528:data<=-16'd6532;
      60529:data<=-16'd6384;
      60530:data<=-16'd6247;
      60531:data<=-16'd5638;
      60532:data<=-16'd5342;
      60533:data<=-16'd4658;
      60534:data<=-16'd4639;
      60535:data<=-16'd4752;
      60536:data<=-16'd3877;
      60537:data<=-16'd4602;
      60538:data<=-16'd5068;
      60539:data<=-16'd4666;
      60540:data<=-16'd6040;
      60541:data<=-16'd1868;
      60542:data<=16'd7793;
      60543:data<=16'd9832;
      60544:data<=16'd6828;
      60545:data<=16'd7570;
      60546:data<=16'd7961;
      60547:data<=16'd7131;
      60548:data<=16'd7824;
      60549:data<=16'd6519;
      60550:data<=16'd3369;
      60551:data<=16'd2604;
      60552:data<=16'd3310;
      60553:data<=16'd3090;
      60554:data<=16'd2726;
      60555:data<=16'd2952;
      60556:data<=16'd2925;
      60557:data<=16'd2754;
      60558:data<=16'd3177;
      60559:data<=16'd3162;
      60560:data<=16'd2406;
      60561:data<=16'd2631;
      60562:data<=16'd2661;
      60563:data<=16'd889;
      60564:data<=16'd258;
      60565:data<=16'd1064;
      60566:data<=16'd842;
      60567:data<=16'd1207;
      60568:data<=16'd1480;
      60569:data<=16'd425;
      60570:data<=16'd1242;
      60571:data<=16'd1579;
      60572:data<=16'd505;
      60573:data<=16'd2387;
      60574:data<=-16'd118;
      60575:data<=-16'd10088;
      60576:data<=-16'd14348;
      60577:data<=-16'd12293;
      60578:data<=-16'd12284;
      60579:data<=-16'd11785;
      60580:data<=-16'd10243;
      60581:data<=-16'd10401;
      60582:data<=-16'd10119;
      60583:data<=-16'd9086;
      60584:data<=-16'd8646;
      60585:data<=-16'd8194;
      60586:data<=-16'd7385;
      60587:data<=-16'd7445;
      60588:data<=-16'd8777;
      60589:data<=-16'd8874;
      60590:data<=-16'd7664;
      60591:data<=-16'd6704;
      60592:data<=-16'd4965;
      60593:data<=-16'd3996;
      60594:data<=-16'd4137;
      60595:data<=-16'd2943;
      60596:data<=-16'd2620;
      60597:data<=-16'd3192;
      60598:data<=-16'd2171;
      60599:data<=-16'd1328;
      60600:data<=-16'd1130;
      60601:data<=-16'd1406;
      60602:data<=-16'd1682;
      60603:data<=-16'd664;
      60604:data<=-16'd520;
      60605:data<=-16'd264;
      60606:data<=16'd332;
      60607:data<=-16'd905;
      60608:data<=16'd3805;
      60609:data<=16'd13461;
      60610:data<=16'd14778;
      60611:data<=16'd11960;
      60612:data<=16'd13229;
      60613:data<=16'd14167;
      60614:data<=16'd13981;
      60615:data<=16'd14107;
      60616:data<=16'd13668;
      60617:data<=16'd13292;
      60618:data<=16'd12854;
      60619:data<=16'd12700;
      60620:data<=16'd12422;
      60621:data<=16'd11599;
      60622:data<=16'd11512;
      60623:data<=16'd11154;
      60624:data<=16'd10998;
      60625:data<=16'd12169;
      60626:data<=16'd12383;
      60627:data<=16'd11928;
      60628:data<=16'd11859;
      60629:data<=16'd11344;
      60630:data<=16'd10766;
      60631:data<=16'd10404;
      60632:data<=16'd10214;
      60633:data<=16'd9250;
      60634:data<=16'd7818;
      60635:data<=16'd7359;
      60636:data<=16'd6532;
      60637:data<=16'd7042;
      60638:data<=16'd8801;
      60639:data<=16'd8378;
      60640:data<=16'd9380;
      60641:data<=16'd7345;
      60642:data<=-16'd2937;
      60643:data<=-16'd7260;
      60644:data<=-16'd4128;
      60645:data<=-16'd4763;
      60646:data<=-16'd4584;
      60647:data<=-16'd3203;
      60648:data<=-16'd4361;
      60649:data<=-16'd3215;
      60650:data<=-16'd1591;
      60651:data<=-16'd1407;
      60652:data<=-16'd391;
      60653:data<=-16'd115;
      60654:data<=16'd70;
      60655:data<=16'd271;
      60656:data<=16'd8;
      60657:data<=16'd678;
      60658:data<=16'd626;
      60659:data<=16'd323;
      60660:data<=16'd326;
      60661:data<=-16'd281;
      60662:data<=16'd1227;
      60663:data<=16'd3110;
      60664:data<=16'd2770;
      60665:data<=16'd2845;
      60666:data<=16'd3196;
      60667:data<=16'd3084;
      60668:data<=16'd2808;
      60669:data<=16'd2889;
      60670:data<=16'd3852;
      60671:data<=16'd3330;
      60672:data<=16'd2886;
      60673:data<=16'd3039;
      60674:data<=16'd2276;
      60675:data<=16'd8810;
      60676:data<=16'd19594;
      60677:data<=16'd20850;
      60678:data<=16'd18178;
      60679:data<=16'd18225;
      60680:data<=16'd17006;
      60681:data<=16'd16416;
      60682:data<=16'd16389;
      60683:data<=16'd15208;
      60684:data<=16'd14986;
      60685:data<=16'd14446;
      60686:data<=16'd13529;
      60687:data<=16'd13725;
      60688:data<=16'd14052;
      60689:data<=16'd14032;
      60690:data<=16'd13336;
      60691:data<=16'd12668;
      60692:data<=16'd12248;
      60693:data<=16'd11402;
      60694:data<=16'd11224;
      60695:data<=16'd10939;
      60696:data<=16'd9897;
      60697:data<=16'd9379;
      60698:data<=16'd9074;
      60699:data<=16'd8989;
      60700:data<=16'd9289;
      60701:data<=16'd10170;
      60702:data<=16'd10530;
      60703:data<=16'd8916;
      60704:data<=16'd8804;
      60705:data<=16'd9100;
      60706:data<=16'd7700;
      60707:data<=16'd9232;
      60708:data<=16'd6432;
      60709:data<=-16'd4073;
      60710:data<=-16'd7497;
      60711:data<=-16'd5491;
      60712:data<=-16'd6187;
      60713:data<=-16'd4128;
      60714:data<=-16'd2399;
      60715:data<=-16'd3735;
      60716:data<=-16'd3251;
      60717:data<=-16'd3509;
      60718:data<=-16'd4866;
      60719:data<=-16'd4918;
      60720:data<=-16'd5048;
      60721:data<=-16'd4713;
      60722:data<=-16'd4369;
      60723:data<=-16'd4634;
      60724:data<=-16'd4488;
      60725:data<=-16'd3759;
      60726:data<=-16'd2258;
      60727:data<=-16'd1915;
      60728:data<=-16'd2403;
      60729:data<=-16'd1580;
      60730:data<=-16'd1698;
      60731:data<=-16'd2326;
      60732:data<=-16'd1915;
      60733:data<=-16'd1794;
      60734:data<=-16'd1616;
      60735:data<=-16'd2246;
      60736:data<=-16'd2675;
      60737:data<=-16'd1219;
      60738:data<=-16'd329;
      60739:data<=16'd611;
      60740:data<=16'd443;
      60741:data<=-16'd428;
      60742:data<=16'd5847;
      60743:data<=16'd13562;
      60744:data<=16'd13314;
      60745:data<=16'd11753;
      60746:data<=16'd11656;
      60747:data<=16'd10537;
      60748:data<=16'd10154;
      60749:data<=16'd9498;
      60750:data<=16'd9288;
      60751:data<=16'd10379;
      60752:data<=16'd10034;
      60753:data<=16'd9276;
      60754:data<=16'd9054;
      60755:data<=16'd8241;
      60756:data<=16'd7506;
      60757:data<=16'd6948;
      60758:data<=16'd6581;
      60759:data<=16'd6830;
      60760:data<=16'd7453;
      60761:data<=16'd7853;
      60762:data<=16'd7924;
      60763:data<=16'd8417;
      60764:data<=16'd8382;
      60765:data<=16'd7600;
      60766:data<=16'd7329;
      60767:data<=16'd6865;
      60768:data<=16'd6787;
      60769:data<=16'd6475;
      60770:data<=16'd4908;
      60771:data<=16'd5136;
      60772:data<=16'd5112;
      60773:data<=16'd4071;
      60774:data<=16'd5695;
      60775:data<=16'd2487;
      60776:data<=-16'd6448;
      60777:data<=-16'd8824;
      60778:data<=-16'd7116;
      60779:data<=-16'd7962;
      60780:data<=-16'd7721;
      60781:data<=-16'd6827;
      60782:data<=-16'd7122;
      60783:data<=-16'd7068;
      60784:data<=-16'd6740;
      60785:data<=-16'd6472;
      60786:data<=-16'd6329;
      60787:data<=-16'd5911;
      60788:data<=-16'd4966;
      60789:data<=-16'd4143;
      60790:data<=-16'd3751;
      60791:data<=-16'd4030;
      60792:data<=-16'd3970;
      60793:data<=-16'd3759;
      60794:data<=-16'd4485;
      60795:data<=-16'd4267;
      60796:data<=-16'd3721;
      60797:data<=-16'd4209;
      60798:data<=-16'd4193;
      60799:data<=-16'd4416;
      60800:data<=-16'd4320;
      60801:data<=-16'd4047;
      60802:data<=-16'd5908;
      60803:data<=-16'd6617;
      60804:data<=-16'd5930;
      60805:data<=-16'd6252;
      60806:data<=-16'd5556;
      60807:data<=-16'd6334;
      60808:data<=-16'd6288;
      60809:data<=16'd1058;
      60810:data<=16'd7602;
      60811:data<=16'd7347;
      60812:data<=16'd5797;
      60813:data<=16'd4296;
      60814:data<=16'd3099;
      60815:data<=16'd3001;
      60816:data<=16'd2560;
      60817:data<=16'd2137;
      60818:data<=16'd1701;
      60819:data<=16'd1293;
      60820:data<=16'd1286;
      60821:data<=16'd884;
      60822:data<=16'd564;
      60823:data<=16'd387;
      60824:data<=16'd306;
      60825:data<=-16'd140;
      60826:data<=-16'd1898;
      60827:data<=-16'd2641;
      60828:data<=-16'd2613;
      60829:data<=-16'd3334;
      60830:data<=-16'd2604;
      60831:data<=-16'd2259;
      60832:data<=-16'd3066;
      60833:data<=-16'd2569;
      60834:data<=-16'd2685;
      60835:data<=-16'd2645;
      60836:data<=-16'd2350;
      60837:data<=-16'd4030;
      60838:data<=-16'd4363;
      60839:data<=-16'd4855;
      60840:data<=-16'd5991;
      60841:data<=-16'd3771;
      60842:data<=-16'd7151;
      60843:data<=-16'd16680;
      60844:data<=-16'd17998;
      60845:data<=-16'd14704;
      60846:data<=-16'd15035;
      60847:data<=-16'd14784;
      60848:data<=-16'd13785;
      60849:data<=-16'd13446;
      60850:data<=-16'd13224;
      60851:data<=-16'd14131;
      60852:data<=-16'd14054;
      60853:data<=-16'd12860;
      60854:data<=-16'd12712;
      60855:data<=-16'd12358;
      60856:data<=-16'd11826;
      60857:data<=-16'd11720;
      60858:data<=-16'd10986;
      60859:data<=-16'd10342;
      60860:data<=-16'd10216;
      60861:data<=-16'd9812;
      60862:data<=-16'd9843;
      60863:data<=-16'd10775;
      60864:data<=-16'd11376;
      60865:data<=-16'd11359;
      60866:data<=-16'd11229;
      60867:data<=-16'd10522;
      60868:data<=-16'd9935;
      60869:data<=-16'd9859;
      60870:data<=-16'd9109;
      60871:data<=-16'd8774;
      60872:data<=-16'd8593;
      60873:data<=-16'd7283;
      60874:data<=-16'd7824;
      60875:data<=-16'd7794;
      60876:data<=-16'd1689;
      60877:data<=16'd4358;
      60878:data<=16'd4639;
      60879:data<=16'd3680;
      60880:data<=16'd3603;
      60881:data<=16'd3271;
      60882:data<=16'd3454;
      60883:data<=16'd3820;
      60884:data<=16'd3576;
      60885:data<=16'd2708;
      60886:data<=16'd1398;
      60887:data<=16'd517;
      60888:data<=-16'd115;
      60889:data<=-16'd1439;
      60890:data<=-16'd2350;
      60891:data<=-16'd1977;
      60892:data<=-16'd1707;
      60893:data<=-16'd1689;
      60894:data<=-16'd1416;
      60895:data<=-16'd1744;
      60896:data<=-16'd1892;
      60897:data<=-16'd1410;
      60898:data<=-16'd1324;
      60899:data<=-16'd908;
      60900:data<=-16'd1359;
      60901:data<=-16'd3196;
      60902:data<=-16'd3046;
      60903:data<=-16'd2649;
      60904:data<=-16'd3627;
      60905:data<=-16'd2977;
      60906:data<=-16'd3151;
      60907:data<=-16'd3253;
      60908:data<=-16'd358;
      60909:data<=-16'd3980;
      60910:data<=-16'd14119;
      60911:data<=-16'd16745;
      60912:data<=-16'd13884;
      60913:data<=-16'd14352;
      60914:data<=-16'd15465;
      60915:data<=-16'd15103;
      60916:data<=-16'd14445;
      60917:data<=-16'd13480;
      60918:data<=-16'd12813;
      60919:data<=-16'd12110;
      60920:data<=-16'd11195;
      60921:data<=-16'd10742;
      60922:data<=-16'd10246;
      60923:data<=-16'd9512;
      60924:data<=-16'd9012;
      60925:data<=-16'd9160;
      60926:data<=-16'd10073;
      60927:data<=-16'd10437;
      60928:data<=-16'd9110;
      60929:data<=-16'd7363;
      60930:data<=-16'd6630;
      60931:data<=-16'd6193;
      60932:data<=-16'd5988;
      60933:data<=-16'd6328;
      60934:data<=-16'd5812;
      60935:data<=-16'd5213;
      60936:data<=-16'd5062;
      60937:data<=-16'd3802;
      60938:data<=-16'd4008;
      60939:data<=-16'd5521;
      60940:data<=-16'd5048;
      60941:data<=-16'd5645;
      60942:data<=-16'd4516;
      60943:data<=16'd3472;
      60944:data<=16'd9468;
      60945:data<=16'd9054;
      60946:data<=16'd8220;
      60947:data<=16'd7674;
      60948:data<=16'd7627;
      60949:data<=16'd8313;
      60950:data<=16'd7310;
      60951:data<=16'd5697;
      60952:data<=16'd4567;
      60953:data<=16'd4316;
      60954:data<=16'd5024;
      60955:data<=16'd4655;
      60956:data<=16'd4323;
      60957:data<=16'd4558;
      60958:data<=16'd3900;
      60959:data<=16'd3999;
      60960:data<=16'd4319;
      60961:data<=16'd3997;
      60962:data<=16'd4235;
      60963:data<=16'd3542;
      60964:data<=16'd2343;
      60965:data<=16'd2253;
      60966:data<=16'd2493;
      60967:data<=16'd2779;
      60968:data<=16'd2749;
      60969:data<=16'd2852;
      60970:data<=16'd1930;
      60971:data<=-16'd505;
      60972:data<=-16'd108;
      60973:data<=16'd673;
      60974:data<=-16'd108;
      60975:data<=16'd1730;
      60976:data<=-16'd2246;
      60977:data<=-16'd13191;
      60978:data<=-16'd15832;
      60979:data<=-16'd13104;
      60980:data<=-16'd13432;
      60981:data<=-16'd12439;
      60982:data<=-16'd11330;
      60983:data<=-16'd11241;
      60984:data<=-16'd9949;
      60985:data<=-16'd9636;
      60986:data<=-16'd9089;
      60987:data<=-16'd7997;
      60988:data<=-16'd8765;
      60989:data<=-16'd9335;
      60990:data<=-16'd8758;
      60991:data<=-16'd7900;
      60992:data<=-16'd7186;
      60993:data<=-16'd7222;
      60994:data<=-16'd6848;
      60995:data<=-16'd6273;
      60996:data<=-16'd6185;
      60997:data<=-16'd5494;
      60998:data<=-16'd4895;
      60999:data<=-16'd5096;
      61000:data<=-16'd5204;
      61001:data<=-16'd4780;
      61002:data<=-16'd4428;
      61003:data<=-16'd4123;
      61004:data<=-16'd2960;
      61005:data<=-16'd2641;
      61006:data<=-16'd2772;
      61007:data<=-16'd1607;
      61008:data<=-16'd2602;
      61009:data<=-16'd1557;
      61010:data<=16'd6887;
      61011:data<=16'd12361;
      61012:data<=16'd12051;
      61013:data<=16'd13870;
      61014:data<=16'd15224;
      61015:data<=16'd14586;
      61016:data<=16'd14885;
      61017:data<=16'd14490;
      61018:data<=16'd13594;
      61019:data<=16'd13074;
      61020:data<=16'd12766;
      61021:data<=16'd12806;
      61022:data<=16'd12040;
      61023:data<=16'd11242;
      61024:data<=16'd10742;
      61025:data<=16'd10367;
      61026:data<=16'd11562;
      61027:data<=16'd12563;
      61028:data<=16'd12393;
      61029:data<=16'd12245;
      61030:data<=16'd11555;
      61031:data<=16'd11083;
      61032:data<=16'd11074;
      61033:data<=16'd11062;
      61034:data<=16'd10960;
      61035:data<=16'd10288;
      61036:data<=16'd10660;
      61037:data<=16'd10257;
      61038:data<=16'd8646;
      61039:data<=16'd10383;
      61040:data<=16'd10807;
      61041:data<=16'd9448;
      61042:data<=16'd11887;
      61043:data<=16'd7899;
      61044:data<=-16'd2546;
      61045:data<=-16'd4722;
      61046:data<=-16'd2857;
      61047:data<=-16'd3263;
      61048:data<=-16'd2604;
      61049:data<=-16'd2766;
      61050:data<=-16'd2940;
      61051:data<=-16'd1306;
      61052:data<=16'd9;
      61053:data<=16'd748;
      61054:data<=-16'd227;
      61055:data<=-16'd1713;
      61056:data<=-16'd1201;
      61057:data<=-16'd699;
      61058:data<=-16'd873;
      61059:data<=-16'd923;
      61060:data<=-16'd694;
      61061:data<=-16'd426;
      61062:data<=-16'd1104;
      61063:data<=-16'd710;
      61064:data<=16'd1190;
      61065:data<=16'd1771;
      61066:data<=16'd1339;
      61067:data<=16'd873;
      61068:data<=16'd860;
      61069:data<=16'd1158;
      61070:data<=16'd1266;
      61071:data<=16'd2038;
      61072:data<=16'd1636;
      61073:data<=16'd1086;
      61074:data<=16'd2250;
      61075:data<=16'd757;
      61076:data<=16'd2523;
      61077:data<=16'd12686;
      61078:data<=16'd17848;
      61079:data<=16'd15638;
      61080:data<=16'd15242;
      61081:data<=16'd14932;
      61082:data<=16'd14093;
      61083:data<=16'd14058;
      61084:data<=16'd13079;
      61085:data<=16'd12460;
      61086:data<=16'd11738;
      61087:data<=16'd10972;
      61088:data<=16'd11762;
      61089:data<=16'd12216;
      61090:data<=16'd12179;
      61091:data<=16'd11729;
      61092:data<=16'd10587;
      61093:data<=16'd10721;
      61094:data<=16'd10780;
      61095:data<=16'd9955;
      61096:data<=16'd10154;
      61097:data<=16'd10840;
      61098:data<=16'd11309;
      61099:data<=16'd10944;
      61100:data<=16'd10157;
      61101:data<=16'd10596;
      61102:data<=16'd11562;
      61103:data<=16'd12331;
      61104:data<=16'd11562;
      61105:data<=16'd9712;
      61106:data<=16'd9993;
      61107:data<=16'd9624;
      61108:data<=16'd8619;
      61109:data<=16'd10226;
      61110:data<=16'd6219;
      61111:data<=-16'd3759;
      61112:data<=-16'd6805;
      61113:data<=-16'd4247;
      61114:data<=-16'd3468;
      61115:data<=-16'd2949;
      61116:data<=-16'd2675;
      61117:data<=-16'd3072;
      61118:data<=-16'd2362;
      61119:data<=-16'd1839;
      61120:data<=-16'd2402;
      61121:data<=-16'd2563;
      61122:data<=-16'd1964;
      61123:data<=-16'd1377;
      61124:data<=-16'd1483;
      61125:data<=-16'd2240;
      61126:data<=-16'd1885;
      61127:data<=16'd71;
      61128:data<=16'd784;
      61129:data<=-16'd55;
      61130:data<=-16'd229;
      61131:data<=-16'd97;
      61132:data<=16'd6;
      61133:data<=-16'd100;
      61134:data<=-16'd751;
      61135:data<=-16'd802;
      61136:data<=-16'd1158;
      61137:data<=-16'd1510;
      61138:data<=-16'd660;
      61139:data<=-16'd1134;
      61140:data<=-16'd1096;
      61141:data<=-16'd32;
      61142:data<=-16'd2272;
      61143:data<=-16'd528;
      61144:data<=16'd8739;
      61145:data<=16'd13069;
      61146:data<=16'd11247;
      61147:data<=16'd10860;
      61148:data<=16'd10572;
      61149:data<=16'd9527;
      61150:data<=16'd9188;
      61151:data<=16'd9564;
      61152:data<=16'd10519;
      61153:data<=16'd10220;
      61154:data<=16'd9098;
      61155:data<=16'd8704;
      61156:data<=16'd8220;
      61157:data<=16'd7877;
      61158:data<=16'd7412;
      61159:data<=16'd6771;
      61160:data<=16'd6865;
      61161:data<=16'd6249;
      61162:data<=16'd5372;
      61163:data<=16'd5683;
      61164:data<=16'd6211;
      61165:data<=16'd6931;
      61166:data<=16'd6962;
      61167:data<=16'd6061;
      61168:data<=16'd5926;
      61169:data<=16'd5752;
      61170:data<=16'd5796;
      61171:data<=16'd5855;
      61172:data<=16'd4472;
      61173:data<=16'd4253;
      61174:data<=16'd3974;
      61175:data<=16'd2948;
      61176:data<=16'd5268;
      61177:data<=16'd2999;
      61178:data<=-16'd7063;
      61179:data<=-16'd10373;
      61180:data<=-16'd6707;
      61181:data<=-16'd5799;
      61182:data<=-16'd5412;
      61183:data<=-16'd4904;
      61184:data<=-16'd5313;
      61185:data<=-16'd4548;
      61186:data<=-16'd4828;
      61187:data<=-16'd5695;
      61188:data<=-16'd4511;
      61189:data<=-16'd3037;
      61190:data<=-16'd2127;
      61191:data<=-16'd2117;
      61192:data<=-16'd2901;
      61193:data<=-16'd2711;
      61194:data<=-16'd2428;
      61195:data<=-16'd2685;
      61196:data<=-16'd2544;
      61197:data<=-16'd2678;
      61198:data<=-16'd2945;
      61199:data<=-16'd2872;
      61200:data<=-16'd3196;
      61201:data<=-16'd3506;
      61202:data<=-16'd3392;
      61203:data<=-16'd3680;
      61204:data<=-16'd3955;
      61205:data<=-16'd3635;
      61206:data<=-16'd3788;
      61207:data<=-16'd3507;
      61208:data<=-16'd2857;
      61209:data<=-16'd4426;
      61210:data<=-16'd2514;
      61211:data<=16'd6363;
      61212:data<=16'd10957;
      61213:data<=16'd8617;
      61214:data<=16'd7326;
      61215:data<=16'd6135;
      61216:data<=16'd4830;
      61217:data<=16'd5438;
      61218:data<=16'd4921;
      61219:data<=16'd3988;
      61220:data<=16'd3806;
      61221:data<=16'd3228;
      61222:data<=16'd2810;
      61223:data<=16'd1249;
      61224:data<=-16'd246;
      61225:data<=16'd224;
      61226:data<=-16'd244;
      61227:data<=-16'd1510;
      61228:data<=-16'd2021;
      61229:data<=-16'd2400;
      61230:data<=-16'd2414;
      61231:data<=-16'd2690;
      61232:data<=-16'd2739;
      61233:data<=-16'd2168;
      61234:data<=-16'd2177;
      61235:data<=-16'd2112;
      61236:data<=-16'd2179;
      61237:data<=-16'd1944;
      61238:data<=-16'd1460;
      61239:data<=-16'd2943;
      61240:data<=-16'd3767;
      61241:data<=-16'd3900;
      61242:data<=-16'd4636;
      61243:data<=-16'd2734;
      61244:data<=-16'd5835;
      61245:data<=-16'd15901;
      61246:data<=-16'd18318;
      61247:data<=-16'd15397;
      61248:data<=-16'd16058;
      61249:data<=-16'd15305;
      61250:data<=-16'd13794;
      61251:data<=-16'd14346;
      61252:data<=-16'd14660;
      61253:data<=-16'd15109;
      61254:data<=-16'd14750;
      61255:data<=-16'd13728;
      61256:data<=-16'd13368;
      61257:data<=-16'd12555;
      61258:data<=-16'd12196;
      61259:data<=-16'd12008;
      61260:data<=-16'd11367;
      61261:data<=-16'd11417;
      61262:data<=-16'd10746;
      61263:data<=-16'd9806;
      61264:data<=-16'd9770;
      61265:data<=-16'd9333;
      61266:data<=-16'd9081;
      61267:data<=-16'd9226;
      61268:data<=-16'd9132;
      61269:data<=-16'd9036;
      61270:data<=-16'd8822;
      61271:data<=-16'd8376;
      61272:data<=-16'd7521;
      61273:data<=-16'd7686;
      61274:data<=-16'd7746;
      61275:data<=-16'd6369;
      61276:data<=-16'd7950;
      61277:data<=-16'd7039;
      61278:data<=16'd1979;
      61279:data<=16'd6537;
      61280:data<=16'd4558;
      61281:data<=16'd4766;
      61282:data<=16'd4305;
      61283:data<=16'd3550;
      61284:data<=16'd4194;
      61285:data<=16'd3295;
      61286:data<=16'd3106;
      61287:data<=16'd3169;
      61288:data<=16'd2484;
      61289:data<=16'd2202;
      61290:data<=16'd652;
      61291:data<=16'd341;
      61292:data<=16'd805;
      61293:data<=-16'd417;
      61294:data<=16'd203;
      61295:data<=16'd525;
      61296:data<=-16'd396;
      61297:data<=16'd352;
      61298:data<=-16'd33;
      61299:data<=16'd103;
      61300:data<=16'd1231;
      61301:data<=-16'd133;
      61302:data<=-16'd1190;
      61303:data<=-16'd1920;
      61304:data<=-16'd2021;
      61305:data<=-16'd804;
      61306:data<=-16'd2543;
      61307:data<=-16'd3867;
      61308:data<=-16'd3930;
      61309:data<=-16'd4764;
      61310:data<=-16'd2156;
      61311:data<=-16'd5148;
      61312:data<=-16'd15605;
      61313:data<=-16'd17540;
      61314:data<=-16'd15390;
      61315:data<=-16'd17103;
      61316:data<=-16'd16286;
      61317:data<=-16'd14971;
      61318:data<=-16'd14645;
      61319:data<=-16'd13315;
      61320:data<=-16'd13277;
      61321:data<=-16'd12704;
      61322:data<=-16'd11623;
      61323:data<=-16'd11458;
      61324:data<=-16'd10417;
      61325:data<=-16'd10038;
      61326:data<=-16'd10511;
      61327:data<=-16'd10671;
      61328:data<=-16'd10936;
      61329:data<=-16'd10040;
      61330:data<=-16'd9092;
      61331:data<=-16'd9359;
      61332:data<=-16'd9270;
      61333:data<=-16'd8689;
      61334:data<=-16'd8122;
      61335:data<=-16'd7884;
      61336:data<=-16'd7752;
      61337:data<=-16'd7494;
      61338:data<=-16'd7160;
      61339:data<=-16'd6745;
      61340:data<=-16'd7996;
      61341:data<=-16'd8341;
      61342:data<=-16'd6299;
      61343:data<=-16'd7319;
      61344:data<=-16'd5291;
      61345:data<=16'd4469;
      61346:data<=16'd8587;
      61347:data<=16'd6320;
      61348:data<=16'd7174;
      61349:data<=16'd8543;
      61350:data<=16'd8801;
      61351:data<=16'd8478;
      61352:data<=16'd6777;
      61353:data<=16'd5968;
      61354:data<=16'd5668;
      61355:data<=16'd5574;
      61356:data<=16'd5686;
      61357:data<=16'd4831;
      61358:data<=16'd4848;
      61359:data<=16'd4834;
      61360:data<=16'd4270;
      61361:data<=16'd4939;
      61362:data<=16'd4701;
      61363:data<=16'd4300;
      61364:data<=16'd4129;
      61365:data<=16'd2343;
      61366:data<=16'd2261;
      61367:data<=16'd3162;
      61368:data<=16'd2719;
      61369:data<=16'd2739;
      61370:data<=16'd2299;
      61371:data<=16'd2629;
      61372:data<=16'd3315;
      61373:data<=16'd2050;
      61374:data<=16'd2561;
      61375:data<=16'd2602;
      61376:data<=16'd1134;
      61377:data<=16'd2396;
      61378:data<=-16'd2027;
      61379:data<=-16'd11849;
      61380:data<=-16'd13655;
      61381:data<=-16'd11347;
      61382:data<=-16'd11438;
      61383:data<=-16'd10580;
      61384:data<=-16'd9796;
      61385:data<=-16'd9383;
      61386:data<=-16'd8458;
      61387:data<=-16'd8341;
      61388:data<=-16'd7746;
      61389:data<=-16'd7353;
      61390:data<=-16'd8787;
      61391:data<=-16'd9908;
      61392:data<=-16'd9639;
      61393:data<=-16'd9148;
      61394:data<=-16'd8769;
      61395:data<=-16'd8184;
      61396:data<=-16'd7559;
      61397:data<=-16'd6678;
      61398:data<=-16'd5908;
      61399:data<=-16'd6414;
      61400:data<=-16'd6581;
      61401:data<=-16'd5824;
      61402:data<=-16'd5629;
      61403:data<=-16'd4874;
      61404:data<=-16'd4490;
      61405:data<=-16'd4642;
      61406:data<=-16'd3303;
      61407:data<=-16'd3277;
      61408:data<=-16'd3136;
      61409:data<=-16'd1557;
      61410:data<=-16'd3316;
      61411:data<=-16'd741;
      61412:data<=16'd9398;
      61413:data<=16'd12885;
      61414:data<=16'd11062;
      61415:data<=16'd12765;
      61416:data<=16'd13156;
      61417:data<=16'd12038;
      61418:data<=16'd12399;
      61419:data<=16'd12125;
      61420:data<=16'd11564;
      61421:data<=16'd10927;
      61422:data<=16'd10346;
      61423:data<=16'd10351;
      61424:data<=16'd9837;
      61425:data<=16'd9568;
      61426:data<=16'd9342;
      61427:data<=16'd9098;
      61428:data<=16'd10173;
      61429:data<=16'd10387;
      61430:data<=16'd9688;
      61431:data<=16'd9853;
      61432:data<=16'd10078;
      61433:data<=16'd11318;
      61434:data<=16'd12401;
      61435:data<=16'd11488;
      61436:data<=16'd10974;
      61437:data<=16'd10759;
      61438:data<=16'd10396;
      61439:data<=16'd10575;
      61440:data<=16'd10531;
      61441:data<=16'd11156;
      61442:data<=16'd10571;
      61443:data<=16'd9415;
      61444:data<=16'd11095;
      61445:data<=16'd7083;
      61446:data<=-16'd3095;
      61447:data<=-16'd5369;
      61448:data<=-16'd2810;
      61449:data<=-16'd3342;
      61450:data<=-16'd2986;
      61451:data<=-16'd2713;
      61452:data<=-16'd2723;
      61453:data<=-16'd669;
      61454:data<=-16'd241;
      61455:data<=-16'd481;
      61456:data<=16'd431;
      61457:data<=16'd187;
      61458:data<=16'd409;
      61459:data<=16'd790;
      61460:data<=16'd23;
      61461:data<=16'd479;
      61462:data<=16'd1033;
      61463:data<=16'd725;
      61464:data<=16'd1486;
      61465:data<=16'd2417;
      61466:data<=16'd2585;
      61467:data<=16'd2438;
      61468:data<=16'd2121;
      61469:data<=16'd2358;
      61470:data<=16'd2641;
      61471:data<=16'd2061;
      61472:data<=16'd2100;
      61473:data<=16'd2922;
      61474:data<=16'd2111;
      61475:data<=16'd963;
      61476:data<=16'd893;
      61477:data<=16'd100;
      61478:data<=16'd3745;
      61479:data<=16'd13302;
      61480:data<=16'd16783;
      61481:data<=16'd14001;
      61482:data<=16'd14087;
      61483:data<=16'd14072;
      61484:data<=16'd12651;
      61485:data<=16'd12622;
      61486:data<=16'd11985;
      61487:data<=16'd11553;
      61488:data<=16'd11254;
      61489:data<=16'd10231;
      61490:data<=16'd10863;
      61491:data<=16'd11423;
      61492:data<=16'd10966;
      61493:data<=16'd10815;
      61494:data<=16'd9952;
      61495:data<=16'd9677;
      61496:data<=16'd9721;
      61497:data<=16'd8645;
      61498:data<=16'd8288;
      61499:data<=16'd8396;
      61500:data<=16'd8288;
      61501:data<=16'd7884;
      61502:data<=16'd7658;
      61503:data<=16'd9233;
      61504:data<=16'd9544;
      61505:data<=16'd8070;
      61506:data<=16'd7915;
      61507:data<=16'd7424;
      61508:data<=16'd7142;
      61509:data<=16'd6686;
      61510:data<=16'd5444;
      61511:data<=16'd6563;
      61512:data<=16'd2488;
      61513:data<=-16'd7350;
      61514:data<=-16'd8624;
      61515:data<=-16'd4945;
      61516:data<=-16'd4660;
      61517:data<=-16'd3791;
      61518:data<=-16'd3209;
      61519:data<=-16'd2936;
      61520:data<=-16'd2040;
      61521:data<=-16'd2679;
      61522:data<=-16'd2297;
      61523:data<=-16'd1962;
      61524:data<=-16'd2617;
      61525:data<=-16'd1621;
      61526:data<=-16'd2015;
      61527:data<=-16'd2523;
      61528:data<=-16'd626;
      61529:data<=-16'd67;
      61530:data<=16'd121;
      61531:data<=16'd579;
      61532:data<=-16'd367;
      61533:data<=-16'd704;
      61534:data<=-16'd549;
      61535:data<=-16'd569;
      61536:data<=-16'd402;
      61537:data<=-16'd738;
      61538:data<=-16'd1121;
      61539:data<=-16'd584;
      61540:data<=16'd1245;
      61541:data<=16'd1839;
      61542:data<=16'd1146;
      61543:data<=16'd1807;
      61544:data<=16'd895;
      61545:data<=16'd3096;
      61546:data<=16'd12533;
      61547:data<=16'd15644;
      61548:data<=16'd11994;
      61549:data<=16'd12486;
      61550:data<=16'd12718;
      61551:data<=16'd11527;
      61552:data<=16'd12008;
      61553:data<=16'd12098;
      61554:data<=16'd12569;
      61555:data<=16'd11541;
      61556:data<=16'd9791;
      61557:data<=16'd10386;
      61558:data<=16'd9485;
      61559:data<=16'd7864;
      61560:data<=16'd7022;
      61561:data<=16'd5629;
      61562:data<=16'd5946;
      61563:data<=16'd5536;
      61564:data<=16'd4444;
      61565:data<=16'd5893;
      61566:data<=16'd6361;
      61567:data<=16'd6102;
      61568:data<=16'd6038;
      61569:data<=16'd5066;
      61570:data<=16'd5354;
      61571:data<=16'd4895;
      61572:data<=16'd4018;
      61573:data<=16'd4255;
      61574:data<=16'd3095;
      61575:data<=16'd2881;
      61576:data<=16'd2416;
      61577:data<=16'd1964;
      61578:data<=16'd4440;
      61579:data<=-16'd405;
      61580:data<=-16'd9797;
      61581:data<=-16'd10176;
      61582:data<=-16'd8401;
      61583:data<=-16'd8760;
      61584:data<=-16'd8319;
      61585:data<=-16'd9454;
      61586:data<=-16'd8884;
      61587:data<=-16'd7567;
      61588:data<=-16'd8310;
      61589:data<=-16'd7565;
      61590:data<=-16'd6766;
      61591:data<=-16'd5903;
      61592:data<=-16'd4748;
      61593:data<=-16'd5541;
      61594:data<=-16'd5121;
      61595:data<=-16'd4672;
      61596:data<=-16'd5344;
      61597:data<=-16'd4219;
      61598:data<=-16'd4073;
      61599:data<=-16'd4825;
      61600:data<=-16'd4831;
      61601:data<=-16'd4576;
      61602:data<=-16'd2892;
      61603:data<=-16'd2569;
      61604:data<=-16'd3101;
      61605:data<=-16'd2572;
      61606:data<=-16'd3143;
      61607:data<=-16'd2461;
      61608:data<=-16'd2293;
      61609:data<=-16'd3177;
      61610:data<=-16'd1513;
      61611:data<=-16'd2758;
      61612:data<=-16'd970;
      61613:data<=16'd9212;
      61614:data<=16'd11991;
      61615:data<=16'd8020;
      61616:data<=16'd7338;
      61617:data<=16'd6458;
      61618:data<=16'd6587;
      61619:data<=16'd6657;
      61620:data<=16'd4939;
      61621:data<=16'd5224;
      61622:data<=16'd4451;
      61623:data<=16'd3789;
      61624:data<=16'd4619;
      61625:data<=16'd3418;
      61626:data<=16'd3750;
      61627:data<=16'd3369;
      61628:data<=16'd415;
      61629:data<=16'd509;
      61630:data<=16'd488;
      61631:data<=-16'd323;
      61632:data<=16'd246;
      61633:data<=-16'd390;
      61634:data<=16'd45;
      61635:data<=16'd456;
      61636:data<=-16'd429;
      61637:data<=-16'd18;
      61638:data<=-16'd710;
      61639:data<=-16'd892;
      61640:data<=-16'd931;
      61641:data<=-16'd3412;
      61642:data<=-16'd3383;
      61643:data<=-16'd3495;
      61644:data<=-16'd4595;
      61645:data<=-16'd3551;
      61646:data<=-16'd8587;
      61647:data<=-16'd15373;
      61648:data<=-16'd14636;
      61649:data<=-16'd13512;
      61650:data<=-16'd13285;
      61651:data<=-16'd12410;
      61652:data<=-16'd13286;
      61653:data<=-16'd13446;
      61654:data<=-16'd13697;
      61655:data<=-16'd13662;
      61656:data<=-16'd12352;
      61657:data<=-16'd12728;
      61658:data<=-16'd12542;
      61659:data<=-16'd11790;
      61660:data<=-16'd11712;
      61661:data<=-16'd10504;
      61662:data<=-16'd10833;
      61663:data<=-16'd10869;
      61664:data<=-16'd8940;
      61665:data<=-16'd9608;
      61666:data<=-16'd11074;
      61667:data<=-16'd11461;
      61668:data<=-16'd11218;
      61669:data<=-16'd10138;
      61670:data<=-16'd10592;
      61671:data<=-16'd10428;
      61672:data<=-16'd9353;
      61673:data<=-16'd9380;
      61674:data<=-16'd8058;
      61675:data<=-16'd8029;
      61676:data<=-16'd8078;
      61677:data<=-16'd6470;
      61678:data<=-16'd9186;
      61679:data<=-16'd7561;
      61680:data<=16'd1853;
      61681:data<=16'd4106;
      61682:data<=16'd1774;
      61683:data<=16'd2453;
      61684:data<=16'd2346;
      61685:data<=16'd2338;
      61686:data<=16'd2105;
      61687:data<=16'd1412;
      61688:data<=16'd2182;
      61689:data<=16'd1835;
      61690:data<=16'd836;
      61691:data<=-16'd246;
      61692:data<=-16'd1181;
      61693:data<=-16'd261;
      61694:data<=-16'd673;
      61695:data<=-16'd1359;
      61696:data<=-16'd469;
      61697:data<=-16'd1236;
      61698:data<=-16'd1257;
      61699:data<=-16'd557;
      61700:data<=-16'd1368;
      61701:data<=-16'd822;
      61702:data<=-16'd687;
      61703:data<=-16'd1898;
      61704:data<=-16'd2491;
      61705:data<=-16'd3159;
      61706:data<=-16'd2682;
      61707:data<=-16'd2441;
      61708:data<=-16'd2933;
      61709:data<=-16'd2356;
      61710:data<=-16'd3322;
      61711:data<=-16'd3218;
      61712:data<=-16'd2620;
      61713:data<=-16'd8334;
      61714:data<=-16'd13571;
      61715:data<=-16'd13500;
      61716:data<=-16'd13758;
      61717:data<=-16'd13788;
      61718:data<=-16'd13377;
      61719:data<=-16'd13042;
      61720:data<=-16'd11464;
      61721:data<=-16'd11441;
      61722:data<=-16'd11902;
      61723:data<=-16'd10827;
      61724:data<=-16'd10160;
      61725:data<=-16'd9441;
      61726:data<=-16'd8856;
      61727:data<=-16'd8802;
      61728:data<=-16'd9085;
      61729:data<=-16'd10181;
      61730:data<=-16'd9800;
      61731:data<=-16'd8511;
      61732:data<=-16'd8363;
      61733:data<=-16'd8047;
      61734:data<=-16'd8146;
      61735:data<=-16'd8067;
      61736:data<=-16'd7107;
      61737:data<=-16'd6977;
      61738:data<=-16'd6499;
      61739:data<=-16'd6119;
      61740:data<=-16'd6482;
      61741:data<=-16'd6443;
      61742:data<=-16'd7306;
      61743:data<=-16'd6514;
      61744:data<=-16'd4786;
      61745:data<=-16'd6290;
      61746:data<=-16'd3284;
      61747:data<=16'd5113;
      61748:data<=16'd7559;
      61749:data<=16'd5736;
      61750:data<=16'd5709;
      61751:data<=16'd6053;
      61752:data<=16'd5815;
      61753:data<=16'd4516;
      61754:data<=16'd3401;
      61755:data<=16'd3676;
      61756:data<=16'd3664;
      61757:data<=16'd3554;
      61758:data<=16'd3375;
      61759:data<=16'd2845;
      61760:data<=16'd3163;
      61761:data<=16'd3482;
      61762:data<=16'd3200;
      61763:data<=16'd3062;
      61764:data<=16'd3013;
      61765:data<=16'd2734;
      61766:data<=16'd1864;
      61767:data<=16'd1480;
      61768:data<=16'd1879;
      61769:data<=16'd1874;
      61770:data<=16'd2093;
      61771:data<=16'd2130;
      61772:data<=16'd1765;
      61773:data<=16'd2108;
      61774:data<=16'd1806;
      61775:data<=16'd1384;
      61776:data<=16'd1619;
      61777:data<=16'd887;
      61778:data<=16'd785;
      61779:data<=-16'd444;
      61780:data<=-16'd6290;
      61781:data<=-16'd11095;
      61782:data<=-16'd11198;
      61783:data<=-16'd10114;
      61784:data<=-16'd9215;
      61785:data<=-16'd8621;
      61786:data<=-16'd8243;
      61787:data<=-16'd7800;
      61788:data<=-16'd7741;
      61789:data<=-16'd7279;
      61790:data<=-16'd7063;
      61791:data<=-16'd7961;
      61792:data<=-16'd8093;
      61793:data<=-16'd7322;
      61794:data<=-16'd7021;
      61795:data<=-16'd7059;
      61796:data<=-16'd6567;
      61797:data<=-16'd5398;
      61798:data<=-16'd4816;
      61799:data<=-16'd4725;
      61800:data<=-16'd4467;
      61801:data<=-16'd4578;
      61802:data<=-16'd4135;
      61803:data<=-16'd3425;
      61804:data<=-16'd3333;
      61805:data<=-16'd2757;
      61806:data<=-16'd2710;
      61807:data<=-16'd2708;
      61808:data<=-16'd1453;
      61809:data<=-16'd1319;
      61810:data<=-16'd785;
      61811:data<=16'd149;
      61812:data<=-16'd1463;
      61813:data<=16'd1391;
      61814:data<=16'd9592;
      61815:data<=16'd12480;
      61816:data<=16'd11571;
      61817:data<=16'd12160;
      61818:data<=16'd11872;
      61819:data<=16'd11662;
      61820:data<=16'd11976;
      61821:data<=16'd11461;
      61822:data<=16'd11655;
      61823:data<=16'd11452;
      61824:data<=16'd10390;
      61825:data<=16'd10522;
      61826:data<=16'd10561;
      61827:data<=16'd9859;
      61828:data<=16'd10358;
      61829:data<=16'd11614;
      61830:data<=16'd11676;
      61831:data<=16'd11082;
      61832:data<=16'd11015;
      61833:data<=16'd10496;
      61834:data<=16'd10014;
      61835:data<=16'd10360;
      61836:data<=16'd9946;
      61837:data<=16'd9646;
      61838:data<=16'd9737;
      61839:data<=16'd8704;
      61840:data<=16'd8734;
      61841:data<=16'd9950;
      61842:data<=16'd10298;
      61843:data<=16'd9973;
      61844:data<=16'd8843;
      61845:data<=16'd8987;
      61846:data<=16'd8593;
      61847:data<=16'd2467;
      61848:data<=-16'd2855;
      61849:data<=-16'd2376;
      61850:data<=-16'd2002;
      61851:data<=-16'd2179;
      61852:data<=-16'd1773;
      61853:data<=-16'd1817;
      61854:data<=-16'd429;
      61855:data<=16'd534;
      61856:data<=-16'd12;
      61857:data<=16'd309;
      61858:data<=16'd543;
      61859:data<=16'd588;
      61860:data<=16'd751;
      61861:data<=16'd321;
      61862:data<=16'd394;
      61863:data<=16'd262;
      61864:data<=-16'd62;
      61865:data<=16'd1078;
      61866:data<=16'd2469;
      61867:data<=16'd2857;
      61868:data<=16'd2323;
      61869:data<=16'd1947;
      61870:data<=16'd2249;
      61871:data<=16'd2167;
      61872:data<=16'd2391;
      61873:data<=16'd2197;
      61874:data<=16'd1421;
      61875:data<=16'd2373;
      61876:data<=16'd2437;
      61877:data<=16'd2058;
      61878:data<=16'd3645;
      61879:data<=16'd3259;
      61880:data<=16'd5709;
      61881:data<=16'd13835;
      61882:data<=16'd16070;
      61883:data<=16'd13292;
      61884:data<=16'd13389;
      61885:data<=16'd13189;
      61886:data<=16'd12502;
      61887:data<=16'd12683;
      61888:data<=16'd11969;
      61889:data<=16'd11649;
      61890:data<=16'd11612;
      61891:data<=16'd11585;
      61892:data<=16'd12111;
      61893:data<=16'd11773;
      61894:data<=16'd11133;
      61895:data<=16'd10850;
      61896:data<=16'd10504;
      61897:data<=16'd10194;
      61898:data<=16'd9300;
      61899:data<=16'd8777;
      61900:data<=16'd9033;
      61901:data<=16'd8478;
      61902:data<=16'd7665;
      61903:data<=16'd8179;
      61904:data<=16'd9709;
      61905:data<=16'd9788;
      61906:data<=16'd8520;
      61907:data<=16'd8405;
      61908:data<=16'd7959;
      61909:data<=16'd7151;
      61910:data<=16'd7112;
      61911:data<=16'd6178;
      61912:data<=16'd6701;
      61913:data<=16'd5943;
      61914:data<=-16'd1347;
      61915:data<=-16'd6223;
      61916:data<=-16'd4611;
      61917:data<=-16'd3688;
      61918:data<=-16'd3391;
      61919:data<=-16'd3046;
      61920:data<=-16'd3601;
      61921:data<=-16'd3400;
      61922:data<=-16'd3568;
      61923:data<=-16'd3776;
      61924:data<=-16'd3338;
      61925:data<=-16'd3313;
      61926:data<=-16'd2939;
      61927:data<=-16'd3119;
      61928:data<=-16'd3212;
      61929:data<=-16'd1955;
      61930:data<=-16'd1726;
      61931:data<=-16'd1660;
      61932:data<=-16'd1078;
      61933:data<=-16'd1378;
      61934:data<=-16'd1439;
      61935:data<=-16'd1692;
      61936:data<=-16'd1838;
      61937:data<=-16'd1583;
      61938:data<=-16'd2270;
      61939:data<=-16'd2000;
      61940:data<=-16'd1648;
      61941:data<=-16'd1651;
      61942:data<=16'd85;
      61943:data<=16'd153;
      61944:data<=16'd99;
      61945:data<=16'd1104;
      61946:data<=-16'd1077;
      61947:data<=16'd1898;
      61948:data<=16'd10531;
      61949:data<=16'd11329;
      61950:data<=16'd9060;
      61951:data<=16'd10114;
      61952:data<=16'd9050;
      61953:data<=16'd8370;
      61954:data<=16'd9582;
      61955:data<=16'd9576;
      61956:data<=16'd9600;
      61957:data<=16'd9333;
      61958:data<=16'd8420;
      61959:data<=16'd7943;
      61960:data<=16'd7685;
      61961:data<=16'd7580;
      61962:data<=16'd6927;
      61963:data<=16'd6496;
      61964:data<=16'd6539;
      61965:data<=16'd5656;
      61966:data<=16'd5847;
      61967:data<=16'd6971;
      61968:data<=16'd6417;
      61969:data<=16'd5909;
      61970:data<=16'd6299;
      61971:data<=16'd6008;
      61972:data<=16'd5250;
      61973:data<=16'd4981;
      61974:data<=16'd4837;
      61975:data<=16'd4147;
      61976:data<=16'd4023;
      61977:data<=16'd3591;
      61978:data<=16'd2675;
      61979:data<=16'd4773;
      61980:data<=16'd4532;
      61981:data<=-16'd2864;
      61982:data<=-16'd7397;
      61983:data<=-16'd6247;
      61984:data<=-16'd6504;
      61985:data<=-16'd6833;
      61986:data<=-16'd5976;
      61987:data<=-16'd6223;
      61988:data<=-16'd6331;
      61989:data<=-16'd5976;
      61990:data<=-16'd5830;
      61991:data<=-16'd5280;
      61992:data<=-16'd4340;
      61993:data<=-16'd3751;
      61994:data<=-16'd3853;
      61995:data<=-16'd3876;
      61996:data<=-16'd3835;
      61997:data<=-16'd3997;
      61998:data<=-16'd3993;
      61999:data<=-16'd4258;
      62000:data<=-16'd3971;
      62001:data<=-16'd3460;
      62002:data<=-16'd4200;
      62003:data<=-16'd4288;
      62004:data<=-16'd4143;
      62005:data<=-16'd4699;
      62006:data<=-16'd3818;
      62007:data<=-16'd3709;
      62008:data<=-16'd4482;
      62009:data<=-16'd3820;
      62010:data<=-16'd4393;
      62011:data<=-16'd4070;
      62012:data<=-16'd2748;
      62013:data<=-16'd5056;
      62014:data<=-16'd2537;
      62015:data<=16'd6435;
      62016:data<=16'd7694;
      62017:data<=16'd3645;
      62018:data<=16'd3682;
      62019:data<=16'd3689;
      62020:data<=16'd2679;
      62021:data<=16'd2966;
      62022:data<=16'd2387;
      62023:data<=16'd1989;
      62024:data<=16'd2507;
      62025:data<=16'd2040;
      62026:data<=16'd1739;
      62027:data<=16'd1845;
      62028:data<=16'd793;
      62029:data<=-16'd547;
      62030:data<=-16'd1236;
      62031:data<=-16'd1457;
      62032:data<=-16'd1448;
      62033:data<=-16'd1545;
      62034:data<=-16'd1400;
      62035:data<=-16'd1707;
      62036:data<=-16'd2761;
      62037:data<=-16'd2312;
      62038:data<=-16'd1533;
      62039:data<=-16'd2364;
      62040:data<=-16'd2278;
      62041:data<=-16'd2614;
      62042:data<=-16'd4787;
      62043:data<=-16'd4807;
      62044:data<=-16'd4593;
      62045:data<=-16'd5682;
      62046:data<=-16'd4203;
      62047:data<=-16'd5448;
      62048:data<=-16'd12301;
      62049:data<=-16'd15564;
      62050:data<=-16'd14422;
      62051:data<=-16'd14204;
      62052:data<=-16'd13734;
      62053:data<=-16'd13345;
      62054:data<=-16'd14442;
      62055:data<=-16'd14918;
      62056:data<=-16'd14307;
      62057:data<=-16'd13858;
      62058:data<=-16'd13694;
      62059:data<=-16'd13245;
      62060:data<=-16'd12747;
      62061:data<=-16'd12522;
      62062:data<=-16'd11723;
      62063:data<=-16'd11041;
      62064:data<=-16'd10994;
      62065:data<=-16'd10398;
      62066:data<=-16'd10551;
      62067:data<=-16'd11333;
      62068:data<=-16'd10906;
      62069:data<=-16'd10968;
      62070:data<=-16'd11162;
      62071:data<=-16'd10248;
      62072:data<=-16'd10034;
      62073:data<=-16'd9773;
      62074:data<=-16'd9186;
      62075:data<=-16'd9019;
      62076:data<=-16'd8220;
      62077:data<=-16'd8126;
      62078:data<=-16'd7928;
      62079:data<=-16'd7743;
      62080:data<=-16'd10314;
      62081:data<=-16'd7635;
      62082:data<=16'd1680;
      62083:data<=16'd4035;
      62084:data<=16'd1380;
      62085:data<=16'd1989;
      62086:data<=16'd2168;
      62087:data<=16'd2261;
      62088:data<=16'd2722;
      62089:data<=16'd1612;
      62090:data<=16'd2346;
      62091:data<=16'd2449;
      62092:data<=-16'd32;
      62093:data<=-16'd240;
      62094:data<=16'd152;
      62095:data<=-16'd331;
      62096:data<=16'd320;
      62097:data<=16'd23;
      62098:data<=-16'd585;
      62099:data<=-16'd135;
      62100:data<=-16'd290;
      62101:data<=-16'd152;
      62102:data<=16'd162;
      62103:data<=-16'd547;
      62104:data<=-16'd1162;
      62105:data<=-16'd1747;
      62106:data<=-16'd2247;
      62107:data<=-16'd1926;
      62108:data<=-16'd1809;
      62109:data<=-16'd1715;
      62110:data<=-16'd1064;
      62111:data<=-16'd1592;
      62112:data<=-16'd2265;
      62113:data<=-16'd763;
      62114:data<=-16'd1889;
      62115:data<=-16'd8483;
      62116:data<=-16'd13207;
      62117:data<=-16'd13397;
      62118:data<=-16'd13180;
      62119:data<=-16'd12569;
      62120:data<=-16'd11729;
      62121:data<=-16'd11586;
      62122:data<=-16'd11022;
      62123:data<=-16'd10728;
      62124:data<=-16'd10543;
      62125:data<=-16'd9682;
      62126:data<=-16'd9083;
      62127:data<=-16'd8578;
      62128:data<=-16'd8299;
      62129:data<=-16'd8278;
      62130:data<=-16'd8291;
      62131:data<=-16'd8887;
      62132:data<=-16'd8605;
      62133:data<=-16'd7650;
      62134:data<=-16'd7473;
      62135:data<=-16'd7110;
      62136:data<=-16'd7087;
      62137:data<=-16'd7006;
      62138:data<=-16'd6375;
      62139:data<=-16'd6394;
      62140:data<=-16'd5379;
      62141:data<=-16'd5207;
      62142:data<=-16'd7025;
      62143:data<=-16'd6407;
      62144:data<=-16'd5691;
      62145:data<=-16'd5538;
      62146:data<=-16'd4193;
      62147:data<=-16'd5744;
      62148:data<=-16'd3142;
      62149:data<=16'd6266;
      62150:data<=16'd8478;
      62151:data<=16'd5882;
      62152:data<=16'd6880;
      62153:data<=16'd6713;
      62154:data<=16'd5811;
      62155:data<=16'd5316;
      62156:data<=16'd4061;
      62157:data<=16'd4863;
      62158:data<=16'd5380;
      62159:data<=16'd4316;
      62160:data<=16'd4261;
      62161:data<=16'd4235;
      62162:data<=16'd4291;
      62163:data<=16'd4193;
      62164:data<=16'd3604;
      62165:data<=16'd4131;
      62166:data<=16'd4134;
      62167:data<=16'd3058;
      62168:data<=16'd2584;
      62169:data<=16'd2458;
      62170:data<=16'd2420;
      62171:data<=16'd2206;
      62172:data<=16'd2622;
      62173:data<=16'd3372;
      62174:data<=16'd2745;
      62175:data<=16'd2535;
      62176:data<=16'd2728;
      62177:data<=16'd2247;
      62178:data<=16'd2443;
      62179:data<=16'd2012;
      62180:data<=16'd1474;
      62181:data<=-16'd182;
      62182:data<=-16'd6343;
      62183:data<=-16'd10220;
      62184:data<=-16'd8745;
      62185:data<=-16'd8715;
      62186:data<=-16'd8860;
      62187:data<=-16'd7413;
      62188:data<=-16'd7429;
      62189:data<=-16'd7470;
      62190:data<=-16'd6939;
      62191:data<=-16'd7306;
      62192:data<=-16'd7644;
      62193:data<=-16'd6965;
      62194:data<=-16'd6325;
      62195:data<=-16'd6523;
      62196:data<=-16'd5570;
      62197:data<=-16'd4335;
      62198:data<=-16'd4748;
      62199:data<=-16'd4400;
      62200:data<=-16'd4052;
      62201:data<=-16'd4290;
      62202:data<=-16'd3310;
      62203:data<=-16'd3330;
      62204:data<=-16'd3130;
      62205:data<=-16'd2059;
      62206:data<=-16'd2787;
      62207:data<=-16'd2111;
      62208:data<=-16'd1272;
      62209:data<=-16'd2408;
      62210:data<=-16'd1491;
      62211:data<=-16'd1005;
      62212:data<=-16'd699;
      62213:data<=16'd825;
      62214:data<=-16'd1163;
      62215:data<=16'd1149;
      62216:data<=16'd10379;
      62217:data<=16'd13473;
      62218:data<=16'd12289;
      62219:data<=16'd12919;
      62220:data<=16'd12372;
      62221:data<=16'd12149;
      62222:data<=16'd12192;
      62223:data<=16'd11737;
      62224:data<=16'd12182;
      62225:data<=16'd11162;
      62226:data<=16'd10281;
      62227:data<=16'd10991;
      62228:data<=16'd10113;
      62229:data<=16'd9697;
      62230:data<=16'd11115;
      62231:data<=16'd11262;
      62232:data<=16'd10657;
      62233:data<=16'd10927;
      62234:data<=16'd10777;
      62235:data<=16'd9979;
      62236:data<=16'd10043;
      62237:data<=16'd9641;
      62238:data<=16'd8511;
      62239:data<=16'd9295;
      62240:data<=16'd9676;
      62241:data<=16'd8868;
      62242:data<=16'd10122;
      62243:data<=16'd11036;
      62244:data<=16'd10592;
      62245:data<=16'd10064;
      62246:data<=16'd9025;
      62247:data<=16'd9755;
      62248:data<=16'd7943;
      62249:data<=16'd432;
      62250:data<=-16'd3234;
      62251:data<=-16'd2200;
      62252:data<=-16'd2591;
      62253:data<=-16'd2250;
      62254:data<=-16'd778;
      62255:data<=16'd337;
      62256:data<=16'd857;
      62257:data<=16'd234;
      62258:data<=16'd500;
      62259:data<=16'd960;
      62260:data<=16'd778;
      62261:data<=16'd1380;
      62262:data<=16'd911;
      62263:data<=16'd675;
      62264:data<=16'd1917;
      62265:data<=16'd1451;
      62266:data<=16'd1057;
      62267:data<=16'd2428;
      62268:data<=16'd3456;
      62269:data<=16'd3506;
      62270:data<=16'd2793;
      62271:data<=16'd3065;
      62272:data<=16'd3339;
      62273:data<=16'd2234;
      62274:data<=16'd2790;
      62275:data<=16'd3287;
      62276:data<=16'd2584;
      62277:data<=16'd2963;
      62278:data<=16'd2082;
      62279:data<=16'd2617;
      62280:data<=16'd4928;
      62281:data<=16'd3259;
      62282:data<=16'd5861;
      62283:data<=16'd14804;
      62284:data<=16'd16154;
      62285:data<=16'd12883;
      62286:data<=16'd13712;
      62287:data<=16'd13614;
      62288:data<=16'd11958;
      62289:data<=16'd11991;
      62290:data<=16'd11822;
      62291:data<=16'd11414;
      62292:data<=16'd12129;
      62293:data<=16'd12766;
      62294:data<=16'd12193;
      62295:data<=16'd11209;
      62296:data<=16'd10513;
      62297:data<=16'd9964;
      62298:data<=16'd9856;
      62299:data<=16'd9814;
      62300:data<=16'd9485;
      62301:data<=16'd9128;
      62302:data<=16'd8238;
      62303:data<=16'd7353;
      62304:data<=16'd7588;
      62305:data<=16'd8825;
      62306:data<=16'd9679;
      62307:data<=16'd8672;
      62308:data<=16'd7589;
      62309:data<=16'd7335;
      62310:data<=16'd6689;
      62311:data<=16'd7297;
      62312:data<=16'd7141;
      62313:data<=16'd5216;
      62314:data<=16'd6375;
      62315:data<=16'd4716;
      62316:data<=-16'd3409;
      62317:data<=-16'd5927;
      62318:data<=-16'd3078;
      62319:data<=-16'd3532;
      62320:data<=-16'd3905;
      62321:data<=-16'd3278;
      62322:data<=-16'd3853;
      62323:data<=-16'd3612;
      62324:data<=-16'd3579;
      62325:data<=-16'd3789;
      62326:data<=-16'd3025;
      62327:data<=-16'd3204;
      62328:data<=-16'd3798;
      62329:data<=-16'd2980;
      62330:data<=-16'd1441;
      62331:data<=-16'd845;
      62332:data<=-16'd1548;
      62333:data<=-16'd2008;
      62334:data<=-16'd1983;
      62335:data<=-16'd1381;
      62336:data<=-16'd364;
      62337:data<=-16'd1122;
      62338:data<=-16'd1865;
      62339:data<=-16'd1162;
      62340:data<=-16'd1798;
      62341:data<=-16'd2032;
      62342:data<=-16'd755;
      62343:data<=-16'd355;
      62344:data<=-16'd165;
      62345:data<=-16'd464;
      62346:data<=-16'd541;
      62347:data<=16'd9;
      62348:data<=-16'd1213;
      62349:data<=16'd1741;
      62350:data<=16'd9949;
      62351:data<=16'd11580;
      62352:data<=16'd8193;
      62353:data<=16'd8244;
      62354:data<=16'd8857;
      62355:data<=16'd8919;
      62356:data<=16'd9379;
      62357:data<=16'd8721;
      62358:data<=16'd8385;
      62359:data<=16'd8231;
      62360:data<=16'd7556;
      62361:data<=16'd7277;
      62362:data<=16'd6219;
      62363:data<=16'd5116;
      62364:data<=16'd5190;
      62365:data<=16'd4827;
      62366:data<=16'd4467;
      62367:data<=16'd5124;
      62368:data<=16'd5436;
      62369:data<=16'd4908;
      62370:data<=16'd4491;
      62371:data<=16'd4212;
      62372:data<=16'd3758;
      62373:data<=16'd3610;
      62374:data<=16'd3280;
      62375:data<=16'd2554;
      62376:data<=16'd2328;
      62377:data<=16'd2246;
      62378:data<=16'd2563;
      62379:data<=16'd2658;
      62380:data<=16'd2152;
      62381:data<=16'd3416;
      62382:data<=16'd1413;
      62383:data<=-16'd6593;
      62384:data<=-16'd9712;
      62385:data<=-16'd7739;
      62386:data<=-16'd8464;
      62387:data<=-16'd8413;
      62388:data<=-16'd7385;
      62389:data<=-16'd7556;
      62390:data<=-16'd7265;
      62391:data<=-16'd8589;
      62392:data<=-16'd8282;
      62393:data<=-16'd4834;
      62394:data<=-16'd4848;
      62395:data<=-16'd5805;
      62396:data<=-16'd4699;
      62397:data<=-16'd4701;
      62398:data<=-16'd4388;
      62399:data<=-16'd4118;
      62400:data<=-16'd4787;
      62401:data<=-16'd4602;
      62402:data<=-16'd4673;
      62403:data<=-16'd4714;
      62404:data<=-16'd4616;
      62405:data<=-16'd5127;
      62406:data<=-16'd4810;
      62407:data<=-16'd4575;
      62408:data<=-16'd4493;
      62409:data<=-16'd4153;
      62410:data<=-16'd4613;
      62411:data<=-16'd4394;
      62412:data<=-16'd4288;
      62413:data<=-16'd4087;
      62414:data<=-16'd3160;
      62415:data<=-16'd4543;
      62416:data<=-16'd1894;
      62417:data<=16'd5635;
      62418:data<=16'd5691;
      62419:data<=16'd2731;
      62420:data<=16'd3918;
      62421:data<=16'd3203;
      62422:data<=16'd2399;
      62423:data<=16'd2622;
      62424:data<=16'd1647;
      62425:data<=16'd2834;
      62426:data<=16'd2845;
      62427:data<=16'd846;
      62428:data<=16'd1395;
      62429:data<=16'd643;
      62430:data<=-16'd1563;
      62431:data<=-16'd1571;
      62432:data<=-16'd1754;
      62433:data<=-16'd2165;
      62434:data<=-16'd1659;
      62435:data<=-16'd1333;
      62436:data<=-16'd1363;
      62437:data<=-16'd1926;
      62438:data<=-16'd2444;
      62439:data<=-16'd2654;
      62440:data<=-16'd2881;
      62441:data<=-16'd2807;
      62442:data<=-16'd3254;
      62443:data<=-16'd4384;
      62444:data<=-16'd4860;
      62445:data<=-16'd4484;
      62446:data<=-16'd4868;
      62447:data<=-16'd5471;
      62448:data<=-16'd4021;
      62449:data<=-16'd5858;
      62450:data<=-16'd13288;
      62451:data<=-16'd16177;
      62452:data<=-16'd14195;
      62453:data<=-16'd14099;
      62454:data<=-16'd13514;
      62455:data<=-16'd13376;
      62456:data<=-16'd14642;
      62457:data<=-16'd14069;
      62458:data<=-16'd14273;
      62459:data<=-16'd14292;
      62460:data<=-16'd12111;
      62461:data<=-16'd11729;
      62462:data<=-16'd11787;
      62463:data<=-16'd11036;
      62464:data<=-16'd11496;
      62465:data<=-16'd10884;
      62466:data<=-16'd9706;
      62467:data<=-16'd10580;
      62468:data<=-16'd11555;
      62469:data<=-16'd10551;
      62470:data<=-16'd9232;
      62471:data<=-16'd9526;
      62472:data<=-16'd9386;
      62473:data<=-16'd8640;
      62474:data<=-16'd8872;
      62475:data<=-16'd7932;
      62476:data<=-16'd7476;
      62477:data<=-16'd8311;
      62478:data<=-16'd6974;
      62479:data<=-16'd6346;
      62480:data<=-16'd6734;
      62481:data<=-16'd6341;
      62482:data<=-16'd7241;
      62483:data<=-16'd3585;
      62484:data<=16'd3703;
      62485:data<=16'd4451;
      62486:data<=16'd3098;
      62487:data<=16'd3993;
      62488:data<=16'd3570;
      62489:data<=16'd3577;
      62490:data<=16'd3397;
      62491:data<=16'd2964;
      62492:data<=16'd3824;
      62493:data<=16'd1950;
      62494:data<=-16'd91;
      62495:data<=16'd1430;
      62496:data<=16'd1369;
      62497:data<=-16'd71;
      62498:data<=16'd572;
      62499:data<=16'd743;
      62500:data<=-16'd138;
      62501:data<=-16'd18;
      62502:data<=16'd6;
      62503:data<=-16'd44;
      62504:data<=16'd1149;
      62505:data<=16'd282;
      62506:data<=-16'd2591;
      62507:data<=-16'd2319;
      62508:data<=-16'd1001;
      62509:data<=-16'd993;
      62510:data<=-16'd666;
      62511:data<=-16'd1394;
      62512:data<=-16'd1224;
      62513:data<=-16'd391;
      62514:data<=-16'd1433;
      62515:data<=-16'd26;
      62516:data<=-16'd1316;
      62517:data<=-16'd9568;
      62518:data<=-16'd12548;
      62519:data<=-16'd10665;
      62520:data<=-16'd11599;
      62521:data<=-16'd10898;
      62522:data<=-16'd9693;
      62523:data<=-16'd10372;
      62524:data<=-16'd9643;
      62525:data<=-16'd8590;
      62526:data<=-16'd7830;
      62527:data<=-16'd7659;
      62528:data<=-16'd7780;
      62529:data<=-16'd6149;
      62530:data<=-16'd6135;
      62531:data<=-16'd7739;
      62532:data<=-16'd7069;
      62533:data<=-16'd6202;
      62534:data<=-16'd5759;
      62535:data<=-16'd4948;
      62536:data<=-16'd4939;
      62537:data<=-16'd5036;
      62538:data<=-16'd5206;
      62539:data<=-16'd5074;
      62540:data<=-16'd4015;
      62541:data<=-16'd2975;
      62542:data<=-16'd2798;
      62543:data<=-16'd4936;
      62544:data<=-16'd6649;
      62545:data<=-16'd5298;
      62546:data<=-16'd4780;
      62547:data<=-16'd4420;
      62548:data<=-16'd3298;
      62549:data<=-16'd3814;
      62550:data<=-16'd105;
      62551:data<=16'd7409;
      62552:data<=16'd8813;
      62553:data<=16'd6757;
      62554:data<=16'd7397;
      62555:data<=16'd7376;
      62556:data<=16'd5513;
      62557:data<=16'd5148;
      62558:data<=16'd6125;
      62559:data<=16'd6072;
      62560:data<=16'd5157;
      62561:data<=16'd4414;
      62562:data<=16'd4698;
      62563:data<=16'd5739;
      62564:data<=16'd4851;
      62565:data<=16'd3805;
      62566:data<=16'd4751;
      62567:data<=16'd4027;
      62568:data<=16'd3127;
      62569:data<=16'd3585;
      62570:data<=16'd2334;
      62571:data<=16'd2372;
      62572:data<=16'd3319;
      62573:data<=16'd2305;
      62574:data<=16'd3075;
      62575:data<=16'd3735;
      62576:data<=16'd2403;
      62577:data<=16'd2322;
      62578:data<=16'd2540;
      62579:data<=16'd3436;
      62580:data<=16'd2880;
      62581:data<=-16'd92;
      62582:data<=16'd1249;
      62583:data<=16'd525;
      62584:data<=-16'd7688;
      62585:data<=-16'd10489;
      62586:data<=-16'd7562;
      62587:data<=-16'd7829;
      62588:data<=-16'd8194;
      62589:data<=-16'd6771;
      62590:data<=-16'd5776;
      62591:data<=-16'd5815;
      62592:data<=-16'd6531;
      62593:data<=-16'd6786;
      62594:data<=-16'd7216;
      62595:data<=-16'd6784;
      62596:data<=-16'd5400;
      62597:data<=-16'd5570;
      62598:data<=-16'd5048;
      62599:data<=-16'd4058;
      62600:data<=-16'd4743;
      62601:data<=-16'd3947;
      62602:data<=-16'd2804;
      62603:data<=-16'd3057;
      62604:data<=-16'd2343;
      62605:data<=-16'd1965;
      62606:data<=-16'd2087;
      62607:data<=-16'd1885;
      62608:data<=-16'd2276;
      62609:data<=-16'd1322;
      62610:data<=-16'd167;
      62611:data<=-16'd1306;
      62612:data<=-16'd2026;
      62613:data<=-16'd1249;
      62614:data<=-16'd667;
      62615:data<=-16'd641;
      62616:data<=16'd757;
      62617:data<=16'd5887;
      62618:data<=16'd11844;
      62619:data<=16'd13964;
      62620:data<=16'd12742;
      62621:data<=16'd11421;
      62622:data<=16'd11309;
      62623:data<=16'd10994;
      62624:data<=16'd10513;
      62625:data<=16'd10618;
      62626:data<=16'd10096;
      62627:data<=16'd9755;
      62628:data<=16'd9934;
      62629:data<=16'd9498;
      62630:data<=16'd9693;
      62631:data<=16'd10003;
      62632:data<=16'd9940;
      62633:data<=16'd10217;
      62634:data<=16'd9263;
      62635:data<=16'd8678;
      62636:data<=16'd9276;
      62637:data<=16'd8692;
      62638:data<=16'd8874;
      62639:data<=16'd9069;
      62640:data<=16'd7382;
      62641:data<=16'd7109;
      62642:data<=16'd7703;
      62643:data<=16'd8204;
      62644:data<=16'd8840;
      62645:data<=16'd7585;
      62646:data<=16'd7632;
      62647:data<=16'd8874;
      62648:data<=16'd8276;
      62649:data<=16'd9336;
      62650:data<=16'd6778;
      62651:data<=-16'd2014;
      62652:data<=-16'd4118;
      62653:data<=-16'd1243;
      62654:data<=-16'd2537;
      62655:data<=-16'd2309;
      62656:data<=-16'd39;
      62657:data<=-16'd147;
      62658:data<=-16'd71;
      62659:data<=16'd91;
      62660:data<=-16'd484;
      62661:data<=-16'd503;
      62662:data<=16'd26;
      62663:data<=16'd1130;
      62664:data<=16'd604;
      62665:data<=-16'd890;
      62666:data<=16'd352;
      62667:data<=16'd1148;
      62668:data<=16'd384;
      62669:data<=16'd2118;
      62670:data<=16'd3577;
      62671:data<=16'd2585;
      62672:data<=16'd2487;
      62673:data<=16'd2817;
      62674:data<=16'd2261;
      62675:data<=16'd2009;
      62676:data<=16'd2021;
      62677:data<=16'd2033;
      62678:data<=16'd1935;
      62679:data<=16'd1706;
      62680:data<=16'd2532;
      62681:data<=16'd4067;
      62682:data<=16'd4137;
      62683:data<=16'd4141;
      62684:data<=16'd8052;
      62685:data<=16'd13295;
      62686:data<=16'd14010;
      62687:data<=16'd12354;
      62688:data<=16'd11852;
      62689:data<=16'd10736;
      62690:data<=16'd9679;
      62691:data<=16'd9561;
      62692:data<=16'd8913;
      62693:data<=16'd9594;
      62694:data<=16'd11207;
      62695:data<=16'd10895;
      62696:data<=16'd10724;
      62697:data<=16'd10781;
      62698:data<=16'd9054;
      62699:data<=16'd8420;
      62700:data<=16'd8755;
      62701:data<=16'd7157;
      62702:data<=16'd6214;
      62703:data<=16'd6924;
      62704:data<=16'd6771;
      62705:data<=16'd7148;
      62706:data<=16'd8994;
      62707:data<=16'd9345;
      62708:data<=16'd7744;
      62709:data<=16'd7316;
      62710:data<=16'd8281;
      62711:data<=16'd7272;
      62712:data<=16'd5680;
      62713:data<=16'd6614;
      62714:data<=16'd6379;
      62715:data<=16'd5139;
      62716:data<=16'd6331;
      62717:data<=16'd3791;
      62718:data<=-16'd2079;
      62719:data<=-16'd2516;
      62720:data<=-16'd1792;
      62721:data<=-16'd3134;
      62722:data<=-16'd1759;
      62723:data<=-16'd1333;
      62724:data<=-16'd2505;
      62725:data<=-16'd1248;
      62726:data<=-16'd1562;
      62727:data<=-16'd3283;
      62728:data<=-16'd2667;
      62729:data<=-16'd2294;
      62730:data<=-16'd2560;
      62731:data<=-16'd1815;
      62732:data<=-16'd857;
      62733:data<=-16'd208;
      62734:data<=16'd190;
      62735:data<=16'd817;
      62736:data<=16'd505;
      62737:data<=-16'd1118;
      62738:data<=-16'd1554;
      62739:data<=-16'd1371;
      62740:data<=-16'd1257;
      62741:data<=-16'd564;
      62742:data<=-16'd1192;
      62743:data<=-16'd1902;
      62744:data<=-16'd810;
      62745:data<=-16'd144;
      62746:data<=-16'd56;
      62747:data<=16'd305;
      62748:data<=16'd238;
      62749:data<=-16'd382;
      62750:data<=16'd83;
      62751:data<=16'd4081;
      62752:data<=16'd8434;
      62753:data<=16'd9015;
      62754:data<=16'd8490;
      62755:data<=16'd8439;
      62756:data<=16'd8743;
      62757:data<=16'd9606;
      62758:data<=16'd8481;
      62759:data<=16'd7013;
      62760:data<=16'd7495;
      62761:data<=16'd6705;
      62762:data<=16'd5568;
      62763:data<=16'd7009;
      62764:data<=16'd8088;
      62765:data<=16'd5976;
      62766:data<=16'd3356;
      62767:data<=16'd3671;
      62768:data<=16'd4570;
      62769:data<=16'd4508;
      62770:data<=16'd5993;
      62771:data<=16'd6408;
      62772:data<=16'd4590;
      62773:data<=16'd4731;
      62774:data<=16'd5089;
      62775:data<=16'd3482;
      62776:data<=16'd3222;
      62777:data<=16'd4381;
      62778:data<=16'd3638;
      62779:data<=16'd1771;
      62780:data<=16'd2432;
      62781:data<=16'd3486;
      62782:data<=16'd2526;
      62783:data<=16'd3107;
      62784:data<=16'd1550;
      62785:data<=-16'd5597;
      62786:data<=-16'd9301;
      62787:data<=-16'd7931;
      62788:data<=-16'd7680;
      62789:data<=-16'd7827;
      62790:data<=-16'd7558;
      62791:data<=-16'd7069;
      62792:data<=-16'd6652;
      62793:data<=-16'd7401;
      62794:data<=-16'd6344;
      62795:data<=-16'd4068;
      62796:data<=-16'd4393;
      62797:data<=-16'd5495;
      62798:data<=-16'd6260;
      62799:data<=-16'd6834;
      62800:data<=-16'd5890;
      62801:data<=-16'd4831;
      62802:data<=-16'd5015;
      62803:data<=-16'd5483;
      62804:data<=-16'd4821;
      62805:data<=-16'd3955;
      62806:data<=-16'd5062;
      62807:data<=-16'd5589;
      62808:data<=-16'd4378;
      62809:data<=-16'd4848;
      62810:data<=-16'd5871;
      62811:data<=-16'd5168;
      62812:data<=-16'd4309;
      62813:data<=-16'd4861;
      62814:data<=-16'd5774;
      62815:data<=-16'd4896;
      62816:data<=-16'd6238;
      62817:data<=-16'd12366;
      62818:data<=-16'd14744;
      62819:data<=-16'd11321;
      62820:data<=-16'd9721;
      62821:data<=-16'd10756;
      62822:data<=-16'd11236;
      62823:data<=-16'd10167;
      62824:data<=-16'd9110;
      62825:data<=-16'd10070;
      62826:data<=-16'd10470;
      62827:data<=-16'd9532;
      62828:data<=-16'd10006;
      62829:data<=-16'd10443;
      62830:data<=-16'd9163;
      62831:data<=-16'd8220;
      62832:data<=-16'd9153;
      62833:data<=-16'd9987;
      62834:data<=-16'd8398;
      62835:data<=-16'd5953;
      62836:data<=-16'd4111;
      62837:data<=-16'd4120;
      62838:data<=-16'd6637;
      62839:data<=-16'd7181;
      62840:data<=-16'd6534;
      62841:data<=-16'd8011;
      62842:data<=-16'd6865;
      62843:data<=-16'd4805;
      62844:data<=-16'd5112;
      62845:data<=-16'd3858;
      62846:data<=-16'd4634;
      62847:data<=-16'd4429;
      62848:data<=16'd4278;
      62849:data<=16'd7401;
      62850:data<=-16'd1647;
      62851:data<=-16'd10730;
      62852:data<=-16'd18346;
      62853:data<=-16'd21466;
      62854:data<=-16'd15875;
      62855:data<=-16'd12000;
      62856:data<=-16'd11791;
      62857:data<=-16'd11972;
      62858:data<=-16'd16351;
      62859:data<=-16'd16110;
      62860:data<=-16'd9166;
      62861:data<=-16'd11929;
      62862:data<=-16'd17829;
      62863:data<=-16'd11617;
      62864:data<=-16'd6623;
      62865:data<=-16'd10481;
      62866:data<=-16'd10746;
      62867:data<=-16'd6466;
      62868:data<=-16'd3259;
      62869:data<=-16'd2170;
      62870:data<=-16'd6109;
      62871:data<=-16'd13089;
      62872:data<=-16'd16768;
      62873:data<=-16'd14657;
      62874:data<=-16'd9218;
      62875:data<=-16'd6021;
      62876:data<=-16'd6419;
      62877:data<=-16'd10348;
      62878:data<=-16'd14316;
      62879:data<=-16'd8316;
      62880:data<=-16'd2134;
      62881:data<=-16'd8752;
      62882:data<=-16'd10924;
      62883:data<=-16'd4278;
      62884:data<=-16'd1092;
      62885:data<=16'd6097;
      62886:data<=16'd11471;
      62887:data<=16'd4608;
      62888:data<=16'd3586;
      62889:data<=16'd10019;
      62890:data<=16'd6488;
      62891:data<=-16'd3198;
      62892:data<=-16'd6270;
      62893:data<=-16'd2419;
      62894:data<=-16'd2074;
      62895:data<=-16'd3140;
      62896:data<=16'd3388;
      62897:data<=16'd4502;
      62898:data<=-16'd1177;
      62899:data<=16'd338;
      62900:data<=16'd946;
      62901:data<=16'd1468;
      62902:data<=16'd5956;
      62903:data<=16'd466;
      62904:data<=-16'd5347;
      62905:data<=-16'd2434;
      62906:data<=-16'd1879;
      62907:data<=-16'd23;
      62908:data<=16'd1157;
      62909:data<=16'd1256;
      62910:data<=16'd6751;
      62911:data<=16'd444;
      62912:data<=-16'd9177;
      62913:data<=-16'd690;
      62914:data<=16'd3136;
      62915:data<=-16'd146;
      62916:data<=16'd3773;
      62917:data<=-16'd596;
      62918:data<=-16'd6091;
      62919:data<=-16'd3096;
      62920:data<=-16'd6983;
      62921:data<=-16'd8117;
      62922:data<=-16'd2008;
      62923:data<=-16'd6780;
      62924:data<=-16'd13576;
      62925:data<=-16'd9291;
      62926:data<=-16'd5879;
      62927:data<=-16'd9627;
      62928:data<=-16'd9841;
      62929:data<=-16'd4880;
      62930:data<=-16'd7056;
      62931:data<=-16'd13408;
      62932:data<=-16'd13022;
      62933:data<=-16'd9360;
      62934:data<=-16'd4206;
      62935:data<=-16'd2453;
      62936:data<=-16'd8869;
      62937:data<=-16'd9144;
      62938:data<=-16'd6067;
      62939:data<=-16'd12880;
      62940:data<=-16'd13494;
      62941:data<=-16'd3845;
      62942:data<=-16'd361;
      62943:data<=-16'd2276;
      62944:data<=-16'd4655;
      62945:data<=-16'd3438;
      62946:data<=16'd528;
      62947:data<=-16'd1823;
      62948:data<=-16'd813;
      62949:data<=16'd4969;
      62950:data<=16'd688;
      62951:data<=16'd1842;
      62952:data<=16'd12605;
      62953:data<=16'd12342;
      62954:data<=16'd13876;
      62955:data<=16'd21140;
      62956:data<=16'd15618;
      62957:data<=16'd9746;
      62958:data<=16'd8619;
      62959:data<=16'd5682;
      62960:data<=16'd12184;
      62961:data<=16'd16149;
      62962:data<=16'd10563;
      62963:data<=16'd15138;
      62964:data<=16'd19064;
      62965:data<=16'd15109;
      62966:data<=16'd17653;
      62967:data<=16'd15898;
      62968:data<=16'd12041;
      62969:data<=16'd18445;
      62970:data<=16'd17399;
      62971:data<=16'd10249;
      62972:data<=16'd11715;
      62973:data<=16'd12977;
      62974:data<=16'd13697;
      62975:data<=16'd15928;
      62976:data<=16'd14041;
      62977:data<=16'd13288;
      62978:data<=16'd11770;
      62979:data<=16'd8006;
      62980:data<=16'd13160;
      62981:data<=16'd20854;
      62982:data<=16'd18575;
      62983:data<=16'd13931;
      62984:data<=16'd13543;
      62985:data<=16'd9970;
      62986:data<=16'd2174;
      62987:data<=16'd1154;
      62988:data<=16'd4977;
      62989:data<=16'd3610;
      62990:data<=16'd3341;
      62991:data<=16'd6737;
      62992:data<=16'd6363;
      62993:data<=16'd5714;
      62994:data<=16'd7227;
      62995:data<=16'd7535;
      62996:data<=16'd6622;
      62997:data<=16'd5159;
      62998:data<=16'd5104;
      62999:data<=16'd3294;
      63000:data<=16'd775;
      63001:data<=16'd6129;
      63002:data<=16'd9085;
      63003:data<=16'd3982;
      63004:data<=16'd4942;
      63005:data<=16'd7185;
      63006:data<=16'd4975;
      63007:data<=16'd7454;
      63008:data<=16'd10179;
      63009:data<=16'd9461;
      63010:data<=16'd8994;
      63011:data<=16'd6760;
      63012:data<=16'd3039;
      63013:data<=-16'd79;
      63014:data<=16'd3046;
      63015:data<=16'd9909;
      63016:data<=16'd8824;
      63017:data<=16'd10375;
      63018:data<=16'd18783;
      63019:data<=16'd18589;
      63020:data<=16'd18906;
      63021:data<=16'd22883;
      63022:data<=16'd16424;
      63023:data<=16'd11019;
      63024:data<=16'd12833;
      63025:data<=16'd11365;
      63026:data<=16'd11218;
      63027:data<=16'd15341;
      63028:data<=16'd16113;
      63029:data<=16'd12185;
      63030:data<=16'd12395;
      63031:data<=16'd18457;
      63032:data<=16'd18137;
      63033:data<=16'd13805;
      63034:data<=16'd12580;
      63035:data<=16'd10043;
      63036:data<=16'd13076;
      63037:data<=16'd16493;
      63038:data<=16'd8123;
      63039:data<=16'd6185;
      63040:data<=16'd12985;
      63041:data<=16'd11354;
      63042:data<=16'd8523;
      63043:data<=16'd8896;
      63044:data<=16'd6764;
      63045:data<=16'd4073;
      63046:data<=16'd3620;
      63047:data<=16'd5606;
      63048:data<=16'd3621;
      63049:data<=16'd1641;
      63050:data<=16'd6112;
      63051:data<=16'd1143;
      63052:data<=-16'd9730;
      63053:data<=-16'd7899;
      63054:data<=-16'd5847;
      63055:data<=-16'd12813;
      63056:data<=-16'd17377;
      63057:data<=-16'd14346;
      63058:data<=-16'd10648;
      63059:data<=-16'd13426;
      63060:data<=-16'd11916;
      63061:data<=-16'd4596;
      63062:data<=-16'd7512;
      63063:data<=-16'd12328;
      63064:data<=-16'd11224;
      63065:data<=-16'd13887;
      63066:data<=-16'd16342;
      63067:data<=-16'd14128;
      63068:data<=-16'd9373;
      63069:data<=-16'd8173;
      63070:data<=-16'd14016;
      63071:data<=-16'd12803;
      63072:data<=-16'd8599;
      63073:data<=-16'd13652;
      63074:data<=-16'd14067;
      63075:data<=-16'd12061;
      63076:data<=-16'd15144;
      63077:data<=-16'd12668;
      63078:data<=-16'd9142;
      63079:data<=-16'd8877;
      63080:data<=-16'd9611;
      63081:data<=-16'd10939;
      63082:data<=-16'd6984;
      63083:data<=-16'd6984;
      63084:data<=-16'd9069;
      63085:data<=16'd240;
      63086:data<=16'd1601;
      63087:data<=-16'd4752;
      63088:data<=16'd1606;
      63089:data<=16'd4366;
      63090:data<=-16'd743;
      63091:data<=16'd616;
      63092:data<=16'd1031;
      63093:data<=-16'd2021;
      63094:data<=-16'd1952;
      63095:data<=-16'd381;
      63096:data<=-16'd1527;
      63097:data<=-16'd3795;
      63098:data<=-16'd3054;
      63099:data<=-16'd4217;
      63100:data<=-16'd4661;
      63101:data<=-16'd1492;
      63102:data<=-16'd7306;
      63103:data<=-16'd12401;
      63104:data<=-16'd6763;
      63105:data<=-16'd6237;
      63106:data<=-16'd6384;
      63107:data<=-16'd2833;
      63108:data<=-16'd5406;
      63109:data<=-16'd7330;
      63110:data<=-16'd8790;
      63111:data<=-16'd9533;
      63112:data<=-16'd4390;
      63113:data<=-16'd5820;
      63114:data<=-16'd7709;
      63115:data<=-16'd1927;
      63116:data<=-16'd5234;
      63117:data<=-16'd12721;
      63118:data<=-16'd15165;
      63119:data<=-16'd18380;
      63120:data<=-16'd17253;
      63121:data<=-16'd16358;
      63122:data<=-16'd20721;
      63123:data<=-16'd17766;
      63124:data<=-16'd11232;
      63125:data<=-16'd12366;
      63126:data<=-16'd14187;
      63127:data<=-16'd11979;
      63128:data<=-16'd13609;
      63129:data<=-16'd15941;
      63130:data<=-16'd8511;
      63131:data<=-16'd5721;
      63132:data<=-16'd15682;
      63133:data<=-16'd17000;
      63134:data<=-16'd13640;
      63135:data<=-16'd17497;
      63136:data<=-16'd12874;
      63137:data<=-16'd6799;
      63138:data<=-16'd12800;
      63139:data<=-16'd14627;
      63140:data<=-16'd9025;
      63141:data<=-16'd6100;
      63142:data<=-16'd6951;
      63143:data<=-16'd10422;
      63144:data<=-16'd10103;
      63145:data<=-16'd7984;
      63146:data<=-16'd9591;
      63147:data<=-16'd5570;
      63148:data<=-16'd218;
      63149:data<=-16'd4246;
      63150:data<=-16'd4637;
      63151:data<=16'd2839;
      63152:data<=16'd7588;
      63153:data<=16'd11623;
      63154:data<=16'd13509;
      63155:data<=16'd9124;
      63156:data<=16'd7611;
      63157:data<=16'd10739;
      63158:data<=16'd12633;
      63159:data<=16'd13044;
      63160:data<=16'd10363;
      63161:data<=16'd9538;
      63162:data<=16'd12936;
      63163:data<=16'd8602;
      63164:data<=16'd3362;
      63165:data<=16'd9612;
      63166:data<=16'd12612;
      63167:data<=16'd9665;
      63168:data<=16'd11741;
      63169:data<=16'd11497;
      63170:data<=16'd10144;
      63171:data<=16'd14389;
      63172:data<=16'd13402;
      63173:data<=16'd7151;
      63174:data<=16'd6476;
      63175:data<=16'd8155;
      63176:data<=16'd6134;
      63177:data<=16'd3527;
      63178:data<=16'd5112;
      63179:data<=16'd8431;
      63180:data<=16'd9711;
      63181:data<=16'd11260;
      63182:data<=16'd12249;
      63183:data<=16'd10117;
      63184:data<=16'd6122;
      63185:data<=16'd1471;
      63186:data<=-16'd365;
      63187:data<=-16'd610;
      63188:data<=-16'd2287;
      63189:data<=-16'd15;
      63190:data<=16'd3562;
      63191:data<=16'd4871;
      63192:data<=16'd8637;
      63193:data<=16'd7433;
      63194:data<=16'd1077;
      63195:data<=-16'd82;
      63196:data<=-16'd1818;
      63197:data<=-16'd1022;
      63198:data<=16'd6945;
      63199:data<=16'd6238;
      63200:data<=16'd270;
      63201:data<=16'd2140;
      63202:data<=16'd6516;
      63203:data<=16'd10323;
      63204:data<=16'd10237;
      63205:data<=16'd6003;
      63206:data<=16'd3519;
      63207:data<=16'd1333;
      63208:data<=16'd5999;
      63209:data<=16'd13148;
      63210:data<=16'd7236;
      63211:data<=16'd4957;
      63212:data<=16'd9690;
      63213:data<=16'd4567;
      63214:data<=16'd5459;
      63215:data<=16'd9467;
      63216:data<=16'd1616;
      63217:data<=16'd6072;
      63218:data<=16'd19229;
      63219:data<=16'd17945;
      63220:data<=16'd16140;
      63221:data<=16'd16766;
      63222:data<=16'd12787;
      63223:data<=16'd14045;
      63224:data<=16'd15905;
      63225:data<=16'd12648;
      63226:data<=16'd12533;
      63227:data<=16'd14421;
      63228:data<=16'd14838;
      63229:data<=16'd14830;
      63230:data<=16'd11714;
      63231:data<=16'd9762;
      63232:data<=16'd16216;
      63233:data<=16'd19349;
      63234:data<=16'd11452;
      63235:data<=16'd9715;
      63236:data<=16'd13341;
      63237:data<=16'd8229;
      63238:data<=16'd6628;
      63239:data<=16'd9649;
      63240:data<=16'd5968;
      63241:data<=16'd6757;
      63242:data<=16'd11218;
      63243:data<=16'd9723;
      63244:data<=16'd7791;
      63245:data<=16'd4924;
      63246:data<=16'd5010;
      63247:data<=16'd8440;
      63248:data<=16'd2781;
      63249:data<=-16'd670;
      63250:data<=16'd3923;
      63251:data<=-16'd1627;
      63252:data<=-16'd11226;
      63253:data<=-16'd12038;
      63254:data<=-16'd10522;
      63255:data<=-16'd10981;
      63256:data<=-16'd11065;
      63257:data<=-16'd7050;
      63258:data<=-16'd6290;
      63259:data<=-16'd13534;
      63260:data<=-16'd12507;
      63261:data<=-16'd7247;
      63262:data<=-16'd13718;
      63263:data<=-16'd16123;
      63264:data<=-16'd9201;
      63265:data<=-16'd9573;
      63266:data<=-16'd11819;
      63267:data<=-16'd9016;
      63268:data<=-16'd10357;
      63269:data<=-16'd12047;
      63270:data<=-16'd6357;
      63271:data<=-16'd4311;
      63272:data<=-16'd9144;
      63273:data<=-16'd7953;
      63274:data<=-16'd5391;
      63275:data<=-16'd9831;
      63276:data<=-16'd11899;
      63277:data<=-16'd10610;
      63278:data<=-16'd10847;
      63279:data<=-16'd12231;
      63280:data<=-16'd14128;
      63281:data<=-16'd8510;
      63282:data<=-16'd3586;
      63283:data<=-16'd11994;
      63284:data<=-16'd11091;
      63285:data<=16'd1498;
      63286:data<=16'd1618;
      63287:data<=16'd1462;
      63288:data<=16'd5802;
      63289:data<=-16'd946;
      63290:data<=-16'd6291;
      63291:data<=-16'd6141;
      63292:data<=-16'd7859;
      63293:data<=-16'd1686;
      63294:data<=16'd3062;
      63295:data<=-16'd4684;
      63296:data<=-16'd7941;
      63297:data<=-16'd4593;
      63298:data<=-16'd5265;
      63299:data<=-16'd4992;
      63300:data<=-16'd3730;
      63301:data<=-16'd5779;
      63302:data<=-16'd4425;
      63303:data<=-16'd852;
      63304:data<=-16'd3968;
      63305:data<=-16'd7582;
      63306:data<=-16'd5523;
      63307:data<=-16'd6213;
      63308:data<=-16'd8795;
      63309:data<=-16'd5979;
      63310:data<=-16'd4652;
      63311:data<=-16'd8251;
      63312:data<=-16'd9630;
      63313:data<=-16'd8184;
      63314:data<=-16'd6570;
      63315:data<=-16'd6972;
      63316:data<=-16'd11198;
      63317:data<=-16'd13700;
      63318:data<=-16'd12941;
      63319:data<=-16'd14657;
      63320:data<=-16'd15177;
      63321:data<=-16'd14205;
      63322:data<=-16'd20524;
      63323:data<=-16'd24095;
      63324:data<=-16'd15279;
      63325:data<=-16'd11797;
      63326:data<=-16'd16930;
      63327:data<=-16'd13388;
      63328:data<=-16'd7817;
      63329:data<=-16'd11866;
      63330:data<=-16'd15107;
      63331:data<=-16'd12516;
      63332:data<=-16'd10745;
      63333:data<=-16'd9843;
      63334:data<=-16'd9135;
      63335:data<=-16'd11203;
      63336:data<=-16'd10140;
      63337:data<=-16'd4128;
      63338:data<=-16'd6169;
      63339:data<=-16'd11496;
      63340:data<=-16'd5762;
      63341:data<=-16'd3354;
      63342:data<=-16'd9063;
      63343:data<=-16'd6763;
      63344:data<=-16'd3375;
      63345:data<=-16'd3459;
      63346:data<=-16'd494;
      63347:data<=-16'd1495;
      63348:data<=-16'd1507;
      63349:data<=16'd2531;
      63350:data<=16'd1445;
      63351:data<=16'd5835;
      63352:data<=16'd13283;
      63353:data<=16'd9589;
      63354:data<=16'd7847;
      63355:data<=16'd9429;
      63356:data<=16'd5808;
      63357:data<=16'd6786;
      63358:data<=16'd11003;
      63359:data<=16'd13987;
      63360:data<=16'd15245;
      63361:data<=16'd8385;
      63362:data<=16'd5269;
      63363:data<=16'd11621;
      63364:data<=16'd13345;
      63365:data<=16'd14757;
      63366:data<=16'd16119;
      63367:data<=16'd8272;
      63368:data<=16'd5491;
      63369:data<=16'd10423;
      63370:data<=16'd7994;
      63371:data<=16'd5142;
      63372:data<=16'd8686;
      63373:data<=16'd10278;
      63374:data<=16'd9838;
      63375:data<=16'd10652;
      63376:data<=16'd12002;
      63377:data<=16'd13412;
      63378:data<=16'd13436;
      63379:data<=16'd13659;
      63380:data<=16'd13493;
      63381:data<=16'd10595;
      63382:data<=16'd11082;
      63383:data<=16'd11544;
      63384:data<=16'd3964;
      63385:data<=16'd610;
      63386:data<=16'd2896;
      63387:data<=-16'd984;
      63388:data<=-16'd1036;
      63389:data<=16'd4244;
      63390:data<=16'd2908;
      63391:data<=16'd2638;
      63392:data<=16'd5046;
      63393:data<=16'd2669;
      63394:data<=16'd2573;
      63395:data<=16'd6743;
      63396:data<=16'd8122;
      63397:data<=16'd5873;
      63398:data<=16'd5564;
      63399:data<=16'd7785;
      63400:data<=16'd3601;
      63401:data<=-16'd711;
      63402:data<=16'd4447;
      63403:data<=16'd6539;
      63404:data<=16'd6024;
      63405:data<=16'd9711;
      63406:data<=16'd6499;
      63407:data<=16'd2237;
      63408:data<=16'd5632;
      63409:data<=16'd6404;
      63410:data<=16'd4813;
      63411:data<=16'd5350;
      63412:data<=16'd6630;
      63413:data<=16'd8699;
      63414:data<=16'd9185;
      63415:data<=16'd8120;
      63416:data<=16'd5735;
      63417:data<=16'd8090;
      63418:data<=16'd19992;
      63419:data<=16'd22703;
      63420:data<=16'd14803;
      63421:data<=16'd16001;
      63422:data<=16'd16797;
      63423:data<=16'd13496;
      63424:data<=16'd16697;
      63425:data<=16'd14724;
      63426:data<=16'd12163;
      63427:data<=16'd20621;
      63428:data<=16'd20967;
      63429:data<=16'd12389;
      63430:data<=16'd12771;
      63431:data<=16'd15703;
      63432:data<=16'd15979;
      63433:data<=16'd16880;
      63434:data<=16'd12342;
      63435:data<=16'd7407;
      63436:data<=16'd9168;
      63437:data<=16'd8915;
      63438:data<=16'd10220;
      63439:data<=16'd16126;
      63440:data<=16'd12502;
      63441:data<=16'd7491;
      63442:data<=16'd10884;
      63443:data<=16'd8983;
      63444:data<=16'd6184;
      63445:data<=16'd7887;
      63446:data<=16'd4390;
      63447:data<=16'd1287;
      63448:data<=16'd1237;
      63449:data<=16'd2270;
      63450:data<=16'd3450;
      63451:data<=-16'd5645;
      63452:data<=-16'd13056;
      63453:data<=-16'd8937;
      63454:data<=-16'd9194;
      63455:data<=-16'd8294;
      63456:data<=-16'd5433;
      63457:data<=-16'd11373;
      63458:data<=-16'd10909;
      63459:data<=-16'd5976;
      63460:data<=-16'd8630;
      63461:data<=-16'd10073;
      63462:data<=-16'd9749;
      63463:data<=-16'd6398;
      63464:data<=-16'd4952;
      63465:data<=-16'd13386;
      63466:data<=-16'd12499;
      63467:data<=-16'd5544;
      63468:data<=-16'd8875;
      63469:data<=-16'd6960;
      63470:data<=-16'd4261;
      63471:data<=-16'd11380;
      63472:data<=-16'd12102;
      63473:data<=-16'd7749;
      63474:data<=-16'd7812;
      63475:data<=-16'd10082;
      63476:data<=-16'd11624;
      63477:data<=-16'd10141;
      63478:data<=-16'd12192;
      63479:data<=-16'd15026;
      63480:data<=-16'd10185;
      63481:data<=-16'd8734;
      63482:data<=-16'd12342;
      63483:data<=-16'd11741;
      63484:data<=-16'd7144;
      63485:data<=16'd332;
      63486:data<=16'd3442;
      63487:data<=16'd2470;
      63488:data<=16'd3550;
      63489:data<=-16'd632;
      63490:data<=-16'd2362;
      63491:data<=16'd2714;
      63492:data<=-16'd2043;
      63493:data<=-16'd4303;
      63494:data<=16'd4664;
      63495:data<=16'd1579;
      63496:data<=-16'd8621;
      63497:data<=-16'd10713;
      63498:data<=-16'd12064;
      63499:data<=-16'd9879;
      63500:data<=-16'd3756;
      63501:data<=-16'd4379;
      63502:data<=-16'd5542;
      63503:data<=-16'd3166;
      63504:data<=-16'd5577;
      63505:data<=-16'd8830;
      63506:data<=-16'd9235;
      63507:data<=-16'd13423;
      63508:data<=-16'd16747;
      63509:data<=-16'd10376;
      63510:data<=-16'd1557;
      63511:data<=-16'd2602;
      63512:data<=-16'd10163;
      63513:data<=-16'd11094;
      63514:data<=-16'd7573;
      63515:data<=-16'd8134;
      63516:data<=-16'd8940;
      63517:data<=-16'd12060;
      63518:data<=-16'd18556;
      63519:data<=-16'd18330;
      63520:data<=-16'd17561;
      63521:data<=-16'd20397;
      63522:data<=-16'd16888;
      63523:data<=-16'd15242;
      63524:data<=-16'd17673;
      63525:data<=-16'd14260;
      63526:data<=-16'd17540;
      63527:data<=-16'd26753;
      63528:data<=-16'd21510;
      63529:data<=-16'd12977;
      63530:data<=-16'd15559;
      63531:data<=-16'd14956;
      63532:data<=-16'd10205;
      63533:data<=-16'd13035;
      63534:data<=-16'd14029;
      63535:data<=-16'd9132;
      63536:data<=-16'd8507;
      63537:data<=-16'd7024;
      63538:data<=-16'd5635;
      63539:data<=-16'd12759;
      63540:data<=-16'd15015;
      63541:data<=-16'd10458;
      63542:data<=-16'd11235;
      63543:data<=-16'd10889;
      63544:data<=-16'd8968;
      63545:data<=-16'd11089;
      63546:data<=-16'd10765;
      63547:data<=-16'd6357;
      63548:data<=-16'd2231;
      63549:data<=-16'd4027;
      63550:data<=-16'd5512;
      63551:data<=16'd6319;
      63552:data<=16'd15938;
      63553:data<=16'd12228;
      63554:data<=16'd10810;
      63555:data<=16'd12557;
      63556:data<=16'd14615;
      63557:data<=16'd17282;
      63558:data<=16'd13759;
      63559:data<=16'd13232;
      63560:data<=16'd17579;
      63561:data<=16'd13596;
      63562:data<=16'd8432;
      63563:data<=16'd9057;
      63564:data<=16'd9929;
      63565:data<=16'd11051;
      63566:data<=16'd11536;
      63567:data<=16'd11100;
      63568:data<=16'd11435;
      63569:data<=16'd10240;
      63570:data<=16'd9749;
      63571:data<=16'd13882;
      63572:data<=16'd15336;
      63573:data<=16'd11033;
      63574:data<=16'd13073;
      63575:data<=16'd15068;
      63576:data<=16'd6693;
      63577:data<=16'd9016;
      63578:data<=16'd17807;
      63579:data<=16'd12666;
      63580:data<=16'd12020;
      63581:data<=16'd13584;
      63582:data<=16'd7874;
      63583:data<=16'd13811;
      63584:data<=16'd14897;
      63585:data<=16'd3360;
      63586:data<=16'd1624;
      63587:data<=16'd45;
      63588:data<=16'd867;
      63589:data<=16'd7354;
      63590:data<=16'd860;
      63591:data<=-16'd1061;
      63592:data<=16'd6282;
      63593:data<=16'd3266;
      63594:data<=-16'd579;
      63595:data<=-16'd863;
      63596:data<=16'd3983;
      63597:data<=16'd10257;
      63598:data<=16'd4024;
      63599:data<=16'd3692;
      63600:data<=16'd9586;
      63601:data<=16'd5554;
      63602:data<=16'd7721;
      63603:data<=16'd7984;
      63604:data<=16'd2126;
      63605:data<=16'd7944;
      63606:data<=16'd7204;
      63607:data<=16'd2206;
      63608:data<=16'd9620;
      63609:data<=16'd10208;
      63610:data<=16'd4572;
      63611:data<=16'd2648;
      63612:data<=16'd1574;
      63613:data<=16'd4507;
      63614:data<=16'd6654;
      63615:data<=16'd10734;
      63616:data<=16'd14963;
      63617:data<=16'd10222;
      63618:data<=16'd11958;
      63619:data<=16'd16152;
      63620:data<=16'd11148;
      63621:data<=16'd13878;
      63622:data<=16'd20134;
      63623:data<=16'd20671;
      63624:data<=16'd19382;
      63625:data<=16'd13941;
      63626:data<=16'd15571;
      63627:data<=16'd20948;
      63628:data<=16'd17515;
      63629:data<=16'd17478;
      63630:data<=16'd16399;
      63631:data<=16'd10288;
      63632:data<=16'd12590;
      63633:data<=16'd14455;
      63634:data<=16'd12968;
      63635:data<=16'd15361;
      63636:data<=16'd15133;
      63637:data<=16'd13092;
      63638:data<=16'd9746;
      63639:data<=16'd3885;
      63640:data<=16'd2475;
      63641:data<=16'd4969;
      63642:data<=16'd7121;
      63643:data<=16'd7868;
      63644:data<=16'd9705;
      63645:data<=16'd10887;
      63646:data<=16'd5946;
      63647:data<=16'd4916;
      63648:data<=16'd5116;
      63649:data<=-16'd3274;
      63650:data<=-16'd591;
      63651:data<=16'd6062;
      63652:data<=-16'd6388;
      63653:data<=-16'd15898;
      63654:data<=-16'd13298;
      63655:data<=-16'd13170;
      63656:data<=-16'd12992;
      63657:data<=-16'd13523;
      63658:data<=-16'd14681;
      63659:data<=-16'd14818;
      63660:data<=-16'd16186;
      63661:data<=-16'd10962;
      63662:data<=-16'd5004;
      63663:data<=-16'd8108;
      63664:data<=-16'd10649;
      63665:data<=-16'd11166;
      63666:data<=-16'd12232;
      63667:data<=-16'd11891;
      63668:data<=-16'd13403;
      63669:data<=-16'd13291;
      63670:data<=-16'd9310;
      63671:data<=-16'd6913;
      63672:data<=-16'd7962;
      63673:data<=-16'd10172;
      63674:data<=-16'd9018;
      63675:data<=-16'd8715;
      63676:data<=-16'd12621;
      63677:data<=-16'd12096;
      63678:data<=-16'd9708;
      63679:data<=-16'd10220;
      63680:data<=-16'd9488;
      63681:data<=-16'd10470;
      63682:data<=-16'd12116;
      63683:data<=-16'd11620;
      63684:data<=-16'd10085;
      63685:data<=-16'd4490;
      63686:data<=-16'd1715;
      63687:data<=-16'd2452;
      63688:data<=16'd2874;
      63689:data<=16'd3545;
      63690:data<=-16'd2491;
      63691:data<=-16'd1924;
      63692:data<=-16'd2723;
      63693:data<=-16'd8510;
      63694:data<=-16'd6845;
      63695:data<=-16'd814;
      63696:data<=-16'd1521;
      63697:data<=-16'd5190;
      63698:data<=-16'd3245;
      63699:data<=-16'd3227;
      63700:data<=-16'd8204;
      63701:data<=-16'd5262;
      63702:data<=-16'd2502;
      63703:data<=-16'd9477;
      63704:data<=-16'd10672;
      63705:data<=-16'd6862;
      63706:data<=-16'd6258;
      63707:data<=-16'd5084;
      63708:data<=-16'd9771;
      63709:data<=-16'd14492;
      63710:data<=-16'd7649;
      63711:data<=-16'd3444;
      63712:data<=-16'd5700;
      63713:data<=-16'd5567;
      63714:data<=-16'd7914;
      63715:data<=-16'd9815;
      63716:data<=-16'd6690;
      63717:data<=-16'd7183;
      63718:data<=-16'd12172;
      63719:data<=-16'd15528;
      63720:data<=-16'd16785;
      63721:data<=-16'd17206;
      63722:data<=-16'd14906;
      63723:data<=-16'd12116;
      63724:data<=-16'd17511;
      63725:data<=-16'd21822;
      63726:data<=-16'd13562;
      63727:data<=-16'd12985;
      63728:data<=-16'd22054;
      63729:data<=-16'd18530;
      63730:data<=-16'd17285;
      63731:data<=-16'd24658;
      63732:data<=-16'd17299;
      63733:data<=-16'd8698;
      63734:data<=-16'd13174;
      63735:data<=-16'd14942;
      63736:data<=-16'd14041;
      63737:data<=-16'd10328;
      63738:data<=-16'd4273;
      63739:data<=-16'd9790;
      63740:data<=-16'd13787;
      63741:data<=-16'd7680;
      63742:data<=-16'd7735;
      63743:data<=-16'd7266;
      63744:data<=-16'd3180;
      63745:data<=-16'd4676;
      63746:data<=-16'd3439;
      63747:data<=-16'd1874;
      63748:data<=-16'd2190;
      63749:data<=16'd610;
      63750:data<=-16'd4965;
      63751:data<=-16'd6764;
      63752:data<=16'd9197;
      63753:data<=16'd17177;
      63754:data<=16'd12975;
      63755:data<=16'd11696;
      63756:data<=16'd11583;
      63757:data<=16'd15123;
      63758:data<=16'd15632;
      63759:data<=16'd8760;
      63760:data<=16'd8643;
      63761:data<=16'd12536;
      63762:data<=16'd15746;
      63763:data<=16'd17749;
      63764:data<=16'd10883;
      63765:data<=16'd8522;
      63766:data<=16'd14765;
      63767:data<=16'd14181;
      63768:data<=16'd13003;
      63769:data<=16'd13535;
      63770:data<=16'd12123;
      63771:data<=16'd12578;
      63772:data<=16'd8247;
      63773:data<=16'd7620;
      63774:data<=16'd14832;
      63775:data<=16'd13295;
      63776:data<=16'd12837;
      63777:data<=16'd14953;
      63778:data<=16'd10328;
      63779:data<=16'd16568;
      63780:data<=16'd19303;
      63781:data<=16'd5172;
      63782:data<=16'd6789;
      63783:data<=16'd17147;
      63784:data<=16'd14164;
      63785:data<=16'd9447;
      63786:data<=16'd1730;
      63787:data<=-16'd1874;
      63788:data<=16'd7291;
      63789:data<=16'd7741;
      63790:data<=16'd2720;
      63791:data<=16'd7912;
      63792:data<=16'd12419;
      63793:data<=16'd13688;
      63794:data<=16'd14431;
      63795:data<=16'd11147;
      63796:data<=16'd9803;
      63797:data<=16'd12216;
      63798:data<=16'd13591;
      63799:data<=16'd13691;
      63800:data<=16'd12554;
      63801:data<=16'd11394;
      63802:data<=16'd12213;
      63803:data<=16'd13180;
      63804:data<=16'd12434;
      63805:data<=16'd12169;
      63806:data<=16'd12933;
      63807:data<=16'd11844;
      63808:data<=16'd11220;
      63809:data<=16'd12674;
      63810:data<=16'd11869;
      63811:data<=16'd10692;
      63812:data<=16'd12305;
      63813:data<=16'd12689;
      63814:data<=16'd11039;
      63815:data<=16'd11394;
      63816:data<=16'd13118;
      63817:data<=16'd11629;
      63818:data<=16'd11238;
      63819:data<=16'd17631;
      63820:data<=16'd21303;
      63821:data<=16'd19188;
      63822:data<=16'd19999;
      63823:data<=16'd20735;
      63824:data<=16'd19754;
      63825:data<=16'd19822;
      63826:data<=16'd16807;
      63827:data<=16'd15720;
      63828:data<=16'd19171;
      63829:data<=16'd17845;
      63830:data<=16'd14427;
      63831:data<=16'd14622;
      63832:data<=16'd14892;
      63833:data<=16'd14416;
      63834:data<=16'd13741;
      63835:data<=16'd13581;
      63836:data<=16'd14216;
      63837:data<=16'd13154;
      63838:data<=16'd12061;
      63839:data<=16'd12240;
      63840:data<=16'd10483;
      63841:data<=16'd8548;
      63842:data<=16'd9508;
      63843:data<=16'd9138;
      63844:data<=16'd6134;
      63845:data<=16'd6090;
      63846:data<=16'd6625;
      63847:data<=16'd3403;
      63848:data<=16'd1695;
      63849:data<=16'd1457;
      63850:data<=16'd790;
      63851:data<=16'd1936;
      63852:data<=-16'd2823;
      63853:data<=-16'd12098;
      63854:data<=-16'd12413;
      63855:data<=-16'd9685;
      63856:data<=-16'd11623;
      63857:data<=-16'd11840;
      63858:data<=-16'd11022;
      63859:data<=-16'd12219;
      63860:data<=-16'd13063;
      63861:data<=-16'd13042;
      63862:data<=-16'd12812;
      63863:data<=-16'd12645;
      63864:data<=-16'd12114;
      63865:data<=-16'd13144;
      63866:data<=-16'd15901;
      63867:data<=-16'd15032;
      63868:data<=-16'd12666;
      63869:data<=-16'd13024;
      63870:data<=-16'd12933;
      63871:data<=-16'd13388;
      63872:data<=-16'd14903;
      63873:data<=-16'd14148;
      63874:data<=-16'd13409;
      63875:data<=-16'd14199;
      63876:data<=-16'd14690;
      63877:data<=-16'd14255;
      63878:data<=-16'd13529;
      63879:data<=-16'd13976;
      63880:data<=-16'd13841;
      63881:data<=-16'd12643;
      63882:data<=-16'd13060;
      63883:data<=-16'd14226;
      63884:data<=-16'd15033;
      63885:data<=-16'd12160;
      63886:data<=-16'd4108;
      63887:data<=-16'd406;
      63888:data<=-16'd2772;
      63889:data<=-16'd3162;
      63890:data<=-16'd3497;
      63891:data<=-16'd5824;
      63892:data<=-16'd6628;
      63893:data<=-16'd6463;
      63894:data<=-16'd5944;
      63895:data<=-16'd5153;
      63896:data<=-16'd5762;
      63897:data<=-16'd6918;
      63898:data<=-16'd7168;
      63899:data<=-16'd7489;
      63900:data<=-16'd7686;
      63901:data<=-16'd6244;
      63902:data<=-16'd5974;
      63903:data<=-16'd8583;
      63904:data<=-16'd9602;
      63905:data<=-16'd8786;
      63906:data<=-16'd8273;
      63907:data<=-16'd6949;
      63908:data<=-16'd7406;
      63909:data<=-16'd10060;
      63910:data<=-16'd10605;
      63911:data<=-16'd9374;
      63912:data<=-16'd8405;
      63913:data<=-16'd7915;
      63914:data<=-16'd7351;
      63915:data<=-16'd8073;
      63916:data<=-16'd11480;
      63917:data<=-16'd11106;
      63918:data<=-16'd7844;
      63919:data<=-16'd12700;
      63920:data<=-16'd19811;
      63921:data<=-16'd20260;
      63922:data<=-16'd20108;
      63923:data<=-16'd19863;
      63924:data<=-16'd17791;
      63925:data<=-16'd18368;
      63926:data<=-16'd19071;
      63927:data<=-16'd16909;
      63928:data<=-16'd16355;
      63929:data<=-16'd18322;
      63930:data<=-16'd18231;
      63931:data<=-16'd15876;
      63932:data<=-16'd14609;
      63933:data<=-16'd13832;
      63934:data<=-16'd13917;
      63935:data<=-16'd15887;
      63936:data<=-16'd15684;
      63937:data<=-16'd13976;
      63938:data<=-16'd14255;
      63939:data<=-16'd13920;
      63940:data<=-16'd12213;
      63941:data<=-16'd10586;
      63942:data<=-16'd9644;
      63943:data<=-16'd9624;
      63944:data<=-16'd8739;
      63945:data<=-16'd8287;
      63946:data<=-16'd7978;
      63947:data<=-16'd5454;
      63948:data<=-16'd4821;
      63949:data<=-16'd4827;
      63950:data<=-16'd3312;
      63951:data<=-16'd5004;
      63952:data<=-16'd2487;
      63953:data<=16'd7377;
      63954:data<=16'd10877;
      63955:data<=16'd9047;
      63956:data<=16'd10158;
      63957:data<=16'd10166;
      63958:data<=16'd9256;
      63959:data<=16'd10393;
      63960:data<=16'd10332;
      63961:data<=16'd9585;
      63962:data<=16'd10971;
      63963:data<=16'd11453;
      63964:data<=16'd10243;
      63965:data<=16'd11485;
      63966:data<=16'd12137;
      63967:data<=16'd10160;
      63968:data<=16'd11174;
      63969:data<=16'd11759;
      63970:data<=16'd9647;
      63971:data<=16'd11065;
      63972:data<=16'd12249;
      63973:data<=16'd11630;
      63974:data<=16'd13071;
      63975:data<=16'd12143;
      63976:data<=16'd10960;
      63977:data<=16'd12410;
      63978:data<=16'd11580;
      63979:data<=16'd11165;
      63980:data<=16'd12169;
      63981:data<=16'd11963;
      63982:data<=16'd11905;
      63983:data<=16'd10331;
      63984:data<=16'd10712;
      63985:data<=16'd13480;
      63986:data<=16'd8868;
      63987:data<=16'd1609;
      63988:data<=16'd328;
      63989:data<=16'd694;
      63990:data<=16'd1559;
      63991:data<=16'd3519;
      63992:data<=16'd4431;
      63993:data<=16'd4070;
      63994:data<=16'd2883;
      63995:data<=16'd2679;
      63996:data<=16'd2796;
      63997:data<=16'd3112;
      63998:data<=16'd5272;
      63999:data<=16'd5409;
      64000:data<=16'd3871;
      64001:data<=16'd4167;
      64002:data<=16'd4440;
      64003:data<=16'd5295;
      64004:data<=16'd5618;
      64005:data<=16'd4625;
      64006:data<=16'd5448;
      64007:data<=16'd4573;
      64008:data<=16'd3189;
      64009:data<=16'd5100;
      64010:data<=16'd4901;
      64011:data<=16'd4626;
      64012:data<=16'd6261;
      64013:data<=16'd5090;
      64014:data<=16'd4681;
      64015:data<=16'd5274;
      64016:data<=16'd5130;
      64017:data<=16'd6391;
      64018:data<=16'd5444;
      64019:data<=16'd6946;
      64020:data<=16'd14084;
      64021:data<=16'd16126;
      64022:data<=16'd15579;
      64023:data<=16'd17660;
      64024:data<=16'd16543;
      64025:data<=16'd15012;
      64026:data<=16'd14507;
      64027:data<=16'd12424;
      64028:data<=16'd13391;
      64029:data<=16'd15632;
      64030:data<=16'd14894;
      64031:data<=16'd14542;
      64032:data<=16'd14795;
      64033:data<=16'd13379;
      64034:data<=16'd12175;
      64035:data<=16'd12954;
      64036:data<=16'd13479;
      64037:data<=16'd12472;
      64038:data<=16'd12208;
      64039:data<=16'd11981;
      64040:data<=16'd10636;
      64041:data<=16'd10181;
      64042:data<=16'd10160;
      64043:data<=16'd9538;
      64044:data<=16'd8436;
      64045:data<=16'd7272;
      64046:data<=16'd6905;
      64047:data<=16'd5529;
      64048:data<=16'd4156;
      64049:data<=16'd4934;
      64050:data<=16'd4170;
      64051:data<=16'd2927;
      64052:data<=16'd2443;
      64053:data<=-16'd3334;
      64054:data<=-16'd10439;
      64055:data<=-16'd11380;
      64056:data<=-16'd10921;
      64057:data<=-16'd11497;
      64058:data<=-16'd10147;
      64059:data<=-16'd9832;
      64060:data<=-16'd11896;
      64061:data<=-16'd11838;
      64062:data<=-16'd10695;
      64063:data<=-16'd11911;
      64064:data<=-16'd12330;
      64065:data<=-16'd11981;
      64066:data<=-16'd13641;
      64067:data<=-16'd14008;
      64068:data<=-16'd13405;
      64069:data<=-16'd14029;
      64070:data<=-16'd13244;
      64071:data<=-16'd12436;
      64072:data<=-16'd13233;
      64073:data<=-16'd14220;
      64074:data<=-16'd15100;
      64075:data<=-16'd14160;
      64076:data<=-16'd13100;
      64077:data<=-16'd13535;
      64078:data<=-16'd13113;
      64079:data<=-16'd14032;
      64080:data<=-16'd14847;
      64081:data<=-16'd13107;
      64082:data<=-16'd13665;
      64083:data<=-16'd13653;
      64084:data<=-16'd11978;
      64085:data<=-16'd14181;
      64086:data<=-16'd12481;
      64087:data<=-16'd4366;
      64088:data<=-16'd980;
      64089:data<=-16'd1929;
      64090:data<=-16'd2153;
      64091:data<=-16'd3143;
      64092:data<=-16'd5121;
      64093:data<=-16'd6220;
      64094:data<=-16'd5119;
      64095:data<=-16'd3557;
      64096:data<=-16'd3422;
      64097:data<=-16'd4179;
      64098:data<=-16'd5275;
      64099:data<=-16'd4934;
      64100:data<=-16'd4498;
      64101:data<=-16'd5785;
      64102:data<=-16'd5415;
      64103:data<=-16'd4963;
      64104:data<=-16'd6276;
      64105:data<=-16'd6067;
      64106:data<=-16'd6441;
      64107:data<=-16'd7233;
      64108:data<=-16'd5715;
      64109:data<=-16'd5626;
      64110:data<=-16'd6755;
      64111:data<=-16'd6751;
      64112:data<=-16'd6675;
      64113:data<=-16'd6008;
      64114:data<=-16'd6031;
      64115:data<=-16'd6698;
      64116:data<=-16'd6701;
      64117:data<=-16'd7736;
      64118:data<=-16'd7776;
      64119:data<=-16'd8034;
      64120:data<=-16'd13230;
      64121:data<=-16'd18331;
      64122:data<=-16'd19382;
      64123:data<=-16'd19132;
      64124:data<=-16'd18607;
      64125:data<=-16'd18571;
      64126:data<=-16'd17493;
      64127:data<=-16'd15546;
      64128:data<=-16'd16506;
      64129:data<=-16'd17020;
      64130:data<=-16'd15288;
      64131:data<=-16'd15749;
      64132:data<=-16'd15964;
      64133:data<=-16'd13993;
      64134:data<=-16'd13581;
      64135:data<=-16'd13758;
      64136:data<=-16'd13297;
      64137:data<=-16'd13834;
      64138:data<=-16'd13514;
      64139:data<=-16'd11935;
      64140:data<=-16'd11785;
      64141:data<=-16'd11568;
      64142:data<=-16'd10322;
      64143:data<=-16'd10316;
      64144:data<=-16'd9670;
      64145:data<=-16'd8448;
      64146:data<=-16'd9224;
      64147:data<=-16'd7169;
      64148:data<=-16'd3488;
      64149:data<=-16'd4783;
      64150:data<=-16'd4407;
      64151:data<=-16'd1811;
      64152:data<=-16'd3946;
      64153:data<=16'd64;
      64154:data<=16'd11420;
      64155:data<=16'd13420;
      64156:data<=16'd10566;
      64157:data<=16'd12243;
      64158:data<=16'd12040;
      64159:data<=16'd11638;
      64160:data<=16'd13884;
      64161:data<=16'd13493;
      64162:data<=16'd13059;
      64163:data<=16'd14396;
      64164:data<=16'd13790;
      64165:data<=16'd13242;
      64166:data<=16'd13934;
      64167:data<=16'd14075;
      64168:data<=16'd13987;
      64169:data<=16'd13797;
      64170:data<=16'd13958;
      64171:data<=16'd13602;
      64172:data<=16'd12577;
      64173:data<=16'd13809;
      64174:data<=16'd14698;
      64175:data<=16'd13063;
      64176:data<=16'd13279;
      64177:data<=16'd13781;
      64178:data<=16'd12719;
      64179:data<=16'd14257;
      64180:data<=16'd15520;
      64181:data<=16'd13591;
      64182:data<=16'd13256;
      64183:data<=16'd13878;
      64184:data<=16'd13082;
      64185:data<=16'd14125;
      64186:data<=16'd14252;
      64187:data<=16'd8308;
      64188:data<=16'd2335;
      64189:data<=16'd1730;
      64190:data<=16'd2074;
      64191:data<=16'd2602;
      64192:data<=16'd4720;
      64193:data<=16'd4628;
      64194:data<=16'd3636;
      64195:data<=16'd4293;
      64196:data<=16'd3438;
      64197:data<=16'd3262;
      64198:data<=16'd5494;
      64199:data<=16'd5410;
      64200:data<=16'd4589;
      64201:data<=16'd5301;
      64202:data<=16'd5048;
      64203:data<=16'd5577;
      64204:data<=16'd6883;
      64205:data<=16'd6686;
      64206:data<=16'd6825;
      64207:data<=16'd6024;
      64208:data<=16'd4212;
      64209:data<=16'd5830;
      64210:data<=16'd8446;
      64211:data<=16'd8668;
      64212:data<=16'd8002;
      64213:data<=16'd7116;
      64214:data<=16'd7952;
      64215:data<=16'd9066;
      64216:data<=16'd8120;
      64217:data<=16'd9676;
      64218:data<=16'd10261;
      64219:data<=16'd6845;
      64220:data<=16'd10666;
      64221:data<=16'd18304;
      64222:data<=16'd18780;
      64223:data<=16'd19438;
      64224:data<=16'd20682;
      64225:data<=16'd17640;
      64226:data<=16'd17438;
      64227:data<=16'd17920;
      64228:data<=16'd15860;
      64229:data<=16'd17887;
      64230:data<=16'd19713;
      64231:data<=16'd17863;
      64232:data<=16'd18017;
      64233:data<=16'd17508;
      64234:data<=16'd15167;
      64235:data<=16'd15728;
      64236:data<=16'd16472;
      64237:data<=16'd15161;
      64238:data<=16'd14665;
      64239:data<=16'd14170;
      64240:data<=16'd12710;
      64241:data<=16'd12425;
      64242:data<=16'd12393;
      64243:data<=16'd11035;
      64244:data<=16'd10060;
      64245:data<=16'd9712;
      64246:data<=16'd9354;
      64247:data<=16'd8449;
      64248:data<=16'd5947;
      64249:data<=16'd4726;
      64250:data<=16'd4792;
      64251:data<=16'd3242;
      64252:data<=16'd3704;
      64253:data<=16'd2616;
      64254:data<=-16'd6029;
      64255:data<=-16'd11952;
      64256:data<=-16'd11212;
      64257:data<=-16'd11339;
      64258:data<=-16'd10872;
      64259:data<=-16'd9897;
      64260:data<=-16'd11568;
      64261:data<=-16'd12527;
      64262:data<=-16'd12187;
      64263:data<=-16'd12205;
      64264:data<=-16'd12123;
      64265:data<=-16'd12272;
      64266:data<=-16'd12792;
      64267:data<=-16'd13436;
      64268:data<=-16'd13168;
      64269:data<=-16'd12580;
      64270:data<=-16'd12941;
      64271:data<=-16'd12298;
      64272:data<=-16'd11711;
      64273:data<=-16'd12766;
      64274:data<=-16'd13320;
      64275:data<=-16'd13655;
      64276:data<=-16'd13235;
      64277:data<=-16'd11876;
      64278:data<=-16'd12003;
      64279:data<=-16'd12787;
      64280:data<=-16'd13960;
      64281:data<=-16'd13819;
      64282:data<=-16'd11586;
      64283:data<=-16'd12301;
      64284:data<=-16'd12554;
      64285:data<=-16'd11057;
      64286:data<=-16'd13649;
      64287:data<=-16'd10977;
      64288:data<=-16'd1792;
      64289:data<=16'd71;
      64290:data<=-16'd1381;
      64291:data<=-16'd1228;
      64292:data<=-16'd3092;
      64293:data<=-16'd2999;
      64294:data<=-16'd2496;
      64295:data<=-16'd3841;
      64296:data<=-16'd2858;
      64297:data<=-16'd2604;
      64298:data<=-16'd4399;
      64299:data<=-16'd4764;
      64300:data<=-16'd4526;
      64301:data<=-16'd4012;
      64302:data<=-16'd3425;
      64303:data<=-16'd3694;
      64304:data<=-16'd4589;
      64305:data<=-16'd6028;
      64306:data<=-16'd6393;
      64307:data<=-16'd5583;
      64308:data<=-16'd5194;
      64309:data<=-16'd5084;
      64310:data<=-16'd5515;
      64311:data<=-16'd6167;
      64312:data<=-16'd6693;
      64313:data<=-16'd7228;
      64314:data<=-16'd6874;
      64315:data<=-16'd6701;
      64316:data<=-16'd7254;
      64317:data<=-16'd8082;
      64318:data<=-16'd9218;
      64319:data<=-16'd8478;
      64320:data<=-16'd8724;
      64321:data<=-16'd13688;
      64322:data<=-16'd17969;
      64323:data<=-16'd19255;
      64324:data<=-16'd19364;
      64325:data<=-16'd18089;
      64326:data<=-16'd17716;
      64327:data<=-16'd17302;
      64328:data<=-16'd15808;
      64329:data<=-16'd16478;
      64330:data<=-16'd16885;
      64331:data<=-16'd15687;
      64332:data<=-16'd15858;
      64333:data<=-16'd15593;
      64334:data<=-16'd14266;
      64335:data<=-16'd13866;
      64336:data<=-16'd14272;
      64337:data<=-16'd14521;
      64338:data<=-16'd13449;
      64339:data<=-16'd12583;
      64340:data<=-16'd12665;
      64341:data<=-16'd11694;
      64342:data<=-16'd10951;
      64343:data<=-16'd10837;
      64344:data<=-16'd10096;
      64345:data<=-16'd9596;
      64346:data<=-16'd8983;
      64347:data<=-16'd7997;
      64348:data<=-16'd5800;
      64349:data<=-16'd3149;
      64350:data<=-16'd3791;
      64351:data<=-16'd3987;
      64352:data<=-16'd2209;
      64353:data<=-16'd3084;
      64354:data<=16'd717;
      64355:data<=16'd10307;
      64356:data<=16'd12771;
      64357:data<=16'd10520;
      64358:data<=16'd10455;
      64359:data<=16'd9730;
      64360:data<=16'd10463;
      64361:data<=16'd12326;
      64362:data<=16'd11811;
      64363:data<=16'd12270;
      64364:data<=16'd12460;
      64365:data<=16'd10366;
      64366:data<=16'd11056;
      64367:data<=16'd13186;
      64368:data<=16'd12798;
      64369:data<=16'd12598;
      64370:data<=16'd12672;
      64371:data<=16'd11523;
      64372:data<=16'd11969;
      64373:data<=16'd14032;
      64374:data<=16'd14179;
      64375:data<=16'd12599;
      64376:data<=16'd12110;
      64377:data<=16'd12410;
      64378:data<=16'd11806;
      64379:data<=16'd12316;
      64380:data<=16'd14343;
      64381:data<=16'd13383;
      64382:data<=16'd10760;
      64383:data<=16'd11126;
      64384:data<=16'd11565;
      64385:data<=16'd11327;
      64386:data<=16'd13315;
      64387:data<=16'd12380;
      64388:data<=16'd5921;
      64389:data<=16'd531;
      64390:data<=-16'd822;
      64391:data<=16'd564;
      64392:data<=16'd2766;
      64393:data<=16'd3450;
      64394:data<=16'd4073;
      64395:data<=16'd5148;
      64396:data<=16'd4331;
      64397:data<=16'd3961;
      64398:data<=16'd5864;
      64399:data<=16'd6587;
      64400:data<=16'd5950;
      64401:data<=16'd6485;
      64402:data<=16'd6423;
      64403:data<=16'd4878;
      64404:data<=16'd5389;
      64405:data<=16'd7286;
      64406:data<=16'd7141;
      64407:data<=16'd7053;
      64408:data<=16'd7397;
      64409:data<=16'd6131;
      64410:data<=16'd6539;
      64411:data<=16'd8178;
      64412:data<=16'd7641;
      64413:data<=16'd7474;
      64414:data<=16'd7377;
      64415:data<=16'd6610;
      64416:data<=16'd7879;
      64417:data<=16'd8214;
      64418:data<=16'd7577;
      64419:data<=16'd8301;
      64420:data<=16'd6921;
      64421:data<=16'd8601;
      64422:data<=16'd16240;
      64423:data<=16'd18632;
      64424:data<=16'd16442;
      64425:data<=16'd16754;
      64426:data<=16'd16020;
      64427:data<=16'd14903;
      64428:data<=16'd15174;
      64429:data<=16'd14383;
      64430:data<=16'd14239;
      64431:data<=16'd14140;
      64432:data<=16'd13182;
      64433:data<=16'd13285;
      64434:data<=16'd12272;
      64435:data<=16'd11112;
      64436:data<=16'd12216;
      64437:data<=16'd12320;
      64438:data<=16'd11514;
      64439:data<=16'd11018;
      64440:data<=16'd9389;
      64441:data<=16'd8372;
      64442:data<=16'd8091;
      64443:data<=16'd7095;
      64444:data<=16'd7203;
      64445:data<=16'd7820;
      64446:data<=16'd6810;
      64447:data<=16'd5315;
      64448:data<=16'd3958;
      64449:data<=16'd2467;
      64450:data<=16'd2173;
      64451:data<=16'd2681;
      64452:data<=16'd2622;
      64453:data<=16'd2655;
      64454:data<=16'd153;
      64455:data<=-16'd6599;
      64456:data<=-16'd10780;
      64457:data<=-16'd10484;
      64458:data<=-16'd10654;
      64459:data<=-16'd10219;
      64460:data<=-16'd9900;
      64461:data<=-16'd12214;
      64462:data<=-16'd12790;
      64463:data<=-16'd11515;
      64464:data<=-16'd11662;
      64465:data<=-16'd11517;
      64466:data<=-16'd11612;
      64467:data<=-16'd12924;
      64468:data<=-16'd13438;
      64469:data<=-16'd13443;
      64470:data<=-16'd13480;
      64471:data<=-16'd12982;
      64472:data<=-16'd12510;
      64473:data<=-16'd12803;
      64474:data<=-16'd13317;
      64475:data<=-16'd12972;
      64476:data<=-16'd12919;
      64477:data<=-16'd13335;
      64478:data<=-16'd12549;
      64479:data<=-16'd12739;
      64480:data<=-16'd14634;
      64481:data<=-16'd14892;
      64482:data<=-16'd13718;
      64483:data<=-16'd12944;
      64484:data<=-16'd12854;
      64485:data<=-16'd13547;
      64486:data<=-16'd14965;
      64487:data<=-16'd15905;
      64488:data<=-16'd12101;
      64489:data<=-16'd4939;
      64490:data<=-16'd2840;
      64491:data<=-16'd4824;
      64492:data<=-16'd5850;
      64493:data<=-16'd7030;
      64494:data<=-16'd6816;
      64495:data<=-16'd5388;
      64496:data<=-16'd5932;
      64497:data<=-16'd5988;
      64498:data<=-16'd5770;
      64499:data<=-16'd7380;
      64500:data<=-16'd7673;
      64501:data<=-16'd6787;
      64502:data<=-16'd6478;
      64503:data<=-16'd5861;
      64504:data<=-16'd6587;
      64505:data<=-16'd8498;
      64506:data<=-16'd8769;
      64507:data<=-16'd8146;
      64508:data<=-16'd7906;
      64509:data<=-16'd8031;
      64510:data<=-16'd8739;
      64511:data<=-16'd9085;
      64512:data<=-16'd8545;
      64513:data<=-16'd7943;
      64514:data<=-16'd7667;
      64515:data<=-16'd7862;
      64516:data<=-16'd8031;
      64517:data<=-16'd7902;
      64518:data<=-16'd8229;
      64519:data<=-16'd7896;
      64520:data<=-16'd6810;
      64521:data<=-16'd8587;
      64522:data<=-16'd13000;
      64523:data<=-16'd16228;
      64524:data<=-16'd17567;
      64525:data<=-16'd17230;
      64526:data<=-16'd16190;
      64527:data<=-16'd15958;
      64528:data<=-16'd15168;
      64529:data<=-16'd14404;
      64530:data<=-16'd15195;
      64531:data<=-16'd14769;
      64532:data<=-16'd13097;
      64533:data<=-16'd13045;
      64534:data<=-16'd13391;
      64535:data<=-16'd13109;
      64536:data<=-16'd13439;
      64537:data<=-16'd13474;
      64538:data<=-16'd12075;
      64539:data<=-16'd10922;
      64540:data<=-16'd10880;
      64541:data<=-16'd10386;
      64542:data<=-16'd9743;
      64543:data<=-16'd9624;
      64544:data<=-16'd8825;
      64545:data<=-16'd8056;
      64546:data<=-16'd7902;
      64547:data<=-16'd7652;
      64548:data<=-16'd7130;
      64549:data<=-16'd4858;
      64550:data<=-16'd2946;
      64551:data<=-16'd3990;
      64552:data<=-16'd3750;
      64553:data<=-16'd2896;
      64554:data<=-16'd3488;
      64555:data<=16'd1192;
      64556:data<=16'd8674;
      64557:data<=16'd9879;
      64558:data<=16'd8463;
      64559:data<=16'd9153;
      64560:data<=16'd9677;
      64561:data<=16'd9721;
      64562:data<=16'd10132;
      64563:data<=16'd10284;
      64564:data<=16'd9856;
      64565:data<=16'd9652;
      64566:data<=16'd10019;
      64567:data<=16'd10416;
      64568:data<=16'd11203;
      64569:data<=16'd11568;
      64570:data<=16'd10957;
      64571:data<=16'd10854;
      64572:data<=16'd10545;
      64573:data<=16'd10279;
      64574:data<=16'd11418;
      64575:data<=16'd11787;
      64576:data<=16'd11245;
      64577:data<=16'd10875;
      64578:data<=16'd10293;
      64579:data<=16'd11098;
      64580:data<=16'd12279;
      64581:data<=16'd12052;
      64582:data<=16'd11784;
      64583:data<=16'd11119;
      64584:data<=16'd10625;
      64585:data<=16'd11062;
      64586:data<=16'd11655;
      64587:data<=16'd12962;
      64588:data<=16'd10928;
      64589:data<=16'd4687;
      64590:data<=16'd2096;
      64591:data<=16'd2532;
      64592:data<=16'd2353;
      64593:data<=16'd3979;
      64594:data<=16'd5039;
      64595:data<=16'd4546;
      64596:data<=16'd4883;
      64597:data<=16'd4294;
      64598:data<=16'd4379;
      64599:data<=16'd6376;
      64600:data<=16'd6704;
      64601:data<=16'd5890;
      64602:data<=16'd5416;
      64603:data<=16'd5001;
      64604:data<=16'd5636;
      64605:data<=16'd6728;
      64606:data<=16'd7186;
      64607:data<=16'd6968;
      64608:data<=16'd6499;
      64609:data<=16'd6385;
      64610:data<=16'd6270;
      64611:data<=16'd6849;
      64612:data<=16'd7758;
      64613:data<=16'd7160;
      64614:data<=16'd6708;
      64615:data<=16'd6787;
      64616:data<=16'd6243;
      64617:data<=16'd6567;
      64618:data<=16'd7084;
      64619:data<=16'd7397;
      64620:data<=16'd7498;
      64621:data<=16'd5789;
      64622:data<=16'd7699;
      64623:data<=16'd14819;
      64624:data<=16'd17318;
      64625:data<=16'd15180;
      64626:data<=16'd15107;
      64627:data<=16'd15013;
      64628:data<=16'd13797;
      64629:data<=16'd13661;
      64630:data<=16'd14183;
      64631:data<=16'd14474;
      64632:data<=16'd13720;
      64633:data<=16'd12715;
      64634:data<=16'd12226;
      64635:data<=16'd11538;
      64636:data<=16'd12158;
      64637:data<=16'd13267;
      64638:data<=16'd12184;
      64639:data<=16'd11092;
      64640:data<=16'd10928;
      64641:data<=16'd10354;
      64642:data<=16'd10378;
      64643:data<=16'd10056;
      64644:data<=16'd8610;
      64645:data<=16'd7909;
      64646:data<=16'd7837;
      64647:data<=16'd7855;
      64648:data<=16'd7206;
      64649:data<=16'd4869;
      64650:data<=16'd3733;
      64651:data<=16'd4529;
      64652:data<=16'd3656;
      64653:data<=16'd2770;
      64654:data<=16'd3480;
      64655:data<=16'd296;
      64656:data<=-16'd6173;
      64657:data<=-16'd8448;
      64658:data<=-16'd7705;
      64659:data<=-16'd8179;
      64660:data<=-16'd8123;
      64661:data<=-16'd8296;
      64662:data<=-16'd9790;
      64663:data<=-16'd9647;
      64664:data<=-16'd9133;
      64665:data<=-16'd9618;
      64666:data<=-16'd8774;
      64667:data<=-16'd8589;
      64668:data<=-16'd10185;
      64669:data<=-16'd10425;
      64670:data<=-16'd9832;
      64671:data<=-16'd9615;
      64672:data<=-16'd8998;
      64673:data<=-16'd9068;
      64674:data<=-16'd10123;
      64675:data<=-16'd10715;
      64676:data<=-16'd10555;
      64677:data<=-16'd10096;
      64678:data<=-16'd9712;
      64679:data<=-16'd9919;
      64680:data<=-16'd10801;
      64681:data<=-16'd11279;
      64682:data<=-16'd10809;
      64683:data<=-16'd10375;
      64684:data<=-16'd10210;
      64685:data<=-16'd9864;
      64686:data<=-16'd9586;
      64687:data<=-16'd10522;
      64688:data<=-16'd11784;
      64689:data<=-16'd8414;
      64690:data<=-16'd1724;
      64691:data<=-16'd59;
      64692:data<=-16'd2403;
      64693:data<=-16'd3119;
      64694:data<=-16'd3368;
      64695:data<=-16'd3617;
      64696:data<=-16'd3213;
      64697:data<=-16'd3280;
      64698:data<=-16'd3523;
      64699:data<=-16'd4232;
      64700:data<=-16'd4843;
      64701:data<=-16'd4416;
      64702:data<=-16'd4540;
      64703:data<=-16'd4601;
      64704:data<=-16'd4211;
      64705:data<=-16'd5283;
      64706:data<=-16'd6234;
      64707:data<=-16'd5900;
      64708:data<=-16'd5671;
      64709:data<=-16'd4965;
      64710:data<=-16'd4159;
      64711:data<=-16'd5084;
      64712:data<=-16'd6376;
      64713:data<=-16'd5814;
      64714:data<=-16'd4969;
      64715:data<=-16'd5379;
      64716:data<=-16'd5394;
      64717:data<=-16'd5301;
      64718:data<=-16'd6119;
      64719:data<=-16'd6543;
      64720:data<=-16'd6278;
      64721:data<=-16'd5421;
      64722:data<=-16'd6746;
      64723:data<=-16'd12469;
      64724:data<=-16'd15905;
      64725:data<=-16'd14689;
      64726:data<=-16'd14415;
      64727:data<=-16'd14117;
      64728:data<=-16'd12669;
      64729:data<=-16'd12355;
      64730:data<=-16'd12469;
      64731:data<=-16'd12883;
      64732:data<=-16'd12700;
      64733:data<=-16'd11773;
      64734:data<=-16'd11691;
      64735:data<=-16'd10768;
      64736:data<=-16'd10354;
      64737:data<=-16'd11492;
      64738:data<=-16'd10739;
      64739:data<=-16'd9909;
      64740:data<=-16'd9878;
      64741:data<=-16'd8862;
      64742:data<=-16'd8942;
      64743:data<=-16'd8745;
      64744:data<=-16'd7623;
      64745:data<=-16'd7624;
      64746:data<=-16'd6966;
      64747:data<=-16'd6454;
      64748:data<=-16'd6273;
      64749:data<=-16'd4244;
      64750:data<=-16'd2886;
      64751:data<=-16'd2793;
      64752:data<=-16'd2544;
      64753:data<=-16'd2206;
      64754:data<=-16'd1665;
      64755:data<=-16'd1377;
      64756:data<=16'd2617;
      64757:data<=16'd9530;
      64758:data<=16'd10646;
      64759:data<=16'd8925;
      64760:data<=16'd9500;
      64761:data<=16'd9506;
      64762:data<=16'd10419;
      64763:data<=16'd11279;
      64764:data<=16'd10091;
      64765:data<=16'd10052;
      64766:data<=16'd9949;
      64767:data<=16'd10108;
      64768:data<=16'd11967;
      64769:data<=16'd11791;
      64770:data<=16'd10818;
      64771:data<=16'd10944;
      64772:data<=16'd10416;
      64773:data<=16'd10527;
      64774:data<=16'd11374;
      64775:data<=16'd11878;
      64776:data<=16'd11958;
      64777:data<=16'd11368;
      64778:data<=16'd11092;
      64779:data<=16'd10748;
      64780:data<=16'd10719;
      64781:data<=16'd11978;
      64782:data<=16'd12239;
      64783:data<=16'd11539;
      64784:data<=16'd10957;
      64785:data<=16'd10301;
      64786:data<=16'd10757;
      64787:data<=16'd11650;
      64788:data<=16'd12076;
      64789:data<=16'd9882;
      64790:data<=16'd3753;
      64791:data<=16'd625;
      64792:data<=16'd2249;
      64793:data<=16'd3243;
      64794:data<=16'd4135;
      64795:data<=16'd4411;
      64796:data<=16'd3603;
      64797:data<=16'd4009;
      64798:data<=16'd3929;
      64799:data<=16'd4405;
      64800:data<=16'd5977;
      64801:data<=16'd5503;
      64802:data<=16'd5092;
      64803:data<=16'd5112;
      64804:data<=16'd4434;
      64805:data<=16'd5492;
      64806:data<=16'd6437;
      64807:data<=16'd5906;
      64808:data<=16'd5841;
      64809:data<=16'd5742;
      64810:data<=16'd5377;
      64811:data<=16'd5274;
      64812:data<=16'd5994;
      64813:data<=16'd6492;
      64814:data<=16'd5624;
      64815:data<=16'd5799;
      64816:data<=16'd6032;
      64817:data<=16'd5383;
      64818:data<=16'd6404;
      64819:data<=16'd6734;
      64820:data<=16'd6554;
      64821:data<=16'd6919;
      64822:data<=16'd5244;
      64823:data<=16'd7711;
      64824:data<=16'd14803;
      64825:data<=16'd16242;
      64826:data<=16'd14289;
      64827:data<=16'd14257;
      64828:data<=16'd13559;
      64829:data<=16'd12340;
      64830:data<=16'd12322;
      64831:data<=16'd13298;
      64832:data<=16'd13068;
      64833:data<=16'd11661;
      64834:data<=16'd11552;
      64835:data<=16'd10777;
      64836:data<=16'd10205;
      64837:data<=16'd11715;
      64838:data<=16'd11373;
      64839:data<=16'd10445;
      64840:data<=16'd10379;
      64841:data<=16'd8933;
      64842:data<=16'd8787;
      64843:data<=16'd9294;
      64844:data<=16'd8528;
      64845:data<=16'd8478;
      64846:data<=16'd7844;
      64847:data<=16'd6931;
      64848:data<=16'd6545;
      64849:data<=16'd4969;
      64850:data<=16'd3630;
      64851:data<=16'd3081;
      64852:data<=16'd2992;
      64853:data<=16'd2764;
      64854:data<=16'd1715;
      64855:data<=16'd1871;
      64856:data<=-16'd1098;
      64857:data<=-16'd8278;
      64858:data<=-16'd10266;
      64859:data<=-16'd8886;
      64860:data<=-16'd9411;
      64861:data<=-16'd9291;
      64862:data<=-16'd10116;
      64863:data<=-16'd10807;
      64864:data<=-16'd9931;
      64865:data<=-16'd10601;
      64866:data<=-16'd10295;
      64867:data<=-16'd9621;
      64868:data<=-16'd11075;
      64869:data<=-16'd11166;
      64870:data<=-16'd10847;
      64871:data<=-16'd11133;
      64872:data<=-16'd10401;
      64873:data<=-16'd10248;
      64874:data<=-16'd10727;
      64875:data<=-16'd11638;
      64876:data<=-16'd12181;
      64877:data<=-16'd11552;
      64878:data<=-16'd11764;
      64879:data<=-16'd11330;
      64880:data<=-16'd10812;
      64881:data<=-16'd12266;
      64882:data<=-16'd12082;
      64883:data<=-16'd11700;
      64884:data<=-16'd12264;
      64885:data<=-16'd10901;
      64886:data<=-16'd11089;
      64887:data<=-16'd12234;
      64888:data<=-16'd12188;
      64889:data<=-16'd12690;
      64890:data<=-16'd8570;
      64891:data<=-16'd1947;
      64892:data<=-16'd1764;
      64893:data<=-16'd4175;
      64894:data<=-16'd4620;
      64895:data<=-16'd4531;
      64896:data<=-16'd4256;
      64897:data<=-16'd4267;
      64898:data<=-16'd3990;
      64899:data<=-16'd4426;
      64900:data<=-16'd5847;
      64901:data<=-16'd5711;
      64902:data<=-16'd5653;
      64903:data<=-16'd5956;
      64904:data<=-16'd5128;
      64905:data<=-16'd5635;
      64906:data<=-16'd6736;
      64907:data<=-16'd6631;
      64908:data<=-16'd6341;
      64909:data<=-16'd5680;
      64910:data<=-16'd5162;
      64911:data<=-16'd5362;
      64912:data<=-16'd6114;
      64913:data<=-16'd6737;
      64914:data<=-16'd6141;
      64915:data<=-16'd5968;
      64916:data<=-16'd5964;
      64917:data<=-16'd5371;
      64918:data<=-16'd6429;
      64919:data<=-16'd7007;
      64920:data<=-16'd6666;
      64921:data<=-16'd7057;
      64922:data<=-16'd5307;
      64923:data<=-16'd6441;
      64924:data<=-16'd13515;
      64925:data<=-16'd16365;
      64926:data<=-16'd14542;
      64927:data<=-16'd14498;
      64928:data<=-16'd13976;
      64929:data<=-16'd12513;
      64930:data<=-16'd12696;
      64931:data<=-16'd13737;
      64932:data<=-16'd13634;
      64933:data<=-16'd12427;
      64934:data<=-16'd12041;
      64935:data<=-16'd11558;
      64936:data<=-16'd10887;
      64937:data<=-16'd11952;
      64938:data<=-16'd11970;
      64939:data<=-16'd10502;
      64940:data<=-16'd10398;
      64941:data<=-16'd10211;
      64942:data<=-16'd9694;
      64943:data<=-16'd9639;
      64944:data<=-16'd9092;
      64945:data<=-16'd8522;
      64946:data<=-16'd7597;
      64947:data<=-16'd6792;
      64948:data<=-16'd6983;
      64949:data<=-16'd6112;
      64950:data<=-16'd4637;
      64951:data<=-16'd4185;
      64952:data<=-16'd3761;
      64953:data<=-16'd3213;
      64954:data<=-16'd2737;
      64955:data<=-16'd2582;
      64956:data<=-16'd1533;
      64957:data<=16'd3237;
      64958:data<=16'd8460;
      64959:data<=16'd9025;
      64960:data<=16'd7630;
      64961:data<=16'd8231;
      64962:data<=16'd9643;
      64963:data<=16'd9917;
      64964:data<=16'd9599;
      64965:data<=16'd9471;
      64966:data<=16'd9018;
      64967:data<=16'd8542;
      64968:data<=16'd9127;
      64969:data<=16'd10301;
      64970:data<=16'd10587;
      64971:data<=16'd10022;
      64972:data<=16'd9632;
      64973:data<=16'd9282;
      64974:data<=16'd9589;
      64975:data<=16'd10790;
      64976:data<=16'd10842;
      64977:data<=16'd10698;
      64978:data<=16'd10951;
      64979:data<=16'd9498;
      64980:data<=16'd9407;
      64981:data<=16'd11435;
      64982:data<=16'd11394;
      64983:data<=16'd10950;
      64984:data<=16'd10768;
      64985:data<=16'd9643;
      64986:data<=16'd10143;
      64987:data<=16'd10501;
      64988:data<=16'd10311;
      64989:data<=16'd11775;
      64990:data<=16'd9151;
      64991:data<=16'd2361;
      64992:data<=-16'd23;
      64993:data<=16'd1865;
      64994:data<=16'd3080;
      64995:data<=16'd2857;
      64996:data<=16'd2714;
      64997:data<=16'd3090;
      64998:data<=16'd2663;
      64999:data<=16'd2840;
      65000:data<=16'd4405;
      65001:data<=16'd4655;
      65002:data<=16'd4269;
      65003:data<=16'd4278;
      65004:data<=16'd3765;
      65005:data<=16'd4232;
      65006:data<=16'd5480;
      65007:data<=16'd5817;
      65008:data<=16'd5733;
      65009:data<=16'd5395;
      65010:data<=16'd4819;
      65011:data<=16'd4695;
      65012:data<=16'd5724;
      65013:data<=16'd6921;
      65014:data<=16'd6263;
      65015:data<=16'd5529;
      65016:data<=16'd5674;
      65017:data<=16'd4839;
      65018:data<=16'd5060;
      65019:data<=16'd6331;
      65020:data<=16'd6179;
      65021:data<=16'd6401;
      65022:data<=16'd5903;
      65023:data<=16'd4902;
      65024:data<=16'd9306;
      65025:data<=16'd15391;
      65026:data<=16'd15685;
      65027:data<=16'd13820;
      65028:data<=16'd13618;
      65029:data<=16'd13245;
      65030:data<=16'd12910;
      65031:data<=16'd13620;
      65032:data<=16'd13706;
      65033:data<=16'd12501;
      65034:data<=16'd11875;
      65035:data<=16'd11776;
      65036:data<=16'd11227;
      65037:data<=16'd11473;
      65038:data<=16'd11958;
      65039:data<=16'd11411;
      65040:data<=16'd10928;
      65041:data<=16'd10284;
      65042:data<=16'd9251;
      65043:data<=16'd8983;
      65044:data<=16'd9000;
      65045:data<=16'd8492;
      65046:data<=16'd7403;
      65047:data<=16'd6680;
      65048:data<=16'd6868;
      65049:data<=16'd6105;
      65050:data<=16'd4613;
      65051:data<=16'd3889;
      65052:data<=16'd3284;
      65053:data<=16'd3115;
      65054:data<=16'd2628;
      65055:data<=16'd1650;
      65056:data<=16'd1817;
      65057:data<=-16'd1266;
      65058:data<=-16'd8032;
      65059:data<=-16'd10088;
      65060:data<=-16'd8366;
      65061:data<=-16'd8520;
      65062:data<=-16'd9406;
      65063:data<=-16'd10296;
      65064:data<=-16'd10551;
      65065:data<=-16'd9841;
      65066:data<=-16'd9908;
      65067:data<=-16'd9567;
      65068:data<=-16'd9345;
      65069:data<=-16'd10666;
      65070:data<=-16'd10980;
      65071:data<=-16'd10655;
      65072:data<=-16'd10511;
      65073:data<=-16'd9386;
      65074:data<=-16'd9618;
      65075:data<=-16'd10980;
      65076:data<=-16'd10784;
      65077:data<=-16'd10477;
      65078:data<=-16'd10399;
      65079:data<=-16'd9371;
      65080:data<=-16'd8969;
      65081:data<=-16'd10163;
      65082:data<=-16'd11200;
      65083:data<=-16'd10836;
      65084:data<=-16'd10340;
      65085:data<=-16'd10149;
      65086:data<=-16'd9709;
      65087:data<=-16'd10110;
      65088:data<=-16'd10818;
      65089:data<=-16'd10983;
      65090:data<=-16'd10229;
      65091:data<=-16'd5598;
      65092:data<=-16'd153;
      65093:data<=-16'd654;
      65094:data<=-16'd3428;
      65095:data<=-16'd3477;
      65096:data<=-16'd3098;
      65097:data<=-16'd2952;
      65098:data<=-16'd2405;
      65099:data<=-16'd2892;
      65100:data<=-16'd4314;
      65101:data<=-16'd5013;
      65102:data<=-16'd4504;
      65103:data<=-16'd3935;
      65104:data<=-16'd3751;
      65105:data<=-16'd3739;
      65106:data<=-16'd4589;
      65107:data<=-16'd5577;
      65108:data<=-16'd5483;
      65109:data<=-16'd5231;
      65110:data<=-16'd5046;
      65111:data<=-16'd4419;
      65112:data<=-16'd4761;
      65113:data<=-16'd6314;
      65114:data<=-16'd6614;
      65115:data<=-16'd5708;
      65116:data<=-16'd5316;
      65117:data<=-16'd4749;
      65118:data<=-16'd5071;
      65119:data<=-16'd6569;
      65120:data<=-16'd6000;
      65121:data<=-16'd5626;
      65122:data<=-16'd6514;
      65123:data<=-16'd4736;
      65124:data<=-16'd6234;
      65125:data<=-16'd13649;
      65126:data<=-16'd16196;
      65127:data<=-16'd13907;
      65128:data<=-16'd13978;
      65129:data<=-16'd13796;
      65130:data<=-16'd12354;
      65131:data<=-16'd12543;
      65132:data<=-16'd13197;
      65133:data<=-16'd12900;
      65134:data<=-16'd12387;
      65135:data<=-16'd12076;
      65136:data<=-16'd11342;
      65137:data<=-16'd10978;
      65138:data<=-16'd11866;
      65139:data<=-16'd11891;
      65140:data<=-16'd10845;
      65141:data<=-16'd10370;
      65142:data<=-16'd9811;
      65143:data<=-16'd9180;
      65144:data<=-16'd8674;
      65145:data<=-16'd7908;
      65146:data<=-16'd7395;
      65147:data<=-16'd6884;
      65148:data<=-16'd6587;
      65149:data<=-16'd6231;
      65150:data<=-16'd4640;
      65151:data<=-16'd3180;
      65152:data<=-16'd2689;
      65153:data<=-16'd2570;
      65154:data<=-16'd2470;
      65155:data<=-16'd1603;
      65156:data<=-16'd896;
      65157:data<=16'd876;
      65158:data<=16'd6084;
      65159:data<=16'd10367;
      65160:data<=16'd10615;
      65161:data<=16'd9961;
      65162:data<=16'd10478;
      65163:data<=16'd11735;
      65164:data<=16'd11929;
      65165:data<=16'd11333;
      65166:data<=16'd11347;
      65167:data<=16'd10713;
      65168:data<=16'd10771;
      65169:data<=16'd12311;
      65170:data<=16'd12522;
      65171:data<=16'd12199;
      65172:data<=16'd11928;
      65173:data<=16'd11060;
      65174:data<=16'd11203;
      65175:data<=16'd11684;
      65176:data<=16'd12029;
      65177:data<=16'd12377;
      65178:data<=16'd11768;
      65179:data<=16'd11295;
      65180:data<=16'd10721;
      65181:data<=16'd10819;
      65182:data<=16'd12640;
      65183:data<=16'd12604;
      65184:data<=16'd11935;
      65185:data<=16'd12187;
      65186:data<=16'd10745;
      65187:data<=16'd11127;
      65188:data<=16'd12515;
      65189:data<=16'd11602;
      65190:data<=16'd12511;
      65191:data<=16'd10481;
      65192:data<=16'd3015;
      65193:data<=16'd1307;
      65194:data<=16'd4431;
      65195:data<=16'd4438;
      65196:data<=16'd3755;
      65197:data<=16'd4188;
      65198:data<=16'd4109;
      65199:data<=16'd3662;
      65200:data<=16'd4272;
      65201:data<=16'd5668;
      65202:data<=16'd5564;
      65203:data<=16'd5328;
      65204:data<=16'd5595;
      65205:data<=16'd4441;
      65206:data<=16'd4672;
      65207:data<=16'd6725;
      65208:data<=16'd6996;
      65209:data<=16'd6402;
      65210:data<=16'd6106;
      65211:data<=16'd5601;
      65212:data<=16'd5996;
      65213:data<=16'd7294;
      65214:data<=16'd7600;
      65215:data<=16'd6590;
      65216:data<=16'd6120;
      65217:data<=16'd5862;
      65218:data<=16'd5492;
      65219:data<=16'd6745;
      65220:data<=16'd7206;
      65221:data<=16'd6313;
      65222:data<=16'd6934;
      65223:data<=16'd6185;
      65224:data<=16'd5820;
      65225:data<=16'd11210;
      65226:data<=16'd16072;
      65227:data<=16'd15553;
      65228:data<=16'd14386;
      65229:data<=16'd14088;
      65230:data<=16'd13182;
      65231:data<=16'd12956;
      65232:data<=16'd14325;
      65233:data<=16'd14452;
      65234:data<=16'd12645;
      65235:data<=16'd12192;
      65236:data<=16'd12023;
      65237:data<=16'd11429;
      65238:data<=16'd12533;
      65239:data<=16'd12519;
      65240:data<=16'd11241;
      65241:data<=16'd11065;
      65242:data<=16'd10082;
      65243:data<=16'd9347;
      65244:data<=16'd9244;
      65245:data<=16'd8152;
      65246:data<=16'd8002;
      65247:data<=16'd7538;
      65248:data<=16'd6431;
      65249:data<=16'd6780;
      65250:data<=16'd5635;
      65251:data<=16'd3518;
      65252:data<=16'd2892;
      65253:data<=16'd2184;
      65254:data<=16'd2103;
      65255:data<=16'd1745;
      65256:data<=16'd487;
      65257:data<=16'd300;
      65258:data<=-16'd2964;
      65259:data<=-16'd9204;
      65260:data<=-16'd10868;
      65261:data<=-16'd9395;
      65262:data<=-16'd10146;
      65263:data<=-16'd11771;
      65264:data<=-16'd11809;
      65265:data<=-16'd11173;
      65266:data<=-16'd11254;
      65267:data<=-16'd11118;
      65268:data<=-16'd10884;
      65269:data<=-16'd11831;
      65270:data<=-16'd12399;
      65271:data<=-16'd11916;
      65272:data<=-16'd11853;
      65273:data<=-16'd11887;
      65274:data<=-16'd11165;
      65275:data<=-16'd10921;
      65276:data<=-16'd12117;
      65277:data<=-16'd12652;
      65278:data<=-16'd12161;
      65279:data<=-16'd12151;
      65280:data<=-16'd11103;
      65281:data<=-16'd10827;
      65282:data<=-16'd12901;
      65283:data<=-16'd12740;
      65284:data<=-16'd11867;
      65285:data<=-16'd12380;
      65286:data<=-16'd10928;
      65287:data<=-16'd10998;
      65288:data<=-16'd12904;
      65289:data<=-16'd12013;
      65290:data<=-16'd11858;
      65291:data<=-16'd11098;
      65292:data<=-16'd5526;
      65293:data<=-16'd1698;
      65294:data<=-16'd2790;
      65295:data<=-16'd4238;
      65296:data<=-16'd4131;
      65297:data<=-16'd3956;
      65298:data<=-16'd4466;
      65299:data<=-16'd3823;
      65300:data<=-16'd3830;
      65301:data<=-16'd6132;
      65302:data<=-16'd6185;
      65303:data<=-16'd5150;
      65304:data<=-16'd5768;
      65305:data<=-16'd5019;
      65306:data<=-16'd5065;
      65307:data<=-16'd6731;
      65308:data<=-16'd6290;
      65309:data<=-16'd5937;
      65310:data<=-16'd6398;
      65311:data<=-16'd5777;
      65312:data<=-16'd5674;
      65313:data<=-16'd6261;
      65314:data<=-16'd6813;
      65315:data<=-16'd6760;
      65316:data<=-16'd6249;
      65317:data<=-16'd6561;
      65318:data<=-16'd6126;
      65319:data<=-16'd6084;
      65320:data<=-16'd7811;
      65321:data<=-16'd7365;
      65322:data<=-16'd6740;
      65323:data<=-16'd7053;
      65324:data<=-16'd4886;
      65325:data<=-16'd7668;
      65326:data<=-16'd15850;
      65327:data<=-16'd17138;
      65328:data<=-16'd14559;
      65329:data<=-16'd15079;
      65330:data<=-16'd14536;
      65331:data<=-16'd13740;
      65332:data<=-16'd14775;
      65333:data<=-16'd14587;
      65334:data<=-16'd13509;
      65335:data<=-16'd12819;
      65336:data<=-16'd12339;
      65337:data<=-16'd12366;
      65338:data<=-16'd12342;
      65339:data<=-16'd12284;
      65340:data<=-16'd12296;
      65341:data<=-16'd11620;
      65342:data<=-16'd10705;
      65343:data<=-16'd10252;
      65344:data<=-16'd9932;
      65345:data<=-16'd9538;
      65346:data<=-16'd9194;
      65347:data<=-16'd8492;
      65348:data<=-16'd7612;
      65349:data<=-16'd7418;
      65350:data<=-16'd6537;
      65351:data<=-16'd4552;
      65352:data<=-16'd3773;
      65353:data<=-16'd3548;
      65354:data<=-16'd3048;
      65355:data<=-16'd2949;
      65356:data<=-16'd1826;
      65357:data<=-16'd614;
      65358:data<=16'd980;
      65359:data<=16'd5993;
      65360:data<=16'd9758;
      65361:data<=16'd9110;
      65362:data<=16'd9182;
      65363:data<=16'd10349;
      65364:data<=16'd10615;
      65365:data<=16'd10742;
      65366:data<=16'd10416;
      65367:data<=16'd10087;
      65368:data<=16'd9632;
      65369:data<=16'd9389;
      65370:data<=16'd10690;
      65371:data<=16'd11071;
      65372:data<=16'd10410;
      65373:data<=16'd10481;
      65374:data<=16'd9596;
      65375:data<=16'd9630;
      65376:data<=16'd11315;
      65377:data<=16'd11038;
      65378:data<=16'd10527;
      65379:data<=16'd10881;
      65380:data<=16'd9912;
      65381:data<=16'd9758;
      65382:data<=16'd11265;
      65383:data<=16'd11603;
      65384:data<=16'd10712;
      65385:data<=16'd10540;
      65386:data<=16'd10460;
      65387:data<=16'd9644;
      65388:data<=16'd10310;
      65389:data<=16'd11130;
      65390:data<=16'd10299;
      65391:data<=16'd11142;
      65392:data<=16'd9192;
      65393:data<=16'd1507;
      65394:data<=-16'd335;
      65395:data<=16'd3626;
      65396:data<=16'd3160;
      65397:data<=16'd2044;
      65398:data<=16'd3057;
      65399:data<=16'd2447;
      65400:data<=16'd2705;
      65401:data<=16'd4253;
      65402:data<=16'd4344;
      65403:data<=16'd4202;
      65404:data<=16'd4399;
      65405:data<=16'd4181;
      65406:data<=16'd4068;
      65407:data<=16'd4687;
      65408:data<=16'd5635;
      65409:data<=16'd5777;
      65410:data<=16'd5392;
      65411:data<=16'd5028;
      65412:data<=16'd4240;
      65413:data<=16'd4344;
      65414:data<=16'd5984;
      65415:data<=16'd6423;
      65416:data<=16'd5328;
      65417:data<=16'd4963;
      65418:data<=16'd4664;
      65419:data<=16'd4761;
      65420:data<=16'd6272;
      65421:data<=16'd6037;
      65422:data<=16'd5075;
      65423:data<=16'd5932;
      65424:data<=16'd4963;
      65425:data<=16'd5736;
      65426:data<=16'd12431;
      65427:data<=16'd15982;
      65428:data<=16'd14468;
      65429:data<=16'd14348;
      65430:data<=16'd13878;
      65431:data<=16'd12704;
      65432:data<=16'd13273;
      65433:data<=16'd13694;
      65434:data<=16'd13312;
      65435:data<=16'd12574;
      65436:data<=16'd11661;
      65437:data<=16'd11065;
      65438:data<=16'd10919;
      65439:data<=16'd11856;
      65440:data<=16'd11943;
      65441:data<=16'd10292;
      65442:data<=16'd9785;
      65443:data<=16'd9734;
      65444:data<=16'd8846;
      65445:data<=16'd8264;
      65446:data<=16'd7764;
      65447:data<=16'd7512;
      65448:data<=16'd7294;
      65449:data<=16'd6760;
      65450:data<=16'd5830;
      65451:data<=16'd3711;
      65452:data<=16'd2830;
      65453:data<=16'd3260;
      65454:data<=16'd2397;
      65455:data<=16'd2426;
      65456:data<=16'd1905;
      65457:data<=-16'd244;
      65458:data<=16'd30;
      65459:data<=-16'd2367;
      65460:data<=-16'd9239;
      65461:data<=-16'd11150;
      65462:data<=-16'd9370;
      65463:data<=-16'd10392;
      65464:data<=-16'd11964;
      65465:data<=-16'd11714;
      65466:data<=-16'd10881;
      65467:data<=-16'd10718;
      65468:data<=-16'd10439;
      65469:data<=-16'd10240;
      65470:data<=-16'd11624;
      65471:data<=-16'd12035;
      65472:data<=-16'd10944;
      65473:data<=-16'd10953;
      65474:data<=-16'd10683;
      65475:data<=-16'd10398;
      65476:data<=-16'd11301;
      65477:data<=-16'd11276;
      65478:data<=-16'd10800;
      65479:data<=-16'd11151;
      65480:data<=-16'd11229;
      65481:data<=-16'd10630;
      65482:data<=-16'd10693;
      65483:data<=-16'd11972;
      65484:data<=-16'd12005;
      65485:data<=-16'd11179;
      65486:data<=-16'd11160;
      65487:data<=-16'd10038;
      65488:data<=-16'd10320;
      65489:data<=-16'd12289;
      65490:data<=-16'd11368;
      65491:data<=-16'd11171;
      65492:data<=-16'd10329;
      65493:data<=-16'd3762;
      65494:data<=-16'd669;
      65495:data<=-16'd3198;
      65496:data<=-16'd3075;
      65497:data<=-16'd2493;
      65498:data<=-16'd3187;
      65499:data<=-16'd2890;
      65500:data<=-16'd3200;
      65501:data<=-16'd3841;
      65502:data<=-16'd4247;
      65503:data<=-16'd4535;
      65504:data<=-16'd4284;
      65505:data<=-16'd4250;
      65506:data<=-16'd3626;
      65507:data<=-16'd3758;
      65508:data<=-16'd5900;
      65509:data<=-16'd6135;
      65510:data<=-16'd5154;
      65511:data<=-16'd5463;
      65512:data<=-16'd4780;
      65513:data<=-16'd4363;
      65514:data<=-16'd5609;
      65515:data<=-16'd5782;
      65516:data<=-16'd5096;
      65517:data<=-16'd5087;
      65518:data<=-16'd4965;
      65519:data<=-16'd4687;
      65520:data<=-16'd5509;
      65521:data<=-16'd6164;
      65522:data<=-16'd5221;
      65523:data<=-16'd5457;
      65524:data<=-16'd5624;
      65525:data<=-16'd3507;
      65526:data<=-16'd6604;
      65527:data<=-16'd14252;
      65528:data<=-16'd15526;
      65529:data<=-16'd13380;
      65530:data<=-16'd13725;
      65531:data<=-16'd13007;
      65532:data<=-16'd12410;
      65533:data<=-16'd13385;
      65534:data<=-16'd12747;
      65535:data<=-16'd11864;
      65536:data<=-16'd11781;
      65537:data<=-16'd10965;
      65538:data<=-16'd10828;
      65539:data<=-16'd11514;
      65540:data<=-16'd11294;
      65541:data<=-16'd10549;
      65542:data<=-16'd9761;
      65543:data<=-16'd8790;
      65544:data<=-16'd8025;
      65545:data<=-16'd7573;
      65546:data<=-16'd7448;
      65547:data<=-16'd7420;
      65548:data<=-16'd6722;
      65549:data<=-16'd5900;
      65550:data<=-16'd5509;
      65551:data<=-16'd4290;
      65552:data<=-16'd2866;
      65553:data<=-16'd2517;
      65554:data<=-16'd1985;
      65555:data<=-16'd1689;
      65556:data<=-16'd1715;
      65557:data<=-16'd235;
      65558:data<=16'd886;
      65559:data<=16'd2598;
      65560:data<=16'd8191;
      65561:data<=16'd11846;
      65562:data<=16'd10619;
      65563:data<=16'd10853;
      65564:data<=16'd12543;
      65565:data<=16'd12454;
      65566:data<=16'd12085;
      65567:data<=16'd11878;
      65568:data<=16'd11544;
      65569:data<=16'd11618;
      65570:data<=16'd12195;
      65571:data<=16'd12845;
      65572:data<=16'd12449;
      65573:data<=16'd12119;
      65574:data<=16'd12243;
      65575:data<=16'd11126;
      65576:data<=16'd11236;
      65577:data<=16'd12928;
      65578:data<=16'd12427;
      65579:data<=16'd11641;
      65580:data<=16'd12155;
      65581:data<=16'd11749;
      65582:data<=16'd11923;
      65583:data<=16'd13107;
      65584:data<=16'd12850;
      65585:data<=16'd12316;
      65586:data<=16'd12522;
      65587:data<=16'd11650;
      65588:data<=16'd11267;
      65589:data<=16'd13082;
      65590:data<=16'd13074;
      65591:data<=16'd11855;
      65592:data<=16'd13153;
      65593:data<=16'd10267;
      65594:data<=16'd2946;
      65595:data<=16'd2416;
      65596:data<=16'd5295;
      65597:data<=16'd4404;
      65598:data<=16'd4402;
      65599:data<=16'd4639;
      65600:data<=16'd3277;
      65601:data<=16'd4253;
      65602:data<=16'd5720;
      65603:data<=16'd5524;
      65604:data<=16'd5498;
      65605:data<=16'd5404;
      65606:data<=16'd5131;
      65607:data<=16'd5526;
      65608:data<=16'd6731;
      65609:data<=16'd7462;
      65610:data<=16'd7018;
      65611:data<=16'd7154;
      65612:data<=16'd7036;
      65613:data<=16'd6108;
      65614:data<=16'd6919;
      65615:data<=16'd7771;
      65616:data<=16'd7142;
      65617:data<=16'd7065;
      65618:data<=16'd6648;
      65619:data<=16'd5929;
      65620:data<=16'd7074;
      65621:data<=16'd8219;
      65622:data<=16'd7177;
      65623:data<=16'd6555;
      65624:data<=16'd7057;
      65625:data<=16'd5711;
      65626:data<=16'd7200;
      65627:data<=16'd14509;
      65628:data<=16'd17352;
      65629:data<=16'd14904;
      65630:data<=16'd15048;
      65631:data<=16'd14516;
      65632:data<=16'd13590;
      65633:data<=16'd15270;
      65634:data<=16'd14662;
      65635:data<=16'd13532;
      65636:data<=16'd14038;
      65637:data<=16'd12830;
      65638:data<=16'd12407;
      65639:data<=16'd13248;
      65640:data<=16'd12933;
      65641:data<=16'd12537;
      65642:data<=16'd11606;
      65643:data<=16'd10671;
      65644:data<=16'd10519;
      65645:data<=16'd9777;
      65646:data<=16'd9039;
      65647:data<=16'd8540;
      65648:data<=16'd8167;
      65649:data<=16'd8053;
      65650:data<=16'd7371;
      65651:data<=16'd6270;
      65652:data<=16'd4649;
      65653:data<=16'd3717;
      65654:data<=16'd3706;
      65655:data<=16'd2784;
      65656:data<=16'd3072;
      65657:data<=16'd2719;
      65658:data<=16'd3;
      65659:data<=16'd385;
      65660:data<=-16'd1510;
      65661:data<=-16'd8614;
      65662:data<=-16'd9908;
      65663:data<=-16'd8335;
      65664:data<=-16'd10381;
      65665:data<=-16'd10857;
      65666:data<=-16'd10413;
      65667:data<=-16'd10520;
      65668:data<=-16'd9902;
      65669:data<=-16'd10020;
      65670:data<=-16'd10270;
      65671:data<=-16'd11229;
      65672:data<=-16'd11749;
      65673:data<=-16'd10373;
      65674:data<=-16'd10652;
      65675:data<=-16'd10683;
      65676:data<=-16'd9650;
      65677:data<=-16'd10985;
      65678:data<=-16'd11059;
      65679:data<=-16'd9988;
      65680:data<=-16'd10574;
      65681:data<=-16'd10003;
      65682:data<=-16'd9894;
      65683:data<=-16'd11291;
      65684:data<=-16'd11450;
      65685:data<=-16'd11242;
      65686:data<=-16'd11089;
      65687:data<=-16'd10428;
      65688:data<=-16'd9887;
      65689:data<=-16'd10662;
      65690:data<=-16'd11928;
      65691:data<=-16'd11368;
      65692:data<=-16'd11605;
      65693:data<=-16'd10188;
      65694:data<=-16'd3039;
      65695:data<=-16'd514;
      65696:data<=-16'd3908;
      65697:data<=-16'd3438;
      65698:data<=-16'd3221;
      65699:data<=-16'd4435;
      65700:data<=-16'd2980;
      65701:data<=-16'd3374;
      65702:data<=-16'd4869;
      65703:data<=-16'd4637;
      65704:data<=-16'd4766;
      65705:data<=-16'd4752;
      65706:data<=-16'd4584;
      65707:data<=-16'd4651;
      65708:data<=-16'd5347;
      65709:data<=-16'd6684;
      65710:data<=-16'd6275;
      65711:data<=-16'd5859;
      65712:data<=-16'd6149;
      65713:data<=-16'd5418;
      65714:data<=-16'd6569;
      65715:data<=-16'd7899;
      65716:data<=-16'd6851;
      65717:data<=-16'd6796;
      65718:data<=-16'd6760;
      65719:data<=-16'd5799;
      65720:data<=-16'd6264;
      65721:data<=-16'd7532;
      65722:data<=-16'd8058;
      65723:data<=-16'd7301;
      65724:data<=-16'd6975;
      65725:data<=-16'd6593;
      65726:data<=-16'd5617;
      65727:data<=-16'd10081;
      65728:data<=-16'd16656;
      65729:data<=-16'd16747;
      65730:data<=-16'd15159;
      65731:data<=-16'd14794;
      65732:data<=-16'd14114;
      65733:data<=-16'd15318;
      65734:data<=-16'd15531;
      65735:data<=-16'd14126;
      65736:data<=-16'd13982;
      65737:data<=-16'd13259;
      65738:data<=-16'd12745;
      65739:data<=-16'd13373;
      65740:data<=-16'd13280;
      65741:data<=-16'd12822;
      65742:data<=-16'd12119;
      65743:data<=-16'd11568;
      65744:data<=-16'd11083;
      65745:data<=-16'd10087;
      65746:data<=-16'd9893;
      65747:data<=-16'd9509;
      65748:data<=-16'd8429;
      65749:data<=-16'd7982;
      65750:data<=-16'd7460;
      65751:data<=-16'd6781;
      65752:data<=-16'd5457;
      65753:data<=-16'd4140;
      65754:data<=-16'd4219;
      65755:data<=-16'd3715;
      65756:data<=-16'd3463;
      65757:data<=-16'd3139;
      65758:data<=-16'd998;
      65759:data<=-16'd913;
      65760:data<=16'd863;
      65761:data<=16'd7406;
      65762:data<=16'd9471;
      65763:data<=16'd8049;
      65764:data<=16'd9266;
      65765:data<=16'd10173;
      65766:data<=16'd10219;
      65767:data<=16'd9873;
      65768:data<=16'd9424;
      65769:data<=16'd9784;
      65770:data<=16'd9407;
      65771:data<=16'd10179;
      65772:data<=16'd11344;
      65773:data<=16'd10467;
      65774:data<=16'd10549;
      65775:data<=16'd10078;
      65776:data<=16'd9119;
      65777:data<=16'd10810;
      65778:data<=16'd11056;
      65779:data<=16'd10255;
      65780:data<=16'd10605;
      65781:data<=16'd9533;
      65782:data<=16'd9454;
      65783:data<=16'd10654;
      65784:data<=16'd10933;
      65785:data<=16'd11248;
      65786:data<=16'd10604;
      65787:data<=16'd10002;
      65788:data<=16'd9850;
      65789:data<=16'd9526;
      65790:data<=16'd10951;
      65791:data<=16'd10860;
      65792:data<=16'd10009;
      65793:data<=16'd11074;
      65794:data<=16'd6749;
      65795:data<=16'd804;
      65796:data<=16'd1950;
      65797:data<=16'd3395;
      65798:data<=16'd2593;
      65799:data<=16'd2828;
      65800:data<=16'd2309;
      65801:data<=16'd2352;
      65802:data<=16'd3838;
      65803:data<=16'd4572;
      65804:data<=16'd4176;
      65805:data<=16'd3494;
      65806:data<=16'd3512;
      65807:data<=16'd3562;
      65808:data<=16'd4309;
      65809:data<=16'd5883;
      65810:data<=16'd5353;
      65811:data<=16'd4872;
      65812:data<=16'd5588;
      65813:data<=16'd4582;
      65814:data<=16'd4608;
      65815:data<=16'd6109;
      65816:data<=16'd6021;
      65817:data<=16'd5791;
      65818:data<=16'd5604;
      65819:data<=16'd4954;
      65820:data<=16'd5186;
      65821:data<=16'd6244;
      65822:data<=16'd6693;
      65823:data<=16'd5644;
      65824:data<=16'd5706;
      65825:data<=16'd6024;
      65826:data<=16'd4264;
      65827:data<=16'd7494;
      65828:data<=16'd14645;
      65829:data<=16'd15635;
      65830:data<=16'd14020;
      65831:data<=16'd13934;
      65832:data<=16'd12885;
      65833:data<=16'd13245;
      65834:data<=16'd14192;
      65835:data<=16'd13467;
      65836:data<=16'd12997;
      65837:data<=16'd12257;
      65838:data<=16'd11403;
      65839:data<=16'd11712;
      65840:data<=16'd12369;
      65841:data<=16'd12348;
      65842:data<=16'd10895;
      65843:data<=16'd9803;
      65844:data<=16'd9941;
      65845:data<=16'd9377;
      65846:data<=16'd8789;
      65847:data<=16'd8340;
      65848:data<=16'd7345;
      65849:data<=16'd6845;
      65850:data<=16'd6408;
      65851:data<=16'd5856;
      65852:data<=16'd4713;
      65853:data<=16'd2843;
      65854:data<=16'd2629;
      65855:data<=16'd2678;
      65856:data<=16'd1923;
      65857:data<=16'd2137;
      65858:data<=16'd889;
      65859:data<=-16'd807;
      65860:data<=-16'd872;
      65861:data<=-16'd4648;
      65862:data<=-16'd10266;
      65863:data<=-16'd10781;
      65864:data<=-16'd9970;
      65865:data<=-16'd11523;
      65866:data<=-16'd12026;
      65867:data<=-16'd11309;
      65868:data<=-16'd11256;
      65869:data<=-16'd10875;
      65870:data<=-16'd10775;
      65871:data<=-16'd12051;
      65872:data<=-16'd12540;
      65873:data<=-16'd12185;
      65874:data<=-16'd12228;
      65875:data<=-16'd11370;
      65876:data<=-16'd11041;
      65877:data<=-16'd12396;
      65878:data<=-16'd12739;
      65879:data<=-16'd12072;
      65880:data<=-16'd11637;
      65881:data<=-16'd11333;
      65882:data<=-16'd11368;
      65883:data<=-16'd11362;
      65884:data<=-16'd11935;
      65885:data<=-16'd12484;
      65886:data<=-16'd11884;
      65887:data<=-16'd11837;
      65888:data<=-16'd11274;
      65889:data<=-16'd10722;
      65890:data<=-16'd12765;
      65891:data<=-16'd12716;
      65892:data<=-16'd11318;
      65893:data<=-16'd12712;
      65894:data<=-16'd9527;
      65895:data<=-16'd3037;
      65896:data<=-16'd3022;
      65897:data<=-16'd4760;
      65898:data<=-16'd3691;
      65899:data<=-16'd3644;
      65900:data<=-16'd3726;
      65901:data<=-16'd3363;
      65902:data<=-16'd4413;
      65903:data<=-16'd5413;
      65904:data<=-16'd5298;
      65905:data<=-16'd5137;
      65906:data<=-16'd5074;
      65907:data<=-16'd4349;
      65908:data<=-16'd4366;
      65909:data<=-16'd6090;
      65910:data<=-16'd6655;
      65911:data<=-16'd6028;
      65912:data<=-16'd6193;
      65913:data<=-16'd5694;
      65914:data<=-16'd5535;
      65915:data<=-16'd6902;
      65916:data<=-16'd7021;
      65917:data<=-16'd6329;
      65918:data<=-16'd6241;
      65919:data<=-16'd5770;
      65920:data<=-16'd5839;
      65921:data<=-16'd6810;
      65922:data<=-16'd7095;
      65923:data<=-16'd6388;
      65924:data<=-16'd6065;
      65925:data<=-16'd6581;
      65926:data<=-16'd5855;
      65927:data<=-16'd6040;
      65928:data<=-16'd11217;
      65929:data<=-16'd15938;
      65930:data<=-16'd15641;
      65931:data<=-16'd14505;
      65932:data<=-16'd13816;
      65933:data<=-16'd13549;
      65934:data<=-16'd14701;
      65935:data<=-16'd14518;
      65936:data<=-16'd13251;
      65937:data<=-16'd12988;
      65938:data<=-16'd12275;
      65939:data<=-16'd12087;
      65940:data<=-16'd13133;
      65941:data<=-16'd12747;
      65942:data<=-16'd11452;
      65943:data<=-16'd10956;
      65944:data<=-16'd10484;
      65945:data<=-16'd9829;
      65946:data<=-16'd9227;
      65947:data<=-16'd8338;
      65948:data<=-16'd7642;
      65949:data<=-16'd7423;
      65950:data<=-16'd7003;
      65951:data<=-16'd6519;
      65952:data<=-16'd5495;
      65953:data<=-16'd3475;
      65954:data<=-16'd2790;
      65955:data<=-16'd2807;
      65956:data<=-16'd1791;
      65957:data<=-16'd2159;
      65958:data<=-16'd1436;
      65959:data<=16'd1248;
      65960:data<=16'd558;
      65961:data<=16'd2443;
      65962:data<=16'd9524;
      65963:data<=16'd11013;
      65964:data<=16'd9806;
      65965:data<=16'd12078;
      65966:data<=16'd12289;
      65967:data<=16'd11676;
      65968:data<=16'd12049;
      65969:data<=16'd10944;
      65970:data<=16'd11435;
      65971:data<=16'd13001;
      65972:data<=16'd13098;
      65973:data<=16'd12921;
      65974:data<=16'd12284;
      65975:data<=16'd12096;
      65976:data<=16'd12098;
      65977:data<=16'd11762;
      65978:data<=16'd13007;
      65979:data<=16'd13268;
      65980:data<=16'd12176;
      65981:data<=16'd12386;
      65982:data<=16'd11731;
      65983:data<=16'd11715;
      65984:data<=16'd13635;
      65985:data<=16'd13574;
      65986:data<=16'd12804;
      65987:data<=16'd12634;
      65988:data<=16'd11546;
      65989:data<=16'd11476;
      65990:data<=16'd12963;
      65991:data<=16'd13612;
      65992:data<=16'd12404;
      65993:data<=16'd11747;
      65994:data<=16'd11637;
      65995:data<=16'd7454;
      65996:data<=16'd3418;
      65997:data<=16'd4786;
      65998:data<=16'd5304;
      65999:data<=16'd4363;
      66000:data<=16'd4927;
      66001:data<=16'd3990;
      66002:data<=16'd4193;
      66003:data<=16'd6417;
      66004:data<=16'd6240;
      66005:data<=16'd5858;
      66006:data<=16'd6072;
      66007:data<=16'd5069;
      66008:data<=16'd5562;
      66009:data<=16'd7218;
      66010:data<=16'd7313;
      66011:data<=16'd6849;
      66012:data<=16'd6818;
      66013:data<=16'd6537;
      66014:data<=16'd6583;
      66015:data<=16'd7677;
      66016:data<=16'd7993;
      66017:data<=16'd7203;
      66018:data<=16'd7269;
      66019:data<=16'd7309;
      66020:data<=16'd6663;
      66021:data<=16'd6919;
      66022:data<=16'd8067;
      66023:data<=16'd8399;
      66024:data<=16'd7298;
      66025:data<=16'd7186;
      66026:data<=16'd7515;
      66027:data<=16'd6492;
      66028:data<=16'd9737;
      66029:data<=16'd16167;
      66030:data<=16'd17080;
      66031:data<=16'd15393;
      66032:data<=16'd15038;
      66033:data<=16'd14474;
      66034:data<=16'd15406;
      66035:data<=16'd15688;
      66036:data<=16'd14299;
      66037:data<=16'd14436;
      66038:data<=16'd13846;
      66039:data<=16'd12962;
      66040:data<=16'd13856;
      66041:data<=16'd13623;
      66042:data<=16'd13042;
      66043:data<=16'd12894;
      66044:data<=16'd11618;
      66045:data<=16'd10886;
      66046:data<=16'd10548;
      66047:data<=16'd9744;
      66048:data<=16'd9315;
      66049:data<=16'd8567;
      66050:data<=16'd8025;
      66051:data<=16'd8319;
      66052:data<=16'd7533;
      66053:data<=16'd5257;
      66054:data<=16'd3849;
      66055:data<=16'd3841;
      66056:data<=16'd3407;
      66057:data<=16'd3309;
      66058:data<=16'd3058;
      66059:data<=16'd581;
      66060:data<=-16'd381;
      66061:data<=-16'd472;
      66062:data<=-16'd4896;
      66063:data<=-16'd8833;
      66064:data<=-16'd9191;
      66065:data<=-16'd10067;
      66066:data<=-16'd10718;
      66067:data<=-16'd10360;
      66068:data<=-16'd10255;
      66069:data<=-16'd10111;
      66070:data<=-16'd10246;
      66071:data<=-16'd10520;
      66072:data<=-16'd11239;
      66073:data<=-16'd11850;
      66074:data<=-16'd11207;
      66075:data<=-16'd10784;
      66076:data<=-16'd10276;
      66077:data<=-16'd10266;
      66078:data<=-16'd11955;
      66079:data<=-16'd11917;
      66080:data<=-16'd11035;
      66081:data<=-16'd11259;
      66082:data<=-16'd10379;
      66083:data<=-16'd10645;
      66084:data<=-16'd12070;
      66085:data<=-16'd11900;
      66086:data<=-16'd11659;
      66087:data<=-16'd11176;
      66088:data<=-16'd10969;
      66089:data<=-16'd11250;
      66090:data<=-16'd10769;
      66091:data<=-16'd11853;
      66092:data<=-16'd11817;
      66093:data<=-16'd10361;
      66094:data<=-16'd11785;
      66095:data<=-16'd8799;
      66096:data<=-16'd2458;
      66097:data<=-16'd3028;
      66098:data<=-16'd4375;
      66099:data<=-16'd3313;
      66100:data<=-16'd4076;
      66101:data<=-16'd3519;
      66102:data<=-16'd3573;
      66103:data<=-16'd5375;
      66104:data<=-16'd4940;
      66105:data<=-16'd4676;
      66106:data<=-16'd4980;
      66107:data<=-16'd4548;
      66108:data<=-16'd5177;
      66109:data<=-16'd5885;
      66110:data<=-16'd6285;
      66111:data<=-16'd6401;
      66112:data<=-16'd6132;
      66113:data<=-16'd6357;
      66114:data<=-16'd5673;
      66115:data<=-16'd5865;
      66116:data<=-16'd7679;
      66117:data<=-16'd7037;
      66118:data<=-16'd6179;
      66119:data<=-16'd6763;
      66120:data<=-16'd6035;
      66121:data<=-16'd6398;
      66122:data<=-16'd7884;
      66123:data<=-16'd7418;
      66124:data<=-16'd6713;
      66125:data<=-16'd7048;
      66126:data<=-16'd7039;
      66127:data<=-16'd6516;
      66128:data<=-16'd8276;
      66129:data<=-16'd12932;
      66130:data<=-16'd15720;
      66131:data<=-16'd15547;
      66132:data<=-16'd14610;
      66133:data<=-16'd13576;
      66134:data<=-16'd14352;
      66135:data<=-16'd15323;
      66136:data<=-16'd14286;
      66137:data<=-16'd13870;
      66138:data<=-16'd13364;
      66139:data<=-16'd12073;
      66140:data<=-16'd12616;
      66141:data<=-16'd13432;
      66142:data<=-16'd12813;
      66143:data<=-16'd11855;
      66144:data<=-16'd11148;
      66145:data<=-16'd10968;
      66146:data<=-16'd10457;
      66147:data<=-16'd9614;
      66148:data<=-16'd9174;
      66149:data<=-16'd8520;
      66150:data<=-16'd8126;
      66151:data<=-16'd7982;
      66152:data<=-16'd6943;
      66153:data<=-16'd5101;
      66154:data<=-16'd3636;
      66155:data<=-16'd3905;
      66156:data<=-16'd3967;
      66157:data<=-16'd2826;
      66158:data<=-16'd2801;
      66159:data<=-16'd1330;
      66160:data<=16'd813;
      66161:data<=-16'd563;
      66162:data<=16'd1676;
      66163:data<=16'd8486;
      66164:data<=16'd9832;
      66165:data<=16'd8895;
      66166:data<=16'd10662;
      66167:data<=16'd10702;
      66168:data<=16'd10043;
      66169:data<=16'd10188;
      66170:data<=16'd9445;
      66171:data<=16'd10126;
      66172:data<=16'd11771;
      66173:data<=16'd11650;
      66174:data<=16'd11060;
      66175:data<=16'd10569;
      66176:data<=16'd10026;
      66177:data<=16'd10669;
      66178:data<=16'd11652;
      66179:data<=16'd11576;
      66180:data<=16'd11119;
      66181:data<=16'd10857;
      66182:data<=16'd10560;
      66183:data<=16'd10372;
      66184:data<=16'd10909;
      66185:data<=16'd11826;
      66186:data<=16'd11644;
      66187:data<=16'd10945;
      66188:data<=16'd10775;
      66189:data<=16'd9862;
      66190:data<=16'd9858;
      66191:data<=16'd11958;
      66192:data<=16'd11670;
      66193:data<=16'd10149;
      66194:data<=16'd11051;
      66195:data<=16'd9194;
      66196:data<=16'd4322;
      66197:data<=16'd2784;
      66198:data<=16'd3136;
      66199:data<=16'd3051;
      66200:data<=16'd3512;
      66201:data<=16'd3304;
      66202:data<=16'd3054;
      66203:data<=16'd4056;
      66204:data<=16'd4851;
      66205:data<=16'd4763;
      66206:data<=16'd4505;
      66207:data<=16'd4441;
      66208:data<=16'd4094;
      66209:data<=16'd4328;
      66210:data<=16'd5843;
      66211:data<=16'd6014;
      66212:data<=16'd5288;
      66213:data<=16'd5583;
      66214:data<=16'd4911;
      66215:data<=16'd5004;
      66216:data<=16'd6830;
      66217:data<=16'd6376;
      66218:data<=16'd5488;
      66219:data<=16'd5894;
      66220:data<=16'd5374;
      66221:data<=16'd5808;
      66222:data<=16'd6683;
      66223:data<=16'd6184;
      66224:data<=16'd6252;
      66225:data<=16'd6100;
      66226:data<=16'd5827;
      66227:data<=16'd6015;
      66228:data<=16'd5315;
      66229:data<=16'd8097;
      66230:data<=16'd14193;
      66231:data<=16'd15664;
      66232:data<=16'd13640;
      66233:data<=16'd12831;
      66234:data<=16'd12960;
      66235:data<=16'd13731;
      66236:data<=16'd13486;
      66237:data<=16'd12286;
      66238:data<=16'd12213;
      66239:data<=16'd11799;
      66240:data<=16'd11311;
      66241:data<=16'd11987;
      66242:data<=16'd11779;
      66243:data<=16'd10895;
      66244:data<=16'd10578;
      66245:data<=16'd10131;
      66246:data<=16'd9494;
      66247:data<=16'd8634;
      66248:data<=16'd7859;
      66249:data<=16'd7652;
      66250:data<=16'd7306;
      66251:data<=16'd6821;
      66252:data<=16'd6261;
      66253:data<=16'd4786;
      66254:data<=16'd3213;
      66255:data<=16'd2952;
      66256:data<=16'd2801;
      66257:data<=16'd2061;
      66258:data<=16'd2237;
      66259:data<=16'd1451;
      66260:data<=-16'd1010;
      66261:data<=-16'd887;
      66262:data<=-16'd1466;
      66263:data<=-16'd6898;
      66264:data<=-16'd10202;
      66265:data<=-16'd10216;
      66266:data<=-16'd11517;
      66267:data<=-16'd11562;
      66268:data<=-16'd10897;
      66269:data<=-16'd11335;
      66270:data<=-16'd10615;
      66271:data<=-16'd10772;
      66272:data<=-16'd12135;
      66273:data<=-16'd12102;
      66274:data<=-16'd11966;
      66275:data<=-16'd11687;
      66276:data<=-16'd11057;
      66277:data<=-16'd11268;
      66278:data<=-16'd11623;
      66279:data<=-16'd12126;
      66280:data<=-16'd12234;
      66281:data<=-16'd11737;
      66282:data<=-16'd11591;
      66283:data<=-16'd11139;
      66284:data<=-16'd11928;
      66285:data<=-16'd13643;
      66286:data<=-16'd12889;
      66287:data<=-16'd11896;
      66288:data<=-16'd11858;
      66289:data<=-16'd11297;
      66290:data<=-16'd11941;
      66291:data<=-16'd12819;
      66292:data<=-16'd12665;
      66293:data<=-16'd12213;
      66294:data<=-16'd11706;
      66295:data<=-16'd12276;
      66296:data<=-16'd9929;
      66297:data<=-16'd4226;
      66298:data<=-16'd3524;
      66299:data<=-16'd5259;
      66300:data<=-16'd4273;
      66301:data<=-16'd4408;
      66302:data<=-16'd4353;
      66303:data<=-16'd4152;
      66304:data<=-16'd6175;
      66305:data<=-16'd5987;
      66306:data<=-16'd5089;
      66307:data<=-16'd6216;
      66308:data<=-16'd5711;
      66309:data<=-16'd5758;
      66310:data<=-16'd7432;
      66311:data<=-16'd6946;
      66312:data<=-16'd6384;
      66313:data<=-16'd6943;
      66314:data<=-16'd6399;
      66315:data<=-16'd6354;
      66316:data<=-16'd7538;
      66317:data<=-16'd7752;
      66318:data<=-16'd7245;
      66319:data<=-16'd7036;
      66320:data<=-16'd6372;
      66321:data<=-16'd6166;
      66322:data<=-16'd7347;
      66323:data<=-16'd7909;
      66324:data<=-16'd7371;
      66325:data<=-16'd6942;
      66326:data<=-16'd6757;
      66327:data<=-16'd6549;
      66328:data<=-16'd6208;
      66329:data<=-16'd8483;
      66330:data<=-16'd13778;
      66331:data<=-16'd16327;
      66332:data<=-16'd15549;
      66333:data<=-16'd14791;
      66334:data<=-16'd14189;
      66335:data<=-16'd14791;
      66336:data<=-16'd15224;
      66337:data<=-16'd14026;
      66338:data<=-16'd13715;
      66339:data<=-16'd12954;
      66340:data<=-16'd11822;
      66341:data<=-16'd12834;
      66342:data<=-16'd12909;
      66343:data<=-16'd11794;
      66344:data<=-16'd11511;
      66345:data<=-16'd10610;
      66346:data<=-16'd10085;
      66347:data<=-16'd10097;
      66348:data<=-16'd9374;
      66349:data<=-16'd8837;
      66350:data<=-16'd8055;
      66351:data<=-16'd7500;
      66352:data<=-16'd7603;
      66353:data<=-16'd6455;
      66354:data<=-16'd4602;
      66355:data<=-16'd3530;
      66356:data<=-16'd3395;
      66357:data<=-16'd3175;
      66358:data<=-16'd2261;
      66359:data<=-16'd1833;
      66360:data<=-16'd335;
      66361:data<=16'd1093;
      66362:data<=-16'd315;
      66363:data<=16'd2437;
      66364:data<=16'd9458;
      66365:data<=16'd10998;
      66366:data<=16'd10285;
      66367:data<=16'd11674;
      66368:data<=16'd11297;
      66369:data<=16'd10892;
      66370:data<=16'd11227;
      66371:data<=16'd10360;
      66372:data<=16'd11021;
      66373:data<=16'd12557;
      66374:data<=16'd12082;
      66375:data<=16'd11474;
      66376:data<=16'd11483;
      66377:data<=16'd10748;
      66378:data<=16'd11082;
      66379:data<=16'd12889;
      66380:data<=16'd12910;
      66381:data<=16'd12169;
      66382:data<=16'd12452;
      66383:data<=16'd11746;
      66384:data<=16'd11909;
      66385:data<=16'd13602;
      66386:data<=16'd13399;
      66387:data<=16'd12900;
      66388:data<=16'd12986;
      66389:data<=16'd12161;
      66390:data<=16'd12178;
      66391:data<=16'd13097;
      66392:data<=16'd13808;
      66393:data<=16'd13315;
      66394:data<=16'd12231;
      66395:data<=16'd13097;
      66396:data<=16'd11304;
      66397:data<=16'd5833;
      66398:data<=16'd4517;
      66399:data<=16'd5257;
      66400:data<=16'd4760;
      66401:data<=16'd5521;
      66402:data<=16'd4863;
      66403:data<=16'd4648;
      66404:data<=16'd6968;
      66405:data<=16'd6875;
      66406:data<=16'd6443;
      66407:data<=16'd7222;
      66408:data<=16'd6302;
      66409:data<=16'd6637;
      66410:data<=16'd8156;
      66411:data<=16'd8122;
      66412:data<=16'd8026;
      66413:data<=16'd7865;
      66414:data<=16'd7285;
      66415:data<=16'd7286;
      66416:data<=16'd8207;
      66417:data<=16'd8918;
      66418:data<=16'd8067;
      66419:data<=16'd7755;
      66420:data<=16'd7846;
      66421:data<=16'd6716;
      66422:data<=16'd7500;
      66423:data<=16'd8912;
      66424:data<=16'd8378;
      66425:data<=16'd8404;
      66426:data<=16'd7826;
      66427:data<=16'd7124;
      66428:data<=16'd8059;
      66429:data<=16'd7821;
      66430:data<=16'd10157;
      66431:data<=16'd16220;
      66432:data<=16'd17371;
      66433:data<=16'd14938;
      66434:data<=16'd15250;
      66435:data<=16'd16178;
      66436:data<=16'd15802;
      66437:data<=16'd14924;
      66438:data<=16'd14110;
      66439:data<=16'd13665;
      66440:data<=16'd13223;
      66441:data<=16'd13414;
      66442:data<=16'd13773;
      66443:data<=16'd12859;
      66444:data<=16'd11734;
      66445:data<=16'd11326;
      66446:data<=16'd11095;
      66447:data<=16'd10712;
      66448:data<=16'd10073;
      66449:data<=16'd9427;
      66450:data<=16'd8931;
      66451:data<=16'd8687;
      66452:data<=16'd8370;
      66453:data<=16'd7145;
      66454:data<=16'd5483;
      66455:data<=16'd4402;
      66456:data<=16'd4035;
      66457:data<=16'd3880;
      66458:data<=16'd3595;
      66459:data<=16'd3145;
      66460:data<=16'd1516;
      66461:data<=16'd118;
      66462:data<=16'd1048;
      66463:data<=-16'd685;
      66464:data<=-16'd6564;
      66465:data<=-16'd9423;
      66466:data<=-16'd9659;
      66467:data<=-16'd10866;
      66468:data<=-16'd10407;
      66469:data<=-16'd9502;
      66470:data<=-16'd10053;
      66471:data<=-16'd9788;
      66472:data<=-16'd9953;
      66473:data<=-16'd11036;
      66474:data<=-16'd10809;
      66475:data<=-16'd10508;
      66476:data<=-16'd10552;
      66477:data<=-16'd9828;
      66478:data<=-16'd9835;
      66479:data<=-16'd10725;
      66480:data<=-16'd10875;
      66481:data<=-16'd10853;
      66482:data<=-16'd11035;
      66483:data<=-16'd10282;
      66484:data<=-16'd9797;
      66485:data<=-16'd10986;
      66486:data<=-16'd11643;
      66487:data<=-16'd11168;
      66488:data<=-16'd11180;
      66489:data<=-16'd10658;
      66490:data<=-16'd9835;
      66491:data<=-16'd10477;
      66492:data<=-16'd11449;
      66493:data<=-16'd11681;
      66494:data<=-16'd11148;
      66495:data<=-16'd10598;
      66496:data<=-16'd10848;
      66497:data<=-16'd8780;
      66498:data<=-16'd4184;
      66499:data<=-16'd2619;
      66500:data<=-16'd3601;
      66501:data<=-16'd3174;
      66502:data<=-16'd2523;
      66503:data<=-16'd3130;
      66504:data<=-16'd4341;
      66505:data<=-16'd5049;
      66506:data<=-16'd4786;
      66507:data<=-16'd4749;
      66508:data<=-16'd4755;
      66509:data<=-16'd4455;
      66510:data<=-16'd5510;
      66511:data<=-16'd6830;
      66512:data<=-16'd6398;
      66513:data<=-16'd5976;
      66514:data<=-16'd6128;
      66515:data<=-16'd5344;
      66516:data<=-16'd5353;
      66517:data<=-16'd6827;
      66518:data<=-16'd6837;
      66519:data<=-16'd6297;
      66520:data<=-16'd6596;
      66521:data<=-16'd5759;
      66522:data<=-16'd5959;
      66523:data<=-16'd7806;
      66524:data<=-16'd7582;
      66525:data<=-16'd7163;
      66526:data<=-16'd7183;
      66527:data<=-16'd5888;
      66528:data<=-16'd6243;
      66529:data<=-16'd7074;
      66530:data<=-16'd8044;
      66531:data<=-16'd12863;
      66532:data<=-16'd16089;
      66533:data<=-16'd14759;
      66534:data<=-16'd14357;
      66535:data<=-16'd14745;
      66536:data<=-16'd14747;
      66537:data<=-16'd14642;
      66538:data<=-16'd13584;
      66539:data<=-16'd13106;
      66540:data<=-16'd12601;
      66541:data<=-16'd12058;
      66542:data<=-16'd13092;
      66543:data<=-16'd12859;
      66544:data<=-16'd11608;
      66545:data<=-16'd11470;
      66546:data<=-16'd10696;
      66547:data<=-16'd9946;
      66548:data<=-16'd9831;
      66549:data<=-16'd9280;
      66550:data<=-16'd8522;
      66551:data<=-16'd7847;
      66552:data<=-16'd8134;
      66553:data<=-16'd7450;
      66554:data<=-16'd5024;
      66555:data<=-16'd4373;
      66556:data<=-16'd3941;
      66557:data<=-16'd2963;
      66558:data<=-16'd3494;
      66559:data<=-16'd2908;
      66560:data<=-16'd1651;
      66561:data<=-16'd453;
      66562:data<=16'd676;
      66563:data<=-16'd928;
      66564:data<=16'd1318;
      66565:data<=16'd8523;
      66566:data<=16'd10340;
      66567:data<=16'd10031;
      66568:data<=16'd11462;
      66569:data<=16'd10470;
      66570:data<=16'd10131;
      66571:data<=16'd10232;
      66572:data<=16'd9527;
      66573:data<=16'd11041;
      66574:data<=16'd11492;
      66575:data<=16'd10784;
      66576:data<=16'd11032;
      66577:data<=16'd9928;
      66578:data<=16'd9770;
      66579:data<=16'd11041;
      66580:data<=16'd11277;
      66581:data<=16'd11307;
      66582:data<=16'd10713;
      66583:data<=16'd10267;
      66584:data<=16'd10113;
      66585:data<=16'd9641;
      66586:data<=16'd10957;
      66587:data<=16'd11518;
      66588:data<=16'd10662;
      66589:data<=16'd10837;
      66590:data<=16'd9565;
      66591:data<=16'd9389;
      66592:data<=16'd11467;
      66593:data<=16'd11197;
      66594:data<=16'd11116;
      66595:data<=16'd10945;
      66596:data<=16'd9517;
      66597:data<=16'd10631;
      66598:data<=16'd8851;
      66599:data<=16'd3404;
      66600:data<=16'd2232;
      66601:data<=16'd2726;
      66602:data<=16'd2352;
      66603:data<=16'd3033;
      66604:data<=16'd3704;
      66605:data<=16'd4595;
      66606:data<=16'd4372;
      66607:data<=16'd3706;
      66608:data<=16'd4629;
      66609:data<=16'd3830;
      66610:data<=16'd3430;
      66611:data<=16'd5550;
      66612:data<=16'd5368;
      66613:data<=16'd4966;
      66614:data<=16'd5887;
      66615:data<=16'd4614;
      66616:data<=16'd4426;
      66617:data<=16'd6449;
      66618:data<=16'd6643;
      66619:data<=16'd5996;
      66620:data<=16'd5962;
      66621:data<=16'd5250;
      66622:data<=16'd4922;
      66623:data<=16'd6334;
      66624:data<=16'd7043;
      66625:data<=16'd6223;
      66626:data<=16'd6299;
      66627:data<=16'd6002;
      66628:data<=16'd5215;
      66629:data<=16'd6129;
      66630:data<=16'd6105;
      66631:data<=16'd7298;
      66632:data<=16'd12995;
      66633:data<=16'd15359;
      66634:data<=16'd13089;
      66635:data<=16'd13399;
      66636:data<=16'd14378;
      66637:data<=16'd13514;
      66638:data<=16'd13066;
      66639:data<=16'd12352;
      66640:data<=16'd11314;
      66641:data<=16'd11606;
      66642:data<=16'd12592;
      66643:data<=16'd12555;
      66644:data<=16'd11539;
      66645:data<=16'd10857;
      66646:data<=16'd10399;
      66647:data<=16'd9897;
      66648:data<=16'd9345;
      66649:data<=16'd8320;
      66650:data<=16'd7859;
      66651:data<=16'd7697;
      66652:data<=16'd7063;
      66653:data<=16'd6781;
      66654:data<=16'd5224;
      66655:data<=16'd3081;
      66656:data<=16'd3121;
      66657:data<=16'd2936;
      66658:data<=16'd2297;
      66659:data<=16'd2397;
      66660:data<=16'd1105;
      66661:data<=16'd123;
      66662:data<=-16'd299;
      66663:data<=-16'd1356;
      66664:data<=-16'd362;
      66665:data<=-16'd2076;
      66666:data<=-16'd9186;
      66667:data<=-16'd12519;
      66668:data<=-16'd11580;
      66669:data<=-16'd11770;
      66670:data<=-16'd11311;
      66671:data<=-16'd10596;
      66672:data<=-16'd11104;
      66673:data<=-16'd11794;
      66674:data<=-16'd12604;
      66675:data<=-16'd12367;
      66676:data<=-16'd11781;
      66677:data<=-16'd11834;
      66678:data<=-16'd11051;
      66679:data<=-16'd11482;
      66680:data<=-16'd13018;
      66681:data<=-16'd12337;
      66682:data<=-16'd12017;
      66683:data<=-16'd12504;
      66684:data<=-16'd10944;
      66685:data<=-16'd10690;
      66686:data<=-16'd12558;
      66687:data<=-16'd12471;
      66688:data<=-16'd11731;
      66689:data<=-16'd11884;
      66690:data<=-16'd11060;
      66691:data<=-16'd11009;
      66692:data<=-16'd12554;
      66693:data<=-16'd12398;
      66694:data<=-16'd11706;
      66695:data<=-16'd12188;
      66696:data<=-16'd11139;
      66697:data<=-16'd10727;
      66698:data<=-16'd12254;
      66699:data<=-16'd9317;
      66700:data<=-16'd3773;
      66701:data<=-16'd3174;
      66702:data<=-16'd4211;
      66703:data<=-16'd3146;
      66704:data<=-16'd3568;
      66705:data<=-16'd5242;
      66706:data<=-16'd5375;
      66707:data<=-16'd5154;
      66708:data<=-16'd5053;
      66709:data<=-16'd4222;
      66710:data<=-16'd4611;
      66711:data<=-16'd6188;
      66712:data<=-16'd6041;
      66713:data<=-16'd5512;
      66714:data<=-16'd5974;
      66715:data<=-16'd5447;
      66716:data<=-16'd5278;
      66717:data<=-16'd6601;
      66718:data<=-16'd7060;
      66719:data<=-16'd6663;
      66720:data<=-16'd6639;
      66721:data<=-16'd6792;
      66722:data<=-16'd6643;
      66723:data<=-16'd6649;
      66724:data<=-16'd7471;
      66725:data<=-16'd7418;
      66726:data<=-16'd6948;
      66727:data<=-16'd7421;
      66728:data<=-16'd6294;
      66729:data<=-16'd6222;
      66730:data<=-16'd8643;
      66731:data<=-16'd7594;
      66732:data<=-16'd8100;
      66733:data<=-16'd14301;
      66734:data<=-16'd16239;
      66735:data<=-16'd14860;
      66736:data<=-16'd16308;
      66737:data<=-16'd16063;
      66738:data<=-16'd14678;
      66739:data<=-16'd14818;
      66740:data<=-16'd14020;
      66741:data<=-16'd13546;
      66742:data<=-16'd14166;
      66743:data<=-16'd14216;
      66744:data<=-16'd13843;
      66745:data<=-16'd13148;
      66746:data<=-16'd12619;
      66747:data<=-16'd12066;
      66748:data<=-16'd11156;
      66749:data<=-16'd10969;
      66750:data<=-16'd10589;
      66751:data<=-16'd9198;
      66752:data<=-16'd8334;
      66753:data<=-16'd8375;
      66754:data<=-16'd7521;
      66755:data<=-16'd5200;
      66756:data<=-16'd4347;
      66757:data<=-16'd4845;
      66758:data<=-16'd4064;
      66759:data<=-16'd4065;
      66760:data<=-16'd3588;
      66761:data<=-16'd787;
      66762:data<=-16'd438;
      66763:data<=-16'd711;
      66764:data<=16'd400;
      66765:data<=-16'd984;
      66766:data<=16'd1583;
      66767:data<=16'd9785;
      66768:data<=16'd12248;
      66769:data<=16'd10214;
      66770:data<=16'd10648;
      66771:data<=16'd10807;
      66772:data<=16'd9956;
      66773:data<=16'd10549;
      66774:data<=16'd11676;
      66775:data<=16'd11735;
      66776:data<=16'd11500;
      66777:data<=16'd11641;
      66778:data<=16'd10709;
      66779:data<=16'd10631;
      66780:data<=16'd12842;
      66781:data<=16'd12912;
      66782:data<=16'd11418;
      66783:data<=16'd11473;
      66784:data<=16'd10894;
      66785:data<=16'd10754;
      66786:data<=16'd12343;
      66787:data<=16'd12398;
      66788:data<=16'd11318;
      66789:data<=16'd11101;
      66790:data<=16'd10986;
      66791:data<=16'd10790;
      66792:data<=16'd11464;
      66793:data<=16'd12384;
      66794:data<=16'd11788;
      66795:data<=16'd11253;
      66796:data<=16'd11265;
      66797:data<=16'd9641;
      66798:data<=16'd10351;
      66799:data<=16'd12601;
      66800:data<=16'd8193;
      66801:data<=16'd2526;
      66802:data<=16'd2544;
      66803:data<=16'd2704;
      66804:data<=16'd2857;
      66805:data<=16'd4810;
      66806:data<=16'd4658;
      66807:data<=16'd3993;
      66808:data<=16'd4460;
      66809:data<=16'd3842;
      66810:data<=16'd3874;
      66811:data<=16'd5351;
      66812:data<=16'd5612;
      66813:data<=16'd4752;
      66814:data<=16'd4758;
      66815:data<=16'd5174;
      66816:data<=16'd4874;
      66817:data<=16'd5286;
      66818:data<=16'd6532;
      66819:data<=16'd6754;
      66820:data<=16'd6557;
      66821:data<=16'd6305;
      66822:data<=16'd5759;
      66823:data<=16'd6297;
      66824:data<=16'd7424;
      66825:data<=16'd7609;
      66826:data<=16'd6910;
      66827:data<=16'd6261;
      66828:data<=16'd6320;
      66829:data<=16'd6545;
      66830:data<=16'd7547;
      66831:data<=16'd8301;
      66832:data<=16'd6717;
      66833:data<=16'd8155;
      66834:data<=16'd13972;
      66835:data<=16'd16023;
      66836:data<=16'd15262;
      66837:data<=16'd16084;
      66838:data<=16'd15617;
      66839:data<=16'd14571;
      66840:data<=16'd14445;
      66841:data<=16'd13775;
      66842:data<=16'd13878;
      66843:data<=16'd14606;
      66844:data<=16'd14402;
      66845:data<=16'd13576;
      66846:data<=16'd12666;
      66847:data<=16'd12442;
      66848:data<=16'd11916;
      66849:data<=16'd10790;
      66850:data<=16'd10566;
      66851:data<=16'd9855;
      66852:data<=16'd8748;
      66853:data<=16'd8830;
      66854:data<=16'd8067;
      66855:data<=16'd5959;
      66856:data<=16'd4655;
      66857:data<=16'd4989;
      66858:data<=16'd5406;
      66859:data<=16'd4394;
      66860:data<=16'd3742;
      66861:data<=16'd2902;
      66862:data<=16'd1027;
      66863:data<=16'd1400;
      66864:data<=16'd1327;
      66865:data<=-16'd115;
      66866:data<=16'd1428;
      66867:data<=-16'd1348;
      66868:data<=-16'd9784;
      66869:data<=-16'd11702;
      66870:data<=-16'd9805;
      66871:data<=-16'd10396;
      66872:data<=-16'd9415;
      66873:data<=-16'd9359;
      66874:data<=-16'd11670;
      66875:data<=-16'd11583;
      66876:data<=-16'd10880;
      66877:data<=-16'd11030;
      66878:data<=-16'd10228;
      66879:data<=-16'd10342;
      66880:data<=-16'd11690;
      66881:data<=-16'd11790;
      66882:data<=-16'd10919;
      66883:data<=-16'd10561;
      66884:data<=-16'd10317;
      66885:data<=-16'd10157;
      66886:data<=-16'd11056;
      66887:data<=-16'd11747;
      66888:data<=-16'd11142;
      66889:data<=-16'd10701;
      66890:data<=-16'd10414;
      66891:data<=-16'd9740;
      66892:data<=-16'd10087;
      66893:data<=-16'd11383;
      66894:data<=-16'd11546;
      66895:data<=-16'd10481;
      66896:data<=-16'd9868;
      66897:data<=-16'd9523;
      66898:data<=-16'd9790;
      66899:data<=-16'd11711;
      66900:data<=-16'd10909;
      66901:data<=-16'd5272;
      66902:data<=-16'd1278;
      66903:data<=-16'd1054;
      66904:data<=-16'd1491;
      66905:data<=-16'd2631;
      66906:data<=-16'd3435;
      66907:data<=-16'd2681;
      66908:data<=-16'd2305;
      66909:data<=-16'd2485;
      66910:data<=-16'd2347;
      66911:data<=-16'd2910;
      66912:data<=-16'd4105;
      66913:data<=-16'd4235;
      66914:data<=-16'd3762;
      66915:data<=-16'd3935;
      66916:data<=-16'd3563;
      66917:data<=-16'd3519;
      66918:data<=-16'd5140;
      66919:data<=-16'd5363;
      66920:data<=-16'd4360;
      66921:data<=-16'd4369;
      66922:data<=-16'd3996;
      66923:data<=-16'd4432;
      66924:data<=-16'd5773;
      66925:data<=-16'd5509;
      66926:data<=-16'd5406;
      66927:data<=-16'd5207;
      66928:data<=-16'd4226;
      66929:data<=-16'd4949;
      66930:data<=-16'd5521;
      66931:data<=-16'd5779;
      66932:data<=-16'd6657;
      66933:data<=-16'd5332;
      66934:data<=-16'd6473;
      66935:data<=-16'd12313;
      66936:data<=-16'd14979;
      66937:data<=-16'd14889;
      66938:data<=-16'd15308;
      66939:data<=-16'd14048;
      66940:data<=-16'd13133;
      66941:data<=-16'd13392;
      66942:data<=-16'd13042;
      66943:data<=-16'd13364;
      66944:data<=-16'd13581;
      66945:data<=-16'd12827;
      66946:data<=-16'd12263;
      66947:data<=-16'd11580;
      66948:data<=-16'd10783;
      66949:data<=-16'd9973;
      66950:data<=-16'd9421;
      66951:data<=-16'd9485;
      66952:data<=-16'd8924;
      66953:data<=-16'd8091;
      66954:data<=-16'd7386;
      66955:data<=-16'd5879;
      66956:data<=-16'd4743;
      66957:data<=-16'd4264;
      66958:data<=-16'd3732;
      66959:data<=-16'd3588;
      66960:data<=-16'd3236;
      66961:data<=-16'd2306;
      66962:data<=-16'd746;
      66963:data<=16'd435;
      66964:data<=-16'd24;
      66965:data<=16'd467;
      66966:data<=16'd1113;
      66967:data<=16'd326;
      66968:data<=16'd4441;
      66969:data<=16'd11573;
      66970:data<=16'd12828;
      66971:data<=16'd11439;
      66972:data<=16'd11515;
      66973:data<=16'd11455;
      66974:data<=16'd12440;
      66975:data<=16'd13164;
      66976:data<=16'd12201;
      66977:data<=16'd12148;
      66978:data<=16'd12348;
      66979:data<=16'd11817;
      66980:data<=16'd12369;
      66981:data<=16'd13229;
      66982:data<=16'd12812;
      66983:data<=16'd12331;
      66984:data<=16'd12176;
      66985:data<=16'd11257;
      66986:data<=16'd11561;
      66987:data<=16'd13611;
      66988:data<=16'd13497;
      66989:data<=16'd12134;
      66990:data<=16'd12052;
      66991:data<=16'd11433;
      66992:data<=16'd11421;
      66993:data<=16'd12595;
      66994:data<=16'd12437;
      66995:data<=16'd11961;
      66996:data<=16'd11559;
      66997:data<=16'd10977;
      66998:data<=16'd11439;
      66999:data<=16'd11923;
      67000:data<=16'd12469;
      67001:data<=16'd11403;
      67002:data<=16'd6068;
      67003:data<=16'd1723;
      67004:data<=16'd1609;
      67005:data<=16'd2607;
      67006:data<=16'd3950;
      67007:data<=16'd4223;
      67008:data<=16'd3272;
      67009:data<=16'd3338;
      67010:data<=16'd3216;
      67011:data<=16'd3409;
      67012:data<=16'd4781;
      67013:data<=16'd4784;
      67014:data<=16'd4208;
      67015:data<=16'd4367;
      67016:data<=16'd4114;
      67017:data<=16'd4173;
      67018:data<=16'd4911;
      67019:data<=16'd5260;
      67020:data<=16'd5145;
      67021:data<=16'd5053;
      67022:data<=16'd4619;
      67023:data<=16'd4118;
      67024:data<=16'd5251;
      67025:data<=16'd6320;
      67026:data<=16'd5714;
      67027:data<=16'd5883;
      67028:data<=16'd5541;
      67029:data<=16'd4373;
      67030:data<=16'd5553;
      67031:data<=16'd6263;
      67032:data<=16'd5897;
      67033:data<=16'd6393;
      67034:data<=16'd5209;
      67035:data<=16'd6714;
      67036:data<=16'd13295;
      67037:data<=16'd16093;
      67038:data<=16'd14566;
      67039:data<=16'd14186;
      67040:data<=16'd13875;
      67041:data<=16'd12982;
      67042:data<=16'd12695;
      67043:data<=16'd13139;
      67044:data<=16'd13420;
      67045:data<=16'd12885;
      67046:data<=16'd12519;
      67047:data<=16'd11664;
      67048:data<=16'd10452;
      67049:data<=16'd10149;
      67050:data<=16'd9303;
      67051:data<=16'd8766;
      67052:data<=16'd8798;
      67053:data<=16'd7662;
      67054:data<=16'd7547;
      67055:data<=16'd6953;
      67056:data<=16'd4253;
      67057:data<=16'd3735;
      67058:data<=16'd3879;
      67059:data<=16'd2914;
      67060:data<=16'd3054;
      67061:data<=16'd1941;
      67062:data<=16'd167;
      67063:data<=-16'd203;
      67064:data<=-16'd760;
      67065:data<=-16'd563;
      67066:data<=-16'd963;
      67067:data<=-16'd2221;
      67068:data<=-16'd1882;
      67069:data<=-16'd5189;
      67070:data<=-16'd11685;
      67071:data<=-16'd13127;
      67072:data<=-16'd11905;
      67073:data<=-16'd12138;
      67074:data<=-16'd12642;
      67075:data<=-16'd13382;
      67076:data<=-16'd13094;
      67077:data<=-16'd12455;
      67078:data<=-16'd12842;
      67079:data<=-16'd12370;
      67080:data<=-16'd12551;
      67081:data<=-16'd13985;
      67082:data<=-16'd13496;
      67083:data<=-16'd12480;
      67084:data<=-16'd12716;
      67085:data<=-16'd12580;
      67086:data<=-16'd12566;
      67087:data<=-16'd13358;
      67088:data<=-16'd13377;
      67089:data<=-16'd12703;
      67090:data<=-16'd12599;
      67091:data<=-16'd12289;
      67092:data<=-16'd11897;
      67093:data<=-16'd12639;
      67094:data<=-16'd12856;
      67095:data<=-16'd12420;
      67096:data<=-16'd12680;
      67097:data<=-16'd11768;
      67098:data<=-16'd10865;
      67099:data<=-16'd12226;
      67100:data<=-16'd13142;
      67101:data<=-16'd12874;
      67102:data<=-16'd10930;
      67103:data<=-16'd5560;
      67104:data<=-16'd1771;
      67105:data<=-16'd3031;
      67106:data<=-16'd4605;
      67107:data<=-16'd4262;
      67108:data<=-16'd4068;
      67109:data<=-16'd4232;
      67110:data<=-16'd3889;
      67111:data<=-16'd3950;
      67112:data<=-16'd4965;
      67113:data<=-16'd5330;
      67114:data<=-16'd5209;
      67115:data<=-16'd5342;
      67116:data<=-16'd4610;
      67117:data<=-16'd4337;
      67118:data<=-16'd5383;
      67119:data<=-16'd5626;
      67120:data<=-16'd5400;
      67121:data<=-16'd5612;
      67122:data<=-16'd5404;
      67123:data<=-16'd4919;
      67124:data<=-16'd5212;
      67125:data<=-16'd6344;
      67126:data<=-16'd6375;
      67127:data<=-16'd5703;
      67128:data<=-16'd6158;
      67129:data<=-16'd5506;
      67130:data<=-16'd5083;
      67131:data<=-16'd7107;
      67132:data<=-16'd6930;
      67133:data<=-16'd6125;
      67134:data<=-16'd7142;
      67135:data<=-16'd5325;
      67136:data<=-16'd6639;
      67137:data<=-16'd14415;
      67138:data<=-16'd16944;
      67139:data<=-16'd14630;
      67140:data<=-16'd14613;
      67141:data<=-16'd13483;
      67142:data<=-16'd12251;
      67143:data<=-16'd13605;
      67144:data<=-16'd13994;
      67145:data<=-16'd13538;
      67146:data<=-16'd13171;
      67147:data<=-16'd12055;
      67148:data<=-16'd11449;
      67149:data<=-16'd10774;
      67150:data<=-16'd9312;
      67151:data<=-16'd8337;
      67152:data<=-16'd7464;
      67153:data<=-16'd6572;
      67154:data<=-16'd6203;
      67155:data<=-16'd5295;
      67156:data<=-16'd3805;
      67157:data<=-16'd3055;
      67158:data<=-16'd2737;
      67159:data<=-16'd2232;
      67160:data<=-16'd2155;
      67161:data<=-16'd1656;
      67162:data<=-16'd2;
      67163:data<=16'd860;
      67164:data<=16'd987;
      67165:data<=16'd1507;
      67166:data<=16'd1271;
      67167:data<=16'd1513;
      67168:data<=16'd2857;
      67169:data<=16'd3322;
      67170:data<=16'd5574;
      67171:data<=16'd10035;
      67172:data<=16'd11028;
      67173:data<=16'd9674;
      67174:data<=16'd10542;
      67175:data<=16'd11564;
      67176:data<=16'd10934;
      67177:data<=16'd10680;
      67178:data<=16'd11130;
      67179:data<=16'd10998;
      67180:data<=16'd10918;
      67181:data<=16'd11696;
      67182:data<=16'd11753;
      67183:data<=16'd11121;
      67184:data<=16'd11260;
      67185:data<=16'd11039;
      67186:data<=16'd10748;
      67187:data<=16'd11715;
      67188:data<=16'd12073;
      67189:data<=16'd11526;
      67190:data<=16'd11441;
      67191:data<=16'd10881;
      67192:data<=16'd10105;
      67193:data<=16'd10671;
      67194:data<=16'd11500;
      67195:data<=16'd11142;
      67196:data<=16'd10789;
      67197:data<=16'd10749;
      67198:data<=16'd9812;
      67199:data<=16'd9973;
      67200:data<=16'd11486;
      67201:data<=16'd11265;
      67202:data<=16'd10971;
      67203:data<=16'd9881;
      67204:data<=16'd4814;
      67205:data<=16'd2256;
      67206:data<=16'd4388;
      67207:data<=16'd4676;
      67208:data<=16'd4598;
      67209:data<=16'd5386;
      67210:data<=16'd4056;
      67211:data<=16'd3556;
      67212:data<=16'd4949;
      67213:data<=16'd5644;
      67214:data<=16'd5621;
      67215:data<=16'd5186;
      67216:data<=16'd4983;
      67217:data<=16'd4834;
      67218:data<=16'd4730;
      67219:data<=16'd5641;
      67220:data<=16'd5667;
      67221:data<=16'd5327;
      67222:data<=16'd6061;
      67223:data<=16'd5225;
      67224:data<=16'd4728;
      67225:data<=16'd6485;
      67226:data<=16'd6766;
      67227:data<=16'd5976;
      67228:data<=16'd5839;
      67229:data<=16'd5427;
      67230:data<=16'd5674;
      67231:data<=16'd6945;
      67232:data<=16'd7527;
      67233:data<=16'd6440;
      67234:data<=16'd5702;
      67235:data<=16'd5849;
      67236:data<=16'd4860;
      67237:data<=16'd7248;
      67238:data<=16'd13207;
      67239:data<=16'd13743;
      67240:data<=16'd11743;
      67241:data<=16'd12266;
      67242:data<=16'd10963;
      67243:data<=16'd10298;
      67244:data<=16'd11825;
      67245:data<=16'd11602;
      67246:data<=16'd11364;
      67247:data<=16'd10912;
      67248:data<=16'd9517;
      67249:data<=16'd9398;
      67250:data<=16'd8942;
      67251:data<=16'd8335;
      67252:data<=16'd8231;
      67253:data<=16'd7303;
      67254:data<=16'd7259;
      67255:data<=16'd6858;
      67256:data<=16'd4819;
      67257:data<=16'd3852;
      67258:data<=16'd3398;
      67259:data<=16'd2924;
      67260:data<=16'd2924;
      67261:data<=16'd2249;
      67262:data<=16'd1152;
      67263:data<=-16'd235;
      67264:data<=-16'd992;
      67265:data<=-16'd726;
      67266:data<=-16'd1087;
      67267:data<=-16'd1086;
      67268:data<=-16'd1406;
      67269:data<=-16'd2708;
      67270:data<=-16'd3177;
      67271:data<=-16'd6311;
      67272:data<=-16'd10571;
      67273:data<=-16'd9937;
      67274:data<=-16'd9427;
      67275:data<=-16'd11324;
      67276:data<=-16'd11365;
      67277:data<=-16'd11373;
      67278:data<=-16'd11480;
      67279:data<=-16'd10395;
      67280:data<=-16'd10572;
      67281:data<=-16'd11646;
      67282:data<=-16'd12028;
      67283:data<=-16'd11671;
      67284:data<=-16'd11122;
      67285:data<=-16'd11038;
      67286:data<=-16'd10953;
      67287:data<=-16'd11524;
      67288:data<=-16'd12320;
      67289:data<=-16'd11724;
      67290:data<=-16'd11449;
      67291:data<=-16'd11538;
      67292:data<=-16'd10580;
      67293:data<=-16'd10436;
      67294:data<=-16'd11332;
      67295:data<=-16'd11450;
      67296:data<=-16'd10878;
      67297:data<=-16'd10496;
      67298:data<=-16'd9982;
      67299:data<=-16'd9670;
      67300:data<=-16'd11200;
      67301:data<=-16'd12135;
      67302:data<=-16'd11132;
      67303:data<=-16'd11492;
      67304:data<=-16'd9467;
      67305:data<=-16'd3977;
      67306:data<=-16'd3582;
      67307:data<=-16'd5890;
      67308:data<=-16'd4911;
      67309:data<=-16'd4607;
      67310:data<=-16'd4851;
      67311:data<=-16'd3765;
      67312:data<=-16'd4156;
      67313:data<=-16'd5344;
      67314:data<=-16'd5474;
      67315:data<=-16'd5280;
      67316:data<=-16'd5215;
      67317:data<=-16'd4830;
      67318:data<=-16'd4746;
      67319:data<=-16'd5941;
      67320:data<=-16'd6208;
      67321:data<=-16'd5278;
      67322:data<=-16'd5488;
      67323:data<=-16'd5203;
      67324:data<=-16'd4981;
      67325:data<=-16'd6422;
      67326:data<=-16'd6578;
      67327:data<=-16'd5999;
      67328:data<=-16'd6024;
      67329:data<=-16'd5388;
      67330:data<=-16'd5372;
      67331:data<=-16'd6068;
      67332:data<=-16'd6625;
      67333:data<=-16'd6768;
      67334:data<=-16'd6100;
      67335:data<=-16'd5924;
      67336:data<=-16'd4864;
      67337:data<=-16'd4658;
      67338:data<=-16'd9881;
      67339:data<=-16'd13711;
      67340:data<=-16'd12187;
      67341:data<=-16'd11317;
      67342:data<=-16'd10551;
      67343:data<=-16'd9990;
      67344:data<=-16'd11676;
      67345:data<=-16'd11681;
      67346:data<=-16'd10636;
      67347:data<=-16'd10602;
      67348:data<=-16'd9814;
      67349:data<=-16'd9245;
      67350:data<=-16'd8737;
      67351:data<=-16'd7494;
      67352:data<=-16'd7043;
      67353:data<=-16'd7206;
      67354:data<=-16'd7254;
      67355:data<=-16'd6346;
      67356:data<=-16'd4299;
      67357:data<=-16'd2939;
      67358:data<=-16'd2575;
      67359:data<=-16'd2322;
      67360:data<=-16'd1988;
      67361:data<=-16'd1727;
      67362:data<=-16'd728;
      67363:data<=16'd1445;
      67364:data<=16'd2008;
      67365:data<=16'd1582;
      67366:data<=16'd2497;
      67367:data<=16'd2027;
      67368:data<=16'd2132;
      67369:data<=16'd4303;
      67370:data<=16'd3946;
      67371:data<=16'd5462;
      67372:data<=16'd10668;
      67373:data<=16'd11539;
      67374:data<=16'd10454;
      67375:data<=16'd11888;
      67376:data<=16'd12549;
      67377:data<=16'd12349;
      67378:data<=16'd12134;
      67379:data<=16'd11590;
      67380:data<=16'd11244;
      67381:data<=16'd11329;
      67382:data<=16'd12548;
      67383:data<=16'd12977;
      67384:data<=16'd11981;
      67385:data<=16'd11911;
      67386:data<=16'd11677;
      67387:data<=16'd11964;
      67388:data<=16'd13585;
      67389:data<=16'd13218;
      67390:data<=16'd12317;
      67391:data<=16'd12490;
      67392:data<=16'd11638;
      67393:data<=16'd11499;
      67394:data<=16'd12754;
      67395:data<=16'd13133;
      67396:data<=16'd12461;
      67397:data<=16'd11544;
      67398:data<=16'd11227;
      67399:data<=16'd11465;
      67400:data<=16'd12304;
      67401:data<=16'd13165;
      67402:data<=16'd12393;
      67403:data<=16'd12172;
      67404:data<=16'd11711;
      67405:data<=16'd7204;
      67406:data<=16'd4378;
      67407:data<=16'd6156;
      67408:data<=16'd6361;
      67409:data<=16'd5702;
      67410:data<=16'd6149;
      67411:data<=16'd5266;
      67412:data<=16'd5134;
      67413:data<=16'd6684;
      67414:data<=16'd6972;
      67415:data<=16'd6422;
      67416:data<=16'd6200;
      67417:data<=16'd5645;
      67418:data<=16'd5664;
      67419:data<=16'd7062;
      67420:data<=16'd7547;
      67421:data<=16'd6363;
      67422:data<=16'd6028;
      67423:data<=16'd6261;
      67424:data<=16'd6020;
      67425:data<=16'd6828;
      67426:data<=16'd7726;
      67427:data<=16'd7283;
      67428:data<=16'd6978;
      67429:data<=16'd6843;
      67430:data<=16'd6024;
      67431:data<=16'd6003;
      67432:data<=16'd7509;
      67433:data<=16'd7887;
      67434:data<=16'd6493;
      67435:data<=16'd6352;
      67436:data<=16'd6253;
      67437:data<=16'd5272;
      67438:data<=16'd8270;
      67439:data<=16'd13103;
      67440:data<=16'd13621;
      67441:data<=16'd12410;
      67442:data<=16'd11920;
      67443:data<=16'd11536;
      67444:data<=16'd12290;
      67445:data<=16'd12387;
      67446:data<=16'd11323;
      67447:data<=16'd11324;
      67448:data<=16'd10939;
      67449:data<=16'd9784;
      67450:data<=16'd9388;
      67451:data<=16'd8836;
      67452:data<=16'd8211;
      67453:data<=16'd7859;
      67454:data<=16'd7250;
      67455:data<=16'd6962;
      67456:data<=16'd5956;
      67457:data<=16'd3909;
      67458:data<=16'd3136;
      67459:data<=16'd3027;
      67460:data<=16'd2523;
      67461:data<=16'd2731;
      67462:data<=16'd2003;
      67463:data<=-16'd306;
      67464:data<=-16'd1293;
      67465:data<=-16'd1303;
      67466:data<=-16'd1528;
      67467:data<=-16'd933;
      67468:data<=-16'd1489;
      67469:data<=-16'd3609;
      67470:data<=-16'd3654;
      67471:data<=-16'd4032;
      67472:data<=-16'd8247;
      67473:data<=-16'd11224;
      67474:data<=-16'd10507;
      67475:data<=-16'd10651;
      67476:data<=-16'd11850;
      67477:data<=-16'd11670;
      67478:data<=-16'd11582;
      67479:data<=-16'd11805;
      67480:data<=-16'd10986;
      67481:data<=-16'd11077;
      67482:data<=-16'd12504;
      67483:data<=-16'd12542;
      67484:data<=-16'd11990;
      67485:data<=-16'd11961;
      67486:data<=-16'd11015;
      67487:data<=-16'd11166;
      67488:data<=-16'd13198;
      67489:data<=-16'd13370;
      67490:data<=-16'd12128;
      67491:data<=-16'd11793;
      67492:data<=-16'd11555;
      67493:data<=-16'd11723;
      67494:data<=-16'd12690;
      67495:data<=-16'd13282;
      67496:data<=-16'd12895;
      67497:data<=-16'd12102;
      67498:data<=-16'd11869;
      67499:data<=-16'd11359;
      67500:data<=-16'd11517;
      67501:data<=-16'd13773;
      67502:data<=-16'd13656;
      67503:data<=-16'd11972;
      67504:data<=-16'd13015;
      67505:data<=-16'd10602;
      67506:data<=-16'd5439;
      67507:data<=-16'd5920;
      67508:data<=-16'd7259;
      67509:data<=-16'd6123;
      67510:data<=-16'd6337;
      67511:data<=-16'd5900;
      67512:data<=-16'd5797;
      67513:data<=-16'd7592;
      67514:data<=-16'd7551;
      67515:data<=-16'd6834;
      67516:data<=-16'd6962;
      67517:data<=-16'd6448;
      67518:data<=-16'd6394;
      67519:data<=-16'd7136;
      67520:data<=-16'd7896;
      67521:data<=-16'd7920;
      67522:data<=-16'd7241;
      67523:data<=-16'd7177;
      67524:data<=-16'd6692;
      67525:data<=-16'd6678;
      67526:data<=-16'd8489;
      67527:data<=-16'd8501;
      67528:data<=-16'd7291;
      67529:data<=-16'd7262;
      67530:data<=-16'd6584;
      67531:data<=-16'd6827;
      67532:data<=-16'd8446;
      67533:data<=-16'd8285;
      67534:data<=-16'd7506;
      67535:data<=-16'd7755;
      67536:data<=-16'd7580;
      67537:data<=-16'd6667;
      67538:data<=-16'd8178;
      67539:data<=-16'd12745;
      67540:data<=-16'd14674;
      67541:data<=-16'd13665;
      67542:data<=-16'd13446;
      67543:data<=-16'd12311;
      67544:data<=-16'd11888;
      67545:data<=-16'd13417;
      67546:data<=-16'd12942;
      67547:data<=-16'd12117;
      67548:data<=-16'd12132;
      67549:data<=-16'd11106;
      67550:data<=-16'd10639;
      67551:data<=-16'd10210;
      67552:data<=-16'd9483;
      67553:data<=-16'd9189;
      67554:data<=-16'd8254;
      67555:data<=-16'd8343;
      67556:data<=-16'd7896;
      67557:data<=-16'd5018;
      67558:data<=-16'd4112;
      67559:data<=-16'd4410;
      67560:data<=-16'd3682;
      67561:data<=-16'd3997;
      67562:data<=-16'd3462;
      67563:data<=-16'd1397;
      67564:data<=-16'd237;
      67565:data<=16'd53;
      67566:data<=16'd223;
      67567:data<=16'd469;
      67568:data<=-16'd5;
      67569:data<=16'd785;
      67570:data<=16'd3316;
      67571:data<=16'd2919;
      67572:data<=16'd4018;
      67573:data<=16'd9439;
      67574:data<=16'd10248;
      67575:data<=16'd9132;
      67576:data<=16'd11236;
      67577:data<=16'd10974;
      67578:data<=16'd10342;
      67579:data<=16'd11072;
      67580:data<=16'd9820;
      67581:data<=16'd10055;
      67582:data<=16'd11699;
      67583:data<=16'd11618;
      67584:data<=16'd11247;
      67585:data<=16'd10517;
      67586:data<=16'd9967;
      67587:data<=16'd10463;
      67588:data<=16'd11082;
      67589:data<=16'd11788;
      67590:data<=16'd11574;
      67591:data<=16'd11071;
      67592:data<=16'd10963;
      67593:data<=16'd9840;
      67594:data<=16'd10308;
      67595:data<=16'd12436;
      67596:data<=16'd12064;
      67597:data<=16'd10907;
      67598:data<=16'd10666;
      67599:data<=16'd9832;
      67600:data<=16'd10075;
      67601:data<=16'd11841;
      67602:data<=16'd12084;
      67603:data<=16'd11033;
      67604:data<=16'd11191;
      67605:data<=16'd10090;
      67606:data<=16'd6146;
      67607:data<=16'd4632;
      67608:data<=16'd5752;
      67609:data<=16'd5181;
      67610:data<=16'd4807;
      67611:data<=16'd5101;
      67612:data<=16'd4387;
      67613:data<=16'd5043;
      67614:data<=16'd6425;
      67615:data<=16'd6061;
      67616:data<=16'd5530;
      67617:data<=16'd5585;
      67618:data<=16'd5143;
      67619:data<=16'd5309;
      67620:data<=16'd6898;
      67621:data<=16'd7283;
      67622:data<=16'd6162;
      67623:data<=16'd6114;
      67624:data<=16'd5946;
      67625:data<=16'd5770;
      67626:data<=16'd7047;
      67627:data<=16'd6913;
      67628:data<=16'd6143;
      67629:data<=16'd6695;
      67630:data<=16'd6194;
      67631:data<=16'd5871;
      67632:data<=16'd6777;
      67633:data<=16'd7160;
      67634:data<=16'd7219;
      67635:data<=16'd6523;
      67636:data<=16'd6003;
      67637:data<=16'd5835;
      67638:data<=16'd5212;
      67639:data<=16'd8291;
      67640:data<=16'd13051;
      67641:data<=16'd13335;
      67642:data<=16'd12134;
      67643:data<=16'd11386;
      67644:data<=16'd10901;
      67645:data<=16'd12269;
      67646:data<=16'd12398;
      67647:data<=16'd11166;
      67648:data<=16'd11157;
      67649:data<=16'd10652;
      67650:data<=16'd9867;
      67651:data<=16'd9100;
      67652:data<=16'd7946;
      67653:data<=16'd8008;
      67654:data<=16'd8088;
      67655:data<=16'd7430;
      67656:data<=16'd6508;
      67657:data<=16'd4513;
      67658:data<=16'd3351;
      67659:data<=16'd3465;
      67660:data<=16'd2804;
      67661:data<=16'd2312;
      67662:data<=16'd2491;
      67663:data<=16'd1619;
      67664:data<=-16'd450;
      67665:data<=-16'd1368;
      67666:data<=-16'd858;
      67667:data<=-16'd1064;
      67668:data<=-16'd967;
      67669:data<=-16'd1366;
      67670:data<=-16'd3532;
      67671:data<=-16'd3342;
      67672:data<=-16'd3689;
      67673:data<=-16'd8234;
      67674:data<=-16'd10146;
      67675:data<=-16'd9818;
      67676:data<=-16'd11462;
      67677:data<=-16'd11571;
      67678:data<=-16'd10822;
      67679:data<=-16'd10934;
      67680:data<=-16'd10316;
      67681:data<=-16'd10378;
      67682:data<=-16'd11317;
      67683:data<=-16'd11943;
      67684:data<=-16'd11843;
      67685:data<=-16'd11206;
      67686:data<=-16'd11088;
      67687:data<=-16'd10278;
      67688:data<=-16'd10175;
      67689:data<=-16'd12170;
      67690:data<=-16'd11835;
      67691:data<=-16'd10584;
      67692:data<=-16'd11088;
      67693:data<=-16'd10252;
      67694:data<=-16'd10457;
      67695:data<=-16'd12363;
      67696:data<=-16'd12069;
      67697:data<=-16'd11312;
      67698:data<=-16'd10728;
      67699:data<=-16'd9950;
      67700:data<=-16'd10704;
      67701:data<=-16'd11709;
      67702:data<=-16'd12258;
      67703:data<=-16'd11808;
      67704:data<=-16'd10930;
      67705:data<=-16'd11502;
      67706:data<=-16'd9229;
      67707:data<=-16'd4857;
      67708:data<=-16'd4969;
      67709:data<=-16'd5714;
      67710:data<=-16'd4481;
      67711:data<=-16'd4648;
      67712:data<=-16'd4405;
      67713:data<=-16'd4569;
      67714:data<=-16'd6470;
      67715:data<=-16'd6299;
      67716:data<=-16'd5236;
      67717:data<=-16'd5409;
      67718:data<=-16'd5184;
      67719:data<=-16'd5583;
      67720:data<=-16'd6664;
      67721:data<=-16'd6623;
      67722:data<=-16'd6513;
      67723:data<=-16'd6648;
      67724:data<=-16'd6006;
      67725:data<=-16'd5717;
      67726:data<=-16'd6463;
      67727:data<=-16'd6989;
      67728:data<=-16'd6898;
      67729:data<=-16'd6482;
      67730:data<=-16'd5777;
      67731:data<=-16'd5413;
      67732:data<=-16'd5982;
      67733:data<=-16'd7063;
      67734:data<=-16'd7119;
      67735:data<=-16'd5990;
      67736:data<=-16'd5897;
      67737:data<=-16'd5920;
      67738:data<=-16'd4928;
      67739:data<=-16'd7100;
      67740:data<=-16'd11712;
      67741:data<=-16'd13198;
      67742:data<=-16'd12446;
      67743:data<=-16'd11606;
      67744:data<=-16'd10910;
      67745:data<=-16'd11597;
      67746:data<=-16'd11985;
      67747:data<=-16'd11057;
      67748:data<=-16'd10652;
      67749:data<=-16'd10232;
      67750:data<=-16'd9389;
      67751:data<=-16'd8736;
      67752:data<=-16'd8029;
      67753:data<=-16'd7629;
      67754:data<=-16'd7203;
      67755:data<=-16'd6751;
      67756:data<=-16'd6636;
      67757:data<=-16'd5260;
      67758:data<=-16'd3196;
      67759:data<=-16'd2611;
      67760:data<=-16'd2593;
      67761:data<=-16'd2319;
      67762:data<=-16'd2138;
      67763:data<=-16'd1178;
      67764:data<=16'd660;
      67765:data<=16'd1651;
      67766:data<=16'd1371;
      67767:data<=16'd1359;
      67768:data<=16'd1585;
      67769:data<=16'd1938;
      67770:data<=16'd3765;
      67771:data<=16'd4657;
      67772:data<=16'd3480;
      67773:data<=16'd5588;
      67774:data<=16'd10329;
      67775:data<=16'd11570;
      67776:data<=16'd11257;
      67777:data<=16'd12527;
      67778:data<=16'd12690;
      67779:data<=16'd11755;
      67780:data<=16'd11535;
      67781:data<=16'd11129;
      67782:data<=16'd11402;
      67783:data<=16'd12892;
      67784:data<=16'd12837;
      67785:data<=16'd11762;
      67786:data<=16'd11764;
      67787:data<=16'd11514;
      67788:data<=16'd11567;
      67789:data<=16'd12813;
      67790:data<=16'd12819;
      67791:data<=16'd12022;
      67792:data<=16'd11900;
      67793:data<=16'd11482;
      67794:data<=16'd11676;
      67795:data<=16'd12825;
      67796:data<=16'd13107;
      67797:data<=16'd12587;
      67798:data<=16'd12093;
      67799:data<=16'd11732;
      67800:data<=16'd11442;
      67801:data<=16'd12070;
      67802:data<=16'd13676;
      67803:data<=16'd13195;
      67804:data<=16'd11773;
      67805:data<=16'd12554;
      67806:data<=16'd11082;
      67807:data<=16'd7018;
      67808:data<=16'd6106;
      67809:data<=16'd6422;
      67810:data<=16'd5974;
      67811:data<=16'd6231;
      67812:data<=16'd5651;
      67813:data<=16'd5711;
      67814:data<=16'd7289;
      67815:data<=16'd7316;
      67816:data<=16'd7001;
      67817:data<=16'd7312;
      67818:data<=16'd6731;
      67819:data<=16'd6605;
      67820:data<=16'd7486;
      67821:data<=16'd8150;
      67822:data<=16'd7999;
      67823:data<=16'd7541;
      67824:data<=16'd7683;
      67825:data<=16'd7333;
      67826:data<=16'd7188;
      67827:data<=16'd8392;
      67828:data<=16'd8211;
      67829:data<=16'd7420;
      67830:data<=16'd7641;
      67831:data<=16'd6822;
      67832:data<=16'd6830;
      67833:data<=16'd8190;
      67834:data<=16'd8167;
      67835:data<=16'd8153;
      67836:data<=16'd7852;
      67837:data<=16'd6616;
      67838:data<=16'd6654;
      67839:data<=16'd7144;
      67840:data<=16'd9271;
      67841:data<=16'd13596;
      67842:data<=16'd14551;
      67843:data<=16'd12536;
      67844:data<=16'd12175;
      67845:data<=16'd12771;
      67846:data<=16'd13173;
      67847:data<=16'd12979;
      67848:data<=16'd12054;
      67849:data<=16'd11558;
      67850:data<=16'd11188;
      67851:data<=16'd10495;
      67852:data<=16'd9767;
      67853:data<=16'd9172;
      67854:data<=16'd8972;
      67855:data<=16'd8569;
      67856:data<=16'd7921;
      67857:data<=16'd6775;
      67858:data<=16'd4702;
      67859:data<=16'd3812;
      67860:data<=16'd4009;
      67861:data<=16'd3460;
      67862:data<=16'd3342;
      67863:data<=16'd3015;
      67864:data<=16'd1363;
      67865:data<=16'd472;
      67866:data<=16'd455;
      67867:data<=16'd206;
      67868:data<=16'd199;
      67869:data<=16'd64;
      67870:data<=-16'd1281;
      67871:data<=-16'd2651;
      67872:data<=-16'd2147;
      67873:data<=-16'd3115;
      67874:data<=-16'd7491;
      67875:data<=-16'd9495;
      67876:data<=-16'd9141;
      67877:data<=-16'd10713;
      67878:data<=-16'd11089;
      67879:data<=-16'd10049;
      67880:data<=-16'd10342;
      67881:data<=-16'd9814;
      67882:data<=-16'd9653;
      67883:data<=-16'd11303;
      67884:data<=-16'd11576;
      67885:data<=-16'd10900;
      67886:data<=-16'd10663;
      67887:data<=-16'd9922;
      67888:data<=-16'd9881;
      67889:data<=-16'd11139;
      67890:data<=-16'd11579;
      67891:data<=-16'd10658;
      67892:data<=-16'd10232;
      67893:data<=-16'd10298;
      67894:data<=-16'd9882;
      67895:data<=-16'd10618;
      67896:data<=-16'd11888;
      67897:data<=-16'd11403;
      67898:data<=-16'd10953;
      67899:data<=-16'd10822;
      67900:data<=-16'd9805;
      67901:data<=-16'd10178;
      67902:data<=-16'd11768;
      67903:data<=-16'd12082;
      67904:data<=-16'd11488;
      67905:data<=-16'd11204;
      67906:data<=-16'd11195;
      67907:data<=-16'd9392;
      67908:data<=-16'd5970;
      67909:data<=-16'd5002;
      67910:data<=-16'd5858;
      67911:data<=-16'd5316;
      67912:data<=-16'd4701;
      67913:data<=-16'd5027;
      67914:data<=-16'd5855;
      67915:data<=-16'd6927;
      67916:data<=-16'd6783;
      67917:data<=-16'd6087;
      67918:data<=-16'd6131;
      67919:data<=-16'd5893;
      67920:data<=-16'd6253;
      67921:data<=-16'd7626;
      67922:data<=-16'd7726;
      67923:data<=-16'd7230;
      67924:data<=-16'd7204;
      67925:data<=-16'd6663;
      67926:data<=-16'd7101;
      67927:data<=-16'd8454;
      67928:data<=-16'd8228;
      67929:data<=-16'd7783;
      67930:data<=-16'd7699;
      67931:data<=-16'd6713;
      67932:data<=-16'd6872;
      67933:data<=-16'd8123;
      67934:data<=-16'd8413;
      67935:data<=-16'd8373;
      67936:data<=-16'd7800;
      67937:data<=-16'd7013;
      67938:data<=-16'd7047;
      67939:data<=-16'd7148;
      67940:data<=-16'd9103;
      67941:data<=-16'd13077;
      67942:data<=-16'd14603;
      67943:data<=-16'd13530;
      67944:data<=-16'd12771;
      67945:data<=-16'd12904;
      67946:data<=-16'd13574;
      67947:data<=-16'd13565;
      67948:data<=-16'd12786;
      67949:data<=-16'd12161;
      67950:data<=-16'd11450;
      67951:data<=-16'd10840;
      67952:data<=-16'd10284;
      67953:data<=-16'd9712;
      67954:data<=-16'd9430;
      67955:data<=-16'd8715;
      67956:data<=-16'd8164;
      67957:data<=-16'd7649;
      67958:data<=-16'd5771;
      67959:data<=-16'd4575;
      67960:data<=-16'd4560;
      67961:data<=-16'd3853;
      67962:data<=-16'd3718;
      67963:data<=-16'd3842;
      67964:data<=-16'd2457;
      67965:data<=-16'd945;
      67966:data<=-16'd500;
      67967:data<=-16'd604;
      67968:data<=-16'd403;
      67969:data<=-16'd59;
      67970:data<=16'd429;
      67971:data<=16'd2184;
      67972:data<=16'd2731;
      67973:data<=16'd1589;
      67974:data<=16'd4228;
      67975:data<=16'd8683;
      67976:data<=16'd9555;
      67977:data<=16'd9796;
      67978:data<=16'd10787;
      67979:data<=16'd10454;
      67980:data<=16'd9988;
      67981:data<=16'd9758;
      67982:data<=16'd9652;
      67983:data<=16'd10543;
      67984:data<=16'd11203;
      67985:data<=16'd10824;
      67986:data<=16'd10292;
      67987:data<=16'd9752;
      67988:data<=16'd9420;
      67989:data<=16'd10141;
      67990:data<=16'd11051;
      67991:data<=16'd10543;
      67992:data<=16'd9912;
      67993:data<=16'd10038;
      67994:data<=16'd9583;
      67995:data<=16'd9831;
      67996:data<=16'd11177;
      67997:data<=16'd11136;
      67998:data<=16'd10557;
      67999:data<=16'd10511;
      68000:data<=16'd10058;
      68001:data<=16'd10246;
      68002:data<=16'd11133;
      68003:data<=16'd11327;
      68004:data<=16'd10957;
      68005:data<=16'd10683;
      68006:data<=16'd10646;
      68007:data<=16'd8983;
      68008:data<=16'd5673;
      68009:data<=16'd4496;
      68010:data<=16'd4802;
      68011:data<=16'd4126;
      68012:data<=16'd3940;
      68013:data<=16'd4040;
      68014:data<=16'd4332;
      68015:data<=16'd5644;
      68016:data<=16'd5664;
      68017:data<=16'd5087;
      68018:data<=16'd5554;
      68019:data<=16'd5037;
      68020:data<=16'd5080;
      68021:data<=16'd6675;
      68022:data<=16'd6687;
      68023:data<=16'd6246;
      68024:data<=16'd6488;
      68025:data<=16'd5671;
      68026:data<=16'd5588;
      68027:data<=16'd6912;
      68028:data<=16'd7241;
      68029:data<=16'd6837;
      68030:data<=16'd6351;
      68031:data<=16'd5439;
      68032:data<=16'd5439;
      68033:data<=16'd6693;
      68034:data<=16'd7131;
      68035:data<=16'd6539;
      68036:data<=16'd6551;
      68037:data<=16'd6475;
      68038:data<=16'd5648;
      68039:data<=16'd5556;
      68040:data<=16'd6529;
      68041:data<=16'd9033;
      68042:data<=16'd12414;
      68043:data<=16'd12725;
      68044:data<=16'd10950;
      68045:data<=16'd11388;
      68046:data<=16'd12357;
      68047:data<=16'd12025;
      68048:data<=16'd11614;
      68049:data<=16'd10713;
      68050:data<=16'd9699;
      68051:data<=16'd9515;
      68052:data<=16'd9201;
      68053:data<=16'd8388;
      68054:data<=16'd7550;
      68055:data<=16'd6963;
      68056:data<=16'd6655;
      68057:data<=16'd6005;
      68058:data<=16'd4622;
      68059:data<=16'd3228;
      68060:data<=16'd2805;
      68061:data<=16'd2598;
      68062:data<=16'd1760;
      68063:data<=16'd1562;
      68064:data<=16'd1306;
      68065:data<=-16'd420;
      68066:data<=-16'd1272;
      68067:data<=-16'd902;
      68068:data<=-16'd1434;
      68069:data<=-16'd1738;
      68070:data<=-16'd1847;
      68071:data<=-16'd3585;
      68072:data<=-16'd4558;
      68073:data<=-16'd3644;
      68074:data<=-16'd5247;
      68075:data<=-16'd9459;
      68076:data<=-16'd11241;
      68077:data<=-16'd11403;
      68078:data<=-16'd12584;
      68079:data<=-16'd12530;
      68080:data<=-16'd11677;
      68081:data<=-16'd11929;
      68082:data<=-16'd11700;
      68083:data<=-16'd11808;
      68084:data<=-16'd12818;
      68085:data<=-16'd12455;
      68086:data<=-16'd12047;
      68087:data<=-16'd12296;
      68088:data<=-16'd11379;
      68089:data<=-16'd11335;
      68090:data<=-16'd12863;
      68091:data<=-16'd12889;
      68092:data<=-16'd12119;
      68093:data<=-16'd12113;
      68094:data<=-16'd11406;
      68095:data<=-16'd11168;
      68096:data<=-16'd12618;
      68097:data<=-16'd12883;
      68098:data<=-16'd12102;
      68099:data<=-16'd12041;
      68100:data<=-16'd11241;
      68101:data<=-16'd11091;
      68102:data<=-16'd12649;
      68103:data<=-16'd12753;
      68104:data<=-16'd11903;
      68105:data<=-16'd11767;
      68106:data<=-16'd11579;
      68107:data<=-16'd11136;
      68108:data<=-16'd8796;
      68109:data<=-16'd5659;
      68110:data<=-16'd5259;
      68111:data<=-16'd5736;
      68112:data<=-16'd5195;
      68113:data<=-16'd4689;
      68114:data<=-16'd4987;
      68115:data<=-16'd6473;
      68116:data<=-16'd6858;
      68117:data<=-16'd6005;
      68118:data<=-16'd6194;
      68119:data<=-16'd5739;
      68120:data<=-16'd5614;
      68121:data<=-16'd7345;
      68122:data<=-16'd7532;
      68123:data<=-16'd6846;
      68124:data<=-16'd6913;
      68125:data<=-16'd6228;
      68126:data<=-16'd6203;
      68127:data<=-16'd7280;
      68128:data<=-16'd7700;
      68129:data<=-16'd7333;
      68130:data<=-16'd6810;
      68131:data<=-16'd6605;
      68132:data<=-16'd6097;
      68133:data<=-16'd6240;
      68134:data<=-16'd7586;
      68135:data<=-16'd7503;
      68136:data<=-16'd6969;
      68137:data<=-16'd6801;
      68138:data<=-16'd5783;
      68139:data<=-16'd6357;
      68140:data<=-16'd7339;
      68141:data<=-16'd8276;
      68142:data<=-16'd12187;
      68143:data<=-16'd13626;
      68144:data<=-16'd11471;
      68145:data<=-16'd12179;
      68146:data<=-16'd13271;
      68147:data<=-16'd12669;
      68148:data<=-16'd12398;
      68149:data<=-16'd11418;
      68150:data<=-16'd10762;
      68151:data<=-16'd10466;
      68152:data<=-16'd9555;
      68153:data<=-16'd9397;
      68154:data<=-16'd8875;
      68155:data<=-16'd7824;
      68156:data<=-16'd7406;
      68157:data<=-16'd6764;
      68158:data<=-16'd5806;
      68159:data<=-16'd4317;
      68160:data<=-16'd3218;
      68161:data<=-16'd3058;
      68162:data<=-16'd2315;
      68163:data<=-16'd2202;
      68164:data<=-16'd1962;
      68165:data<=-16'd100;
      68166:data<=16'd651;
      68167:data<=16'd1064;
      68168:data<=16'd1642;
      68169:data<=16'd913;
      68170:data<=16'd1671;
      68171:data<=16'd3433;
      68172:data<=16'd4102;
      68173:data<=16'd4270;
      68174:data<=16'd4214;
      68175:data<=16'd7133;
      68176:data<=16'd11254;
      68177:data<=16'd11576;
      68178:data<=16'd11873;
      68179:data<=16'd12818;
      68180:data<=16'd12073;
      68181:data<=16'd12220;
      68182:data<=16'd11846;
      68183:data<=16'd11358;
      68184:data<=16'd13085;
      68185:data<=16'd13182;
      68186:data<=16'd12261;
      68187:data<=16'd12481;
      68188:data<=16'd11559;
      68189:data<=16'd11438;
      68190:data<=16'd13050;
      68191:data<=16'd13280;
      68192:data<=16'd12527;
      68193:data<=16'd12239;
      68194:data<=16'd11882;
      68195:data<=16'd11734;
      68196:data<=16'd12880;
      68197:data<=16'd13628;
      68198:data<=16'd12598;
      68199:data<=16'd12384;
      68200:data<=16'd12334;
      68201:data<=16'd11130;
      68202:data<=16'd11796;
      68203:data<=16'd13091;
      68204:data<=16'd12857;
      68205:data<=16'd12645;
      68206:data<=16'd12096;
      68207:data<=16'd11424;
      68208:data<=16'd10110;
      68209:data<=16'd7134;
      68210:data<=16'd5836;
      68211:data<=16'd6249;
      68212:data<=16'd5618;
      68213:data<=16'd4968;
      68214:data<=16'd5251;
      68215:data<=16'd6567;
      68216:data<=16'd7374;
      68217:data<=16'd6516;
      68218:data<=16'd6319;
      68219:data<=16'd6310;
      68220:data<=16'd5982;
      68221:data<=16'd7241;
      68222:data<=16'd8008;
      68223:data<=16'd7485;
      68224:data<=16'd7606;
      68225:data<=16'd7420;
      68226:data<=16'd6622;
      68227:data<=16'd6790;
      68228:data<=16'd8081;
      68229:data<=16'd8560;
      68230:data<=16'd7908;
      68231:data<=16'd7682;
      68232:data<=16'd6766;
      68233:data<=16'd6536;
      68234:data<=16'd8716;
      68235:data<=16'd8869;
      68236:data<=16'd7741;
      68237:data<=16'd8000;
      68238:data<=16'd6990;
      68239:data<=16'd7080;
      68240:data<=16'd8537;
      68241:data<=16'd8533;
      68242:data<=16'd11050;
      68243:data<=16'd14202;
      68244:data<=16'd13443;
      68245:data<=16'd12853;
      68246:data<=16'd13632;
      68247:data<=16'd13952;
      68248:data<=16'd13850;
      68249:data<=16'd12824;
      68250:data<=16'd12028;
      68251:data<=16'd11611;
      68252:data<=16'd10915;
      68253:data<=16'd10555;
      68254:data<=16'd9776;
      68255:data<=16'd8907;
      68256:data<=16'd8570;
      68257:data<=16'd8266;
      68258:data<=16'd7479;
      68259:data<=16'd5344;
      68260:data<=16'd4196;
      68261:data<=16'd4514;
      68262:data<=16'd3577;
      68263:data<=16'd3645;
      68264:data<=16'd3850;
      68265:data<=16'd1471;
      68266:data<=16'd502;
      68267:data<=16'd684;
      68268:data<=-16'd105;
      68269:data<=-16'd138;
      68270:data<=-16'd467;
      68271:data<=-16'd1180;
      68272:data<=-16'd2259;
      68273:data<=-16'd3486;
      68274:data<=-16'd2711;
      68275:data<=-16'd4232;
      68276:data<=-16'd8595;
      68277:data<=-16'd9999;
      68278:data<=-16'd10881;
      68279:data<=-16'd12037;
      68280:data<=-16'd11173;
      68281:data<=-16'd11054;
      68282:data<=-16'd10831;
      68283:data<=-16'd10571;
      68284:data<=-16'd12143;
      68285:data<=-16'd12289;
      68286:data<=-16'd11555;
      68287:data<=-16'd11570;
      68288:data<=-16'd10737;
      68289:data<=-16'd10769;
      68290:data<=-16'd11888;
      68291:data<=-16'd12188;
      68292:data<=-16'd11932;
      68293:data<=-16'd11656;
      68294:data<=-16'd11546;
      68295:data<=-16'd10781;
      68296:data<=-16'd10748;
      68297:data<=-16'd12530;
      68298:data<=-16'd12640;
      68299:data<=-16'd11790;
      68300:data<=-16'd11618;
      68301:data<=-16'd10217;
      68302:data<=-16'd10423;
      68303:data<=-16'd12373;
      68304:data<=-16'd12202;
      68305:data<=-16'd11591;
      68306:data<=-16'd11241;
      68307:data<=-16'd10610;
      68308:data<=-16'd10310;
      68309:data<=-16'd8105;
      68310:data<=-16'd5180;
      68311:data<=-16'd4602;
      68312:data<=-16'd4855;
      68313:data<=-16'd4499;
      68314:data<=-16'd4071;
      68315:data<=-16'd4868;
      68316:data<=-16'd6143;
      68317:data<=-16'd5783;
      68318:data<=-16'd5548;
      68319:data<=-16'd5698;
      68320:data<=-16'd4742;
      68321:data<=-16'd5281;
      68322:data<=-16'd6892;
      68323:data<=-16'd6807;
      68324:data<=-16'd6466;
      68325:data<=-16'd6294;
      68326:data<=-16'd5644;
      68327:data<=-16'd6046;
      68328:data<=-16'd7365;
      68329:data<=-16'd7512;
      68330:data<=-16'd6772;
      68331:data<=-16'd6704;
      68332:data<=-16'd6399;
      68333:data<=-16'd6279;
      68334:data<=-16'd7753;
      68335:data<=-16'd8000;
      68336:data<=-16'd7142;
      68337:data<=-16'd7617;
      68338:data<=-16'd6945;
      68339:data<=-16'd6325;
      68340:data<=-16'd7694;
      68341:data<=-16'd7645;
      68342:data<=-16'd8798;
      68343:data<=-16'd12939;
      68344:data<=-16'd13813;
      68345:data<=-16'd12217;
      68346:data<=-16'd12898;
      68347:data<=-16'd13941;
      68348:data<=-16'd13585;
      68349:data<=-16'd12695;
      68350:data<=-16'd11975;
      68351:data<=-16'd11705;
      68352:data<=-16'd11157;
      68353:data<=-16'd10282;
      68354:data<=-16'd9709;
      68355:data<=-16'd9209;
      68356:data<=-16'd8783;
      68357:data<=-16'd8533;
      68358:data<=-16'd7538;
      68359:data<=-16'd5606;
      68360:data<=-16'd4487;
      68361:data<=-16'd4516;
      68362:data<=-16'd4112;
      68363:data<=-16'd3639;
      68364:data<=-16'd3453;
      68365:data<=-16'd2366;
      68366:data<=-16'd1064;
      68367:data<=-16'd516;
      68368:data<=-16'd58;
      68369:data<=16'd356;
      68370:data<=16'd388;
      68371:data<=16'd869;
      68372:data<=16'd2537;
      68373:data<=16'd3432;
      68374:data<=16'd2544;
      68375:data<=16'd3500;
      68376:data<=16'd7153;
      68377:data<=16'd10067;
      68378:data<=16'd11521;
      68379:data<=16'd11888;
      68380:data<=16'd11491;
      68381:data<=16'd11464;
      68382:data<=16'd11151;
      68383:data<=16'd11021;
      68384:data<=16'd12181;
      68385:data<=16'd12583;
      68386:data<=16'd11855;
      68387:data<=16'd11661;
      68388:data<=16'd11354;
      68389:data<=16'd10701;
      68390:data<=16'd11159;
      68391:data<=16'd12424;
      68392:data<=16'd12464;
      68393:data<=16'd11621;
      68394:data<=16'd11379;
      68395:data<=16'd10810;
      68396:data<=16'd10837;
      68397:data<=16'd12463;
      68398:data<=16'd12522;
      68399:data<=16'd11562;
      68400:data<=16'd11543;
      68401:data<=16'd10510;
      68402:data<=16'd10486;
      68403:data<=16'd12304;
      68404:data<=16'd12122;
      68405:data<=16'd11417;
      68406:data<=16'd11286;
      68407:data<=16'd10337;
      68408:data<=16'd10533;
      68409:data<=16'd9650;
      68410:data<=16'd5797;
      68411:data<=16'd4002;
      68412:data<=16'd4523;
      68413:data<=16'd3999;
      68414:data<=16'd3345;
      68415:data<=16'd3914;
      68416:data<=16'd5162;
      68417:data<=16'd5295;
      68418:data<=16'd4525;
      68419:data<=16'd4622;
      68420:data<=16'd4411;
      68421:data<=16'd4511;
      68422:data<=16'd6043;
      68423:data<=16'd6017;
      68424:data<=16'd5244;
      68425:data<=16'd5786;
      68426:data<=16'd5377;
      68427:data<=16'd4937;
      68428:data<=16'd6061;
      68429:data<=16'd6507;
      68430:data<=16'd6135;
      68431:data<=16'd6087;
      68432:data<=16'd5670;
      68433:data<=16'd5089;
      68434:data<=16'd5830;
      68435:data<=16'd7125;
      68436:data<=16'd6884;
      68437:data<=16'd6267;
      68438:data<=16'd6111;
      68439:data<=16'd5491;
      68440:data<=16'd5967;
      68441:data<=16'd6818;
      68442:data<=16'd7263;
      68443:data<=16'd10340;
      68444:data<=16'd12821;
      68445:data<=16'd11582;
      68446:data<=16'd11661;
      68447:data<=16'd12965;
      68448:data<=16'd12443;
      68449:data<=16'd12055;
      68450:data<=16'd11712;
      68451:data<=16'd10753;
      68452:data<=16'd10204;
      68453:data<=16'd9506;
      68454:data<=16'd8883;
      68455:data<=16'd8557;
      68456:data<=16'd7782;
      68457:data<=16'd7203;
      68458:data<=16'd7050;
      68459:data<=16'd6008;
      68460:data<=16'd4111;
      68461:data<=16'd3316;
      68462:data<=16'd3274;
      68463:data<=16'd2613;
      68464:data<=16'd2670;
      68465:data<=16'd2261;
      68466:data<=16'd117;
      68467:data<=-16'd629;
      68468:data<=-16'd529;
      68469:data<=-16'd1034;
      68470:data<=-16'd801;
      68471:data<=-16'd1656;
      68472:data<=-16'd3322;
      68473:data<=-16'd3879;
      68474:data<=-16'd4146;
      68475:data<=-16'd3582;
      68476:data<=-16'd5049;
      68477:data<=-16'd9981;
      68478:data<=-16'd12245;
      68479:data<=-16'd12014;
      68480:data<=-16'd12642;
      68481:data<=-16'd12367;
      68482:data<=-16'd11849;
      68483:data<=-16'd11734;
      68484:data<=-16'd12073;
      68485:data<=-16'd13561;
      68486:data<=-16'd13432;
      68487:data<=-16'd12416;
      68488:data<=-16'd12508;
      68489:data<=-16'd11749;
      68490:data<=-16'd12070;
      68491:data<=-16'd13803;
      68492:data<=-16'd13344;
      68493:data<=-16'd12471;
      68494:data<=-16'd12522;
      68495:data<=-16'd11963;
      68496:data<=-16'd12073;
      68497:data<=-16'd13071;
      68498:data<=-16'd13077;
      68499:data<=-16'd12417;
      68500:data<=-16'd12375;
      68501:data<=-16'd12010;
      68502:data<=-16'd11229;
      68503:data<=-16'd12138;
      68504:data<=-16'd13195;
      68505:data<=-16'd12539;
      68506:data<=-16'd11984;
      68507:data<=-16'd11465;
      68508:data<=-16'd11176;
      68509:data<=-16'd11082;
      68510:data<=-16'd8355;
      68511:data<=-16'd5426;
      68512:data<=-16'd5410;
      68513:data<=-16'd5285;
      68514:data<=-16'd4523;
      68515:data<=-16'd5059;
      68516:data<=-16'd5996;
      68517:data<=-16'd6043;
      68518:data<=-16'd5702;
      68519:data<=-16'd5915;
      68520:data<=-16'd5712;
      68521:data<=-16'd5535;
      68522:data<=-16'd6831;
      68523:data<=-16'd7256;
      68524:data<=-16'd6581;
      68525:data<=-16'd6570;
      68526:data<=-16'd6119;
      68527:data<=-16'd6155;
      68528:data<=-16'd7219;
      68529:data<=-16'd7551;
      68530:data<=-16'd7435;
      68531:data<=-16'd7028;
      68532:data<=-16'd6626;
      68533:data<=-16'd6511;
      68534:data<=-16'd6698;
      68535:data<=-16'd8047;
      68536:data<=-16'd8076;
      68537:data<=-16'd6960;
      68538:data<=-16'd7573;
      68539:data<=-16'd6781;
      68540:data<=-16'd6208;
      68541:data<=-16'd8137;
      68542:data<=-16'd7371;
      68543:data<=-16'd8179;
      68544:data<=-16'd13051;
      68545:data<=-16'd13305;
      68546:data<=-16'd11887;
      68547:data<=-16'd13658;
      68548:data<=-16'd13843;
      68549:data<=-16'd13010;
      68550:data<=-16'd12596;
      68551:data<=-16'd11550;
      68552:data<=-16'd11367;
      68553:data<=-16'd10978;
      68554:data<=-16'd9882;
      68555:data<=-16'd9444;
      68556:data<=-16'd8751;
      68557:data<=-16'd8258;
      68558:data<=-16'd8296;
      68559:data<=-16'd6889;
      68560:data<=-16'd4604;
      68561:data<=-16'd3835;
      68562:data<=-16'd3967;
      68563:data<=-16'd3448;
      68564:data<=-16'd3125;
      68565:data<=-16'd2393;
      68566:data<=-16'd440;
      68567:data<=16'd249;
      68568:data<=16'd109;
      68569:data<=16'd790;
      68570:data<=16'd977;
      68571:data<=16'd1394;
      68572:data<=16'd2557;
      68573:data<=16'd3539;
      68574:data<=16'd4081;
      68575:data<=16'd3406;
      68576:data<=16'd4375;
      68577:data<=16'd8451;
      68578:data<=16'd11374;
      68579:data<=16'd12555;
      68580:data<=16'd12815;
      68581:data<=16'd12070;
      68582:data<=16'd12101;
      68583:data<=16'd11922;
      68584:data<=16'd12201;
      68585:data<=16'd13902;
      68586:data<=16'd13561;
      68587:data<=16'd12601;
      68588:data<=16'd12596;
      68589:data<=16'd11640;
      68590:data<=16'd12125;
      68591:data<=16'd13483;
      68592:data<=16'd13253;
      68593:data<=16'd13038;
      68594:data<=16'd12528;
      68595:data<=16'd12085;
      68596:data<=16'd12496;
      68597:data<=16'd12816;
      68598:data<=16'd13593;
      68599:data<=16'd13435;
      68600:data<=16'd12719;
      68601:data<=16'd12942;
      68602:data<=16'd11903;
      68603:data<=16'd12257;
      68604:data<=16'd14295;
      68605:data<=16'd13339;
      68606:data<=16'd12888;
      68607:data<=16'd13251;
      68608:data<=16'd11764;
      68609:data<=16'd12652;
      68610:data<=16'd12225;
      68611:data<=16'd7462;
      68612:data<=16'd5921;
      68613:data<=16'd6667;
      68614:data<=16'd5624;
      68615:data<=16'd5724;
      68616:data<=16'd6887;
      68617:data<=16'd7318;
      68618:data<=16'd7203;
      68619:data<=16'd6924;
      68620:data<=16'd6795;
      68621:data<=16'd6569;
      68622:data<=16'd7313;
      68623:data<=16'd8536;
      68624:data<=16'd8181;
      68625:data<=16'd7900;
      68626:data<=16'd8084;
      68627:data<=16'd7338;
      68628:data<=16'd7541;
      68629:data<=16'd8722;
      68630:data<=16'd8828;
      68631:data<=16'd8531;
      68632:data<=16'd8317;
      68633:data<=16'd7650;
      68634:data<=16'd7764;
      68635:data<=16'd8954;
      68636:data<=16'd9053;
      68637:data<=16'd8537;
      68638:data<=16'd8739;
      68639:data<=16'd7908;
      68640:data<=16'd7550;
      68641:data<=16'd8992;
      68642:data<=16'd8687;
      68643:data<=16'd9047;
      68644:data<=16'd12892;
      68645:data<=16'd14530;
      68646:data<=16'd13473;
      68647:data<=16'd13975;
      68648:data<=16'd14571;
      68649:data<=16'd14069;
      68650:data<=16'd13500;
      68651:data<=16'd12875;
      68652:data<=16'd12216;
      68653:data<=16'd11271;
      68654:data<=16'd10502;
      68655:data<=16'd10295;
      68656:data<=16'd9738;
      68657:data<=16'd9037;
      68658:data<=16'd8489;
      68659:data<=16'd7347;
      68660:data<=16'd5783;
      68661:data<=16'd4877;
      68662:data<=16'd4846;
      68663:data<=16'd4513;
      68664:data<=16'd3911;
      68665:data<=16'd3586;
      68666:data<=16'd2317;
      68667:data<=16'd928;
      68668:data<=16'd755;
      68669:data<=16'd328;
      68670:data<=16'd70;
      68671:data<=16'd246;
      68672:data<=-16'd1061;
      68673:data<=-16'd2469;
      68674:data<=-16'd2681;
      68675:data<=-16'd2698;
      68676:data<=-16'd2382;
      68677:data<=-16'd4170;
      68678:data<=-16'd9266;
      68679:data<=-16'd12035;
      68680:data<=-16'd10988;
      68681:data<=-16'd10745;
      68682:data<=-16'd11110;
      68683:data<=-16'd10557;
      68684:data<=-16'd10956;
      68685:data<=-16'd11840;
      68686:data<=-16'd11825;
      68687:data<=-16'd11697;
      68688:data<=-16'd11403;
      68689:data<=-16'd10772;
      68690:data<=-16'd10655;
      68691:data<=-16'd11380;
      68692:data<=-16'd12110;
      68693:data<=-16'd11590;
      68694:data<=-16'd10975;
      68695:data<=-16'd11207;
      68696:data<=-16'd10648;
      68697:data<=-16'd10795;
      68698:data<=-16'd12343;
      68699:data<=-16'd11937;
      68700:data<=-16'd11122;
      68701:data<=-16'd11306;
      68702:data<=-16'd10293;
      68703:data<=-16'd10757;
      68704:data<=-16'd12490;
      68705:data<=-16'd11873;
      68706:data<=-16'd11586;
      68707:data<=-16'd11586;
      68708:data<=-16'd10339;
      68709:data<=-16'd11085;
      68710:data<=-16'd10933;
      68711:data<=-16'd7006;
      68712:data<=-16'd4646;
      68713:data<=-16'd4825;
      68714:data<=-16'd4532;
      68715:data<=-16'd4303;
      68716:data<=-16'd5053;
      68717:data<=-16'd6099;
      68718:data<=-16'd6006;
      68719:data<=-16'd5544;
      68720:data<=-16'd5824;
      68721:data<=-16'd5278;
      68722:data<=-16'd5407;
      68723:data<=-16'd7201;
      68724:data<=-16'd7300;
      68725:data<=-16'd6677;
      68726:data<=-16'd6784;
      68727:data<=-16'd5990;
      68728:data<=-16'd6228;
      68729:data<=-16'd7606;
      68730:data<=-16'd7602;
      68731:data<=-16'd7283;
      68732:data<=-16'd6945;
      68733:data<=-16'd6193;
      68734:data<=-16'd6411;
      68735:data<=-16'd7503;
      68736:data<=-16'd8047;
      68737:data<=-16'd7247;
      68738:data<=-16'd6852;
      68739:data<=-16'd7442;
      68740:data<=-16'd6630;
      68741:data<=-16'd6639;
      68742:data<=-16'd8043;
      68743:data<=-16'd7115;
      68744:data<=-16'd8407;
      68745:data<=-16'd13035;
      68746:data<=-16'd13397;
      68747:data<=-16'd12255;
      68748:data<=-16'd13759;
      68749:data<=-16'd13759;
      68750:data<=-16'd12787;
      68751:data<=-16'd12225;
      68752:data<=-16'd10939;
      68753:data<=-16'd10543;
      68754:data<=-16'd10416;
      68755:data<=-16'd9658;
      68756:data<=-16'd9241;
      68757:data<=-16'd8187;
      68758:data<=-16'd7365;
      68759:data<=-16'd7285;
      68760:data<=-16'd5667;
      68761:data<=-16'd4049;
      68762:data<=-16'd4146;
      68763:data<=-16'd3845;
      68764:data<=-16'd3325;
      68765:data<=-16'd3368;
      68766:data<=-16'd2114;
      68767:data<=-16'd343;
      68768:data<=-16'd118;
      68769:data<=16'd18;
      68770:data<=16'd382;
      68771:data<=16'd102;
      68772:data<=16'd1089;
      68773:data<=16'd2752;
      68774:data<=16'd3112;
      68775:data<=16'd3186;
      68776:data<=16'd2881;
      68777:data<=16'd3999;
      68778:data<=16'd8636;
      68779:data<=16'd11823;
      68780:data<=16'd11606;
      68781:data<=16'd11502;
      68782:data<=16'd11186;
      68783:data<=16'd10637;
      68784:data<=16'd10953;
      68785:data<=16'd11470;
      68786:data<=16'd12116;
      68787:data<=16'd11835;
      68788:data<=16'd11129;
      68789:data<=16'd11286;
      68790:data<=16'd10636;
      68791:data<=16'd10560;
      68792:data<=16'd11843;
      68793:data<=16'd11432;
      68794:data<=16'd10906;
      68795:data<=16'd11207;
      68796:data<=16'd10317;
      68797:data<=16'd10446;
      68798:data<=16'd11814;
      68799:data<=16'd11831;
      68800:data<=16'd11397;
      68801:data<=16'd11010;
      68802:data<=16'd10141;
      68803:data<=16'd10305;
      68804:data<=16'd11873;
      68805:data<=16'd12304;
      68806:data<=16'd11232;
      68807:data<=16'd11142;
      68808:data<=16'd10936;
      68809:data<=16'd10210;
      68810:data<=16'd11388;
      68811:data<=16'd10241;
      68812:data<=16'd5371;
      68813:data<=16'd4076;
      68814:data<=16'd5107;
      68815:data<=16'd3914;
      68816:data<=16'd4108;
      68817:data<=16'd5738;
      68818:data<=16'd5764;
      68819:data<=16'd5570;
      68820:data<=16'd5465;
      68821:data<=16'd4845;
      68822:data<=16'd5151;
      68823:data<=16'd6451;
      68824:data<=16'd6965;
      68825:data<=16'd6437;
      68826:data<=16'd6125;
      68827:data<=16'd5879;
      68828:data<=16'd5671;
      68829:data<=16'd6649;
      68830:data<=16'd7436;
      68831:data<=16'd6643;
      68832:data<=16'd6235;
      68833:data<=16'd6593;
      68834:data<=16'd6155;
      68835:data<=16'd6196;
      68836:data<=16'd7313;
      68837:data<=16'd7078;
      68838:data<=16'd6294;
      68839:data<=16'd6458;
      68840:data<=16'd5604;
      68841:data<=16'd5539;
      68842:data<=16'd7285;
      68843:data<=16'd6799;
      68844:data<=16'd7257;
      68845:data<=16'd11215;
      68846:data<=16'd12269;
      68847:data<=16'd11511;
      68848:data<=16'd12781;
      68849:data<=16'd12651;
      68850:data<=16'd11643;
      68851:data<=16'd11220;
      68852:data<=16'd9993;
      68853:data<=16'd9687;
      68854:data<=16'd9629;
      68855:data<=16'd8466;
      68856:data<=16'd8062;
      68857:data<=16'd7527;
      68858:data<=16'd6614;
      68859:data<=16'd6517;
      68860:data<=16'd5336;
      68861:data<=16'd3439;
      68862:data<=16'd2919;
      68863:data<=16'd2640;
      68864:data<=16'd2109;
      68865:data<=16'd2074;
      68866:data<=16'd1253;
      68867:data<=-16'd523;
      68868:data<=-16'd1095;
      68869:data<=-16'd1113;
      68870:data<=-16'd1773;
      68871:data<=-16'd1506;
      68872:data<=-16'd1797;
      68873:data<=-16'd3697;
      68874:data<=-16'd4082;
      68875:data<=-16'd4053;
      68876:data<=-16'd4523;
      68877:data<=-16'd3662;
      68878:data<=-16'd5858;
      68879:data<=-16'd11415;
      68880:data<=-16'd13036;
      68881:data<=-16'd11855;
      68882:data<=-16'd12289;
      68883:data<=-16'd12342;
      68884:data<=-16'd11497;
      68885:data<=-16'd11847;
      68886:data<=-16'd12795;
      68887:data<=-16'd12815;
      68888:data<=-16'd12492;
      68889:data<=-16'd12278;
      68890:data<=-16'd11386;
      68891:data<=-16'd11294;
      68892:data<=-16'd12713;
      68893:data<=-16'd13001;
      68894:data<=-16'd12301;
      68895:data<=-16'd12117;
      68896:data<=-16'd11620;
      68897:data<=-16'd11526;
      68898:data<=-16'd12624;
      68899:data<=-16'd13063;
      68900:data<=-16'd12284;
      68901:data<=-16'd11894;
      68902:data<=-16'd11858;
      68903:data<=-16'd11317;
      68904:data<=-16'd11843;
      68905:data<=-16'd13085;
      68906:data<=-16'd12777;
      68907:data<=-16'd12590;
      68908:data<=-16'd12330;
      68909:data<=-16'd10910;
      68910:data<=-16'd11913;
      68911:data<=-16'd12182;
      68912:data<=-16'd7708;
      68913:data<=-16'd5422;
      68914:data<=-16'd6102;
      68915:data<=-16'd4980;
      68916:data<=-16'd5333;
      68917:data<=-16'd7080;
      68918:data<=-16'd6895;
      68919:data<=-16'd6751;
      68920:data<=-16'd6695;
      68921:data<=-16'd5985;
      68922:data<=-16'd6291;
      68923:data<=-16'd7297;
      68924:data<=-16'd7926;
      68925:data<=-16'd7739;
      68926:data<=-16'd7250;
      68927:data<=-16'd7180;
      68928:data<=-16'd6874;
      68929:data<=-16'd7209;
      68930:data<=-16'd8379;
      68931:data<=-16'd8247;
      68932:data<=-16'd7597;
      68933:data<=-16'd7363;
      68934:data<=-16'd6619;
      68935:data<=-16'd6849;
      68936:data<=-16'd8470;
      68937:data<=-16'd8824;
      68938:data<=-16'd7688;
      68939:data<=-16'd7150;
      68940:data<=-16'd7042;
      68941:data<=-16'd6940;
      68942:data<=-16'd8214;
      68943:data<=-16'd8684;
      68944:data<=-16'd7101;
      68945:data<=-16'd8943;
      68946:data<=-16'd13183;
      68947:data<=-16'd13546;
      68948:data<=-16'd12983;
      68949:data<=-16'd13853;
      68950:data<=-16'd13267;
      68951:data<=-16'd12425;
      68952:data<=-16'd11897;
      68953:data<=-16'd10907;
      68954:data<=-16'd10586;
      68955:data<=-16'd10143;
      68956:data<=-16'd9438;
      68957:data<=-16'd8849;
      68958:data<=-16'd7859;
      68959:data<=-16'd7674;
      68960:data<=-16'd6977;
      68961:data<=-16'd4813;
      68962:data<=-16'd4208;
      68963:data<=-16'd4128;
      68964:data<=-16'd3136;
      68965:data<=-16'd3262;
      68966:data<=-16'd2723;
      68967:data<=-16'd610;
      68968:data<=16'd111;
      68969:data<=16'd67;
      68970:data<=16'd752;
      68971:data<=16'd770;
      68972:data<=16'd635;
      68973:data<=16'd1891;
      68974:data<=16'd3019;
      68975:data<=16'd3230;
      68976:data<=16'd3557;
      68977:data<=16'd3110;
      68978:data<=16'd3918;
      68979:data<=16'd8781;
      68980:data<=16'd12239;
      68981:data<=16'd11556;
      68982:data<=16'd11520;
      68983:data<=16'd11492;
      68984:data<=16'd10234;
      68985:data<=16'd10815;
      68986:data<=16'd12176;
      68987:data<=16'd12313;
      68988:data<=16'd11888;
      68989:data<=16'd11194;
      68990:data<=16'd10869;
      68991:data<=16'd11142;
      68992:data<=16'd11776;
      68993:data<=16'd12240;
      68994:data<=16'd11708;
      68995:data<=16'd11388;
      68996:data<=16'd11415;
      68997:data<=16'd10771;
      68998:data<=16'd11176;
      68999:data<=16'd12196;
      69000:data<=16'd11828;
      69001:data<=16'd11568;
      69002:data<=16'd11438;
      69003:data<=16'd10295;
      69004:data<=16'd10618;
      69005:data<=16'd12578;
      69006:data<=16'd12659;
      69007:data<=16'd11753;
      69008:data<=16'd11805;
      69009:data<=16'd10871;
      69010:data<=16'd10843;
      69011:data<=16'd12743;
      69012:data<=16'd10310;
      69013:data<=16'd5318;
      69014:data<=16'd4752;
      69015:data<=16'd5307;
      69016:data<=16'd4857;
      69017:data<=16'd6028;
      69018:data<=16'd6672;
      69019:data<=16'd6231;
      69020:data<=16'd6364;
      69021:data<=16'd6161;
      69022:data<=16'd5809;
      69023:data<=16'd6329;
      69024:data<=16'd7532;
      69025:data<=16'd7978;
      69026:data<=16'd7326;
      69027:data<=16'd7109;
      69028:data<=16'd6654;
      69029:data<=16'd6636;
      69030:data<=16'd8451;
      69031:data<=16'd8563;
      69032:data<=16'd7075;
      69033:data<=16'd7051;
      69034:data<=16'd6865;
      69035:data<=16'd7054;
      69036:data<=16'd8448;
      69037:data<=16'd8410;
      69038:data<=16'd7551;
      69039:data<=16'd7368;
      69040:data<=16'd7113;
      69041:data<=16'd6839;
      69042:data<=16'd7547;
      69043:data<=16'd8351;
      69044:data<=16'd7285;
      69045:data<=16'd8025;
      69046:data<=16'd12289;
      69047:data<=16'd13430;
      69048:data<=16'd12451;
      69049:data<=16'd13878;
      69050:data<=16'd13668;
      69051:data<=16'd12026;
      69052:data<=16'd11802;
      69053:data<=16'd11226;
      69054:data<=16'd10733;
      69055:data<=16'd10232;
      69056:data<=16'd9298;
      69057:data<=16'd8989;
      69058:data<=16'd8176;
      69059:data<=16'd7538;
      69060:data<=16'd7012;
      69061:data<=16'd5016;
      69062:data<=16'd4077;
      69063:data<=16'd4100;
      69064:data<=16'd3231;
      69065:data<=16'd3058;
      69066:data<=16'd2942;
      69067:data<=16'd1754;
      69068:data<=16'd476;
      69069:data<=-16'd230;
      69070:data<=-16'd411;
      69071:data<=-16'd675;
      69072:data<=-16'd262;
      69073:data<=-16'd593;
      69074:data<=-16'd3037;
      69075:data<=-16'd3503;
      69076:data<=-16'd2805;
      69077:data<=-16'd3204;
      69078:data<=-16'd2547;
      69079:data<=-16'd5544;
      69080:data<=-16'd11562;
      69081:data<=-16'd12066;
      69082:data<=-16'd10715;
      69083:data<=-16'd11059;
      69084:data<=-16'd10053;
      69085:data<=-16'd10354;
      69086:data<=-16'd11885;
      69087:data<=-16'd11790;
      69088:data<=-16'd11358;
      69089:data<=-16'd11074;
      69090:data<=-16'd10853;
      69091:data<=-16'd10395;
      69092:data<=-16'd10307;
      69093:data<=-16'd11470;
      69094:data<=-16'd11485;
      69095:data<=-16'd11033;
      69096:data<=-16'd11215;
      69097:data<=-16'd9917;
      69098:data<=-16'd10058;
      69099:data<=-16'd12110;
      69100:data<=-16'd11805;
      69101:data<=-16'd10998;
      69102:data<=-16'd10895;
      69103:data<=-16'd9818;
      69104:data<=-16'd10014;
      69105:data<=-16'd11784;
      69106:data<=-16'd12017;
      69107:data<=-16'd10963;
      69108:data<=-16'd10807;
      69109:data<=-16'd10461;
      69110:data<=-16'd9978;
      69111:data<=-16'd11615;
      69112:data<=-16'd10745;
      69113:data<=-16'd5560;
      69114:data<=-16'd3968;
      69115:data<=-16'd4957;
      69116:data<=-16'd3677;
      69117:data<=-16'd4187;
      69118:data<=-16'd5915;
      69119:data<=-16'd5645;
      69120:data<=-16'd5536;
      69121:data<=-16'd5221;
      69122:data<=-16'd4390;
      69123:data<=-16'd5224;
      69124:data<=-16'd6655;
      69125:data<=-16'd6751;
      69126:data<=-16'd6175;
      69127:data<=-16'd5988;
      69128:data<=-16'd5676;
      69129:data<=-16'd5789;
      69130:data<=-16'd7034;
      69131:data<=-16'd7000;
      69132:data<=-16'd6038;
      69133:data<=-16'd6172;
      69134:data<=-16'd5712;
      69135:data<=-16'd5371;
      69136:data<=-16'd6428;
      69137:data<=-16'd6933;
      69138:data<=-16'd6746;
      69139:data<=-16'd6229;
      69140:data<=-16'd5695;
      69141:data<=-16'd5679;
      69142:data<=-16'd5873;
      69143:data<=-16'd6910;
      69144:data<=-16'd6769;
      69145:data<=-16'd5695;
      69146:data<=-16'd8704;
      69147:data<=-16'd12129;
      69148:data<=-16'd11838;
      69149:data<=-16'd12264;
      69150:data<=-16'd12686;
      69151:data<=-16'd11353;
      69152:data<=-16'd10941;
      69153:data<=-16'd10586;
      69154:data<=-16'd9824;
      69155:data<=-16'd9241;
      69156:data<=-16'd8352;
      69157:data<=-16'd8156;
      69158:data<=-16'd7655;
      69159:data<=-16'd6595;
      69160:data<=-16'd6391;
      69161:data<=-16'd5163;
      69162:data<=-16'd3262;
      69163:data<=-16'd2787;
      69164:data<=-16'd2285;
      69165:data<=-16'd1883;
      69166:data<=-16'd2416;
      69167:data<=-16'd1506;
      69168:data<=16'd705;
      69169:data<=16'd1152;
      69170:data<=16'd872;
      69171:data<=16'd1469;
      69172:data<=16'd1048;
      69173:data<=16'd1568;
      69174:data<=16'd4132;
      69175:data<=16'd4144;
      69176:data<=16'd3542;
      69177:data<=16'd4350;
      69178:data<=16'd3090;
      69179:data<=16'd4989;
      69180:data<=16'd11465;
      69181:data<=16'd13209;
      69182:data<=16'd11603;
      69183:data<=16'd11944;
      69184:data<=16'd11705;
      69185:data<=16'd10983;
      69186:data<=16'd11582;
      69187:data<=16'd12584;
      69188:data<=16'd12795;
      69189:data<=16'd12178;
      69190:data<=16'd11829;
      69191:data<=16'd11218;
      69192:data<=16'd11160;
      69193:data<=16'd12772;
      69194:data<=16'd12833;
      69195:data<=16'd11752;
      69196:data<=16'd11781;
      69197:data<=16'd11121;
      69198:data<=16'd11294;
      69199:data<=16'd12883;
      69200:data<=16'd12665;
      69201:data<=16'd11799;
      69202:data<=16'd11618;
      69203:data<=16'd11229;
      69204:data<=16'd11291;
      69205:data<=16'd12008;
      69206:data<=16'd12680;
      69207:data<=16'd12469;
      69208:data<=16'd11991;
      69209:data<=16'd11740;
      69210:data<=16'd10698;
      69211:data<=16'd11297;
      69212:data<=16'd12505;
      69213:data<=16'd8931;
      69214:data<=16'd5018;
      69215:data<=16'd5045;
      69216:data<=16'd4849;
      69217:data<=16'd5172;
      69218:data<=16'd6816;
      69219:data<=16'd6502;
      69220:data<=16'd5765;
      69221:data<=16'd5885;
      69222:data<=16'd5702;
      69223:data<=16'd6075;
      69224:data<=16'd6815;
      69225:data<=16'd6910;
      69226:data<=16'd6637;
      69227:data<=16'd6511;
      69228:data<=16'd6299;
      69229:data<=16'd5805;
      69230:data<=16'd6488;
      69231:data<=16'd7700;
      69232:data<=16'd7021;
      69233:data<=16'd6050;
      69234:data<=16'd6072;
      69235:data<=16'd5770;
      69236:data<=16'd6037;
      69237:data<=16'd7080;
      69238:data<=16'd6925;
      69239:data<=16'd5985;
      69240:data<=16'd6003;
      69241:data<=16'd6041;
      69242:data<=16'd5429;
      69243:data<=16'd6290;
      69244:data<=16'd6886;
      69245:data<=16'd5137;
      69246:data<=16'd6655;
      69247:data<=16'd11361;
      69248:data<=16'd12208;
      69249:data<=16'd11518;
      69250:data<=16'd12377;
      69251:data<=16'd11764;
      69252:data<=16'd10730;
      69253:data<=16'd10404;
      69254:data<=16'd9715;
      69255:data<=16'd9391;
      69256:data<=16'd8758;
      69257:data<=16'd7929;
      69258:data<=16'd7665;
      69259:data<=16'd6980;
      69260:data<=16'd6528;
      69261:data<=16'd5535;
      69262:data<=16'd3254;
      69263:data<=16'd2573;
      69264:data<=16'd2643;
      69265:data<=16'd1914;
      69266:data<=16'd2140;
      69267:data<=16'd1463;
      69268:data<=-16'd717;
      69269:data<=-16'd1240;
      69270:data<=-16'd969;
      69271:data<=-16'd1347;
      69272:data<=-16'd1474;
      69273:data<=-16'd2059;
      69274:data<=-16'd3438;
      69275:data<=-16'd4153;
      69276:data<=-16'd4100;
      69277:data<=-16'd4356;
      69278:data<=-16'd4144;
      69279:data<=-16'd4099;
      69280:data<=-16'd7965;
      69281:data<=-16'd12815;
      69282:data<=-16'd12760;
      69283:data<=-16'd11555;
      69284:data<=-16'd12022;
      69285:data<=-16'd11112;
      69286:data<=-16'd11221;
      69287:data<=-16'd13247;
      69288:data<=-16'd12977;
      69289:data<=-16'd11899;
      69290:data<=-16'd12128;
      69291:data<=-16'd11872;
      69292:data<=-16'd12110;
      69293:data<=-16'd13224;
      69294:data<=-16'd12928;
      69295:data<=-16'd12119;
      69296:data<=-16'd12263;
      69297:data<=-16'd12044;
      69298:data<=-16'd11615;
      69299:data<=-16'd12464;
      69300:data<=-16'd13405;
      69301:data<=-16'd12900;
      69302:data<=-16'd12257;
      69303:data<=-16'd12132;
      69304:data<=-16'd11414;
      69305:data<=-16'd11650;
      69306:data<=-16'd13591;
      69307:data<=-16'd13462;
      69308:data<=-16'd11972;
      69309:data<=-16'd12489;
      69310:data<=-16'd12019;
      69311:data<=-16'd11458;
      69312:data<=-16'd13756;
      69313:data<=-16'd11914;
      69314:data<=-16'd6123;
      69315:data<=-16'd5292;
      69316:data<=-16'd6304;
      69317:data<=-16'd5636;
      69318:data<=-16'd6789;
      69319:data<=-16'd7442;
      69320:data<=-16'd6584;
      69321:data<=-16'd6758;
      69322:data<=-16'd6492;
      69323:data<=-16'd6078;
      69324:data<=-16'd6910;
      69325:data<=-16'd7562;
      69326:data<=-16'd7436;
      69327:data<=-16'd7087;
      69328:data<=-16'd7021;
      69329:data<=-16'd6754;
      69330:data<=-16'd6599;
      69331:data<=-16'd7677;
      69332:data<=-16'd7958;
      69333:data<=-16'd7162;
      69334:data<=-16'd7074;
      69335:data<=-16'd6391;
      69336:data<=-16'd6159;
      69337:data<=-16'd7335;
      69338:data<=-16'd7239;
      69339:data<=-16'd6611;
      69340:data<=-16'd6393;
      69341:data<=-16'd5688;
      69342:data<=-16'd5767;
      69343:data<=-16'd6660;
      69344:data<=-16'd6957;
      69345:data<=-16'd6132;
      69346:data<=-16'd6317;
      69347:data<=-16'd9820;
      69348:data<=-16'd12396;
      69349:data<=-16'd11994;
      69350:data<=-16'd12446;
      69351:data<=-16'd12569;
      69352:data<=-16'd11359;
      69353:data<=-16'd11000;
      69354:data<=-16'd10519;
      69355:data<=-16'd9665;
      69356:data<=-16'd8880;
      69357:data<=-16'd8293;
      69358:data<=-16'd8395;
      69359:data<=-16'd7712;
      69360:data<=-16'd6977;
      69361:data<=-16'd6385;
      69362:data<=-16'd4096;
      69363:data<=-16'd3071;
      69364:data<=-16'd3466;
      69365:data<=-16'd2399;
      69366:data<=-16'd2106;
      69367:data<=-16'd2109;
      69368:data<=-16'd464;
      69369:data<=16'd610;
      69370:data<=16'd638;
      69371:data<=16'd734;
      69372:data<=16'd961;
      69373:data<=16'd728;
      69374:data<=16'd1204;
      69375:data<=16'd3377;
      69376:data<=16'd3507;
      69377:data<=16'd2726;
      69378:data<=16'd3791;
      69379:data<=16'd2772;
      69380:data<=16'd4466;
      69381:data<=16'd11400;
      69382:data<=16'd12680;
      69383:data<=16'd10507;
      69384:data<=16'd11433;
      69385:data<=16'd10818;
      69386:data<=16'd10575;
      69387:data<=16'd12289;
      69388:data<=16'd12025;
      69389:data<=16'd11715;
      69390:data<=16'd11734;
      69391:data<=16'd11060;
      69392:data<=16'd11223;
      69393:data<=16'd11729;
      69394:data<=16'd12289;
      69395:data<=16'd11843;
      69396:data<=16'd10863;
      69397:data<=16'd11339;
      69398:data<=16'd10783;
      69399:data<=16'd10410;
      69400:data<=16'd12317;
      69401:data<=16'd12084;
      69402:data<=16'd10833;
      69403:data<=16'd11321;
      69404:data<=16'd10796;
      69405:data<=16'd10745;
      69406:data<=16'd12360;
      69407:data<=16'd12354;
      69408:data<=16'd11414;
      69409:data<=16'd11492;
      69410:data<=16'd11129;
      69411:data<=16'd10693;
      69412:data<=16'd12076;
      69413:data<=16'd11787;
      69414:data<=16'd7391;
      69415:data<=16'd4429;
      69416:data<=16'd4613;
      69417:data<=16'd4566;
      69418:data<=16'd5125;
      69419:data<=16'd6097;
      69420:data<=16'd5783;
      69421:data<=16'd5353;
      69422:data<=16'd5172;
      69423:data<=16'd5065;
      69424:data<=16'd5294;
      69425:data<=16'd5791;
      69426:data<=16'd6203;
      69427:data<=16'd5962;
      69428:data<=16'd5971;
      69429:data<=16'd5943;
      69430:data<=16'd5524;
      69431:data<=16'd6523;
      69432:data<=16'd7154;
      69433:data<=16'd6560;
      69434:data<=16'd6610;
      69435:data<=16'd5774;
      69436:data<=16'd5506;
      69437:data<=16'd6890;
      69438:data<=16'd6598;
      69439:data<=16'd6041;
      69440:data<=16'd5917;
      69441:data<=16'd5271;
      69442:data<=16'd5768;
      69443:data<=16'd5712;
      69444:data<=16'd5833;
      69445:data<=16'd6724;
      69446:data<=16'd5310;
      69447:data<=16'd6649;
      69448:data<=16'd11288;
      69449:data<=16'd12003;
      69450:data<=16'd11764;
      69451:data<=16'd12604;
      69452:data<=16'd11685;
      69453:data<=16'd11022;
      69454:data<=16'd10493;
      69455:data<=16'd9693;
      69456:data<=16'd9518;
      69457:data<=16'd8836;
      69458:data<=16'd8564;
      69459:data<=16'd8093;
      69460:data<=16'd7003;
      69461:data<=16'd6783;
      69462:data<=16'd5125;
      69463:data<=16'd3306;
      69464:data<=16'd3767;
      69465:data<=16'd3054;
      69466:data<=16'd1962;
      69467:data<=16'd2487;
      69468:data<=16'd1610;
      69469:data<=-16'd224;
      69470:data<=-16'd294;
      69471:data<=16'd193;
      69472:data<=-16'd519;
      69473:data<=-16'd840;
      69474:data<=-16'd834;
      69475:data<=-16'd2549;
      69476:data<=-16'd3104;
      69477:data<=-16'd2294;
      69478:data<=-16'd3099;
      69479:data<=-16'd2578;
      69480:data<=-16'd3265;
      69481:data<=-16'd8789;
      69482:data<=-16'd11643;
      69483:data<=-16'd10696;
      69484:data<=-16'd10840;
      69485:data<=-16'd10548;
      69486:data<=-16'd10222;
      69487:data<=-16'd11188;
      69488:data<=-16'd11882;
      69489:data<=-16'd11564;
      69490:data<=-16'd10636;
      69491:data<=-16'd10760;
      69492:data<=-16'd10815;
      69493:data<=-16'd10445;
      69494:data<=-16'd11887;
      69495:data<=-16'd11844;
      69496:data<=-16'd10443;
      69497:data<=-16'd11136;
      69498:data<=-16'd10605;
      69499:data<=-16'd10125;
      69500:data<=-16'd11746;
      69501:data<=-16'd11464;
      69502:data<=-16'd10972;
      69503:data<=-16'd11192;
      69504:data<=-16'd10161;
      69505:data<=-16'd10404;
      69506:data<=-16'd11617;
      69507:data<=-16'd12145;
      69508:data<=-16'd11826;
      69509:data<=-16'd10780;
      69510:data<=-16'd11041;
      69511:data<=-16'd10907;
      69512:data<=-16'd10668;
      69513:data<=-16'd12511;
      69514:data<=-16'd10164;
      69515:data<=-16'd4833;
      69516:data<=-16'd4182;
      69517:data<=-16'd4473;
      69518:data<=-16'd4176;
      69519:data<=-16'd5601;
      69520:data<=-16'd5721;
      69521:data<=-16'd5470;
      69522:data<=-16'd5799;
      69523:data<=-16'd4916;
      69524:data<=-16'd5169;
      69525:data<=-16'd6560;
      69526:data<=-16'd6613;
      69527:data<=-16'd6070;
      69528:data<=-16'd5706;
      69529:data<=-16'd5453;
      69530:data<=-16'd5651;
      69531:data<=-16'd6478;
      69532:data<=-16'd6931;
      69533:data<=-16'd6338;
      69534:data<=-16'd6015;
      69535:data<=-16'd5911;
      69536:data<=-16'd5442;
      69537:data<=-16'd5606;
      69538:data<=-16'd6182;
      69539:data<=-16'd6608;
      69540:data<=-16'd6429;
      69541:data<=-16'd5498;
      69542:data<=-16'd5059;
      69543:data<=-16'd5216;
      69544:data<=-16'd6049;
      69545:data<=-16'd6757;
      69546:data<=-16'd5607;
      69547:data<=-16'd5915;
      69548:data<=-16'd9197;
      69549:data<=-16'd11398;
      69550:data<=-16'd12145;
      69551:data<=-16'd12132;
      69552:data<=-16'd11232;
      69553:data<=-16'd10733;
      69554:data<=-16'd9876;
      69555:data<=-16'd9203;
      69556:data<=-16'd9179;
      69557:data<=-16'd7993;
      69558:data<=-16'd7571;
      69559:data<=-16'd7809;
      69560:data<=-16'd6484;
      69561:data<=-16'd6070;
      69562:data<=-16'd5611;
      69563:data<=-16'd3462;
      69564:data<=-16'd3022;
      69565:data<=-16'd3140;
      69566:data<=-16'd1798;
      69567:data<=-16'd1330;
      69568:data<=-16'd1021;
      69569:data<=16'd343;
      69570:data<=16'd945;
      69571:data<=16'd805;
      69572:data<=16'd1312;
      69573:data<=16'd1765;
      69574:data<=16'd1823;
      69575:data<=16'd3157;
      69576:data<=16'd4379;
      69577:data<=16'd3573;
      69578:data<=16'd3739;
      69579:data<=16'd4350;
      69580:data<=16'd3344;
      69581:data<=16'd6134;
      69582:data<=16'd11923;
      69583:data<=16'd12665;
      69584:data<=16'd11012;
      69585:data<=16'd11649;
      69586:data<=16'd11442;
      69587:data<=16'd11091;
      69588:data<=16'd12471;
      69589:data<=16'd12480;
      69590:data<=16'd11699;
      69591:data<=16'd11890;
      69592:data<=16'd11270;
      69593:data<=16'd11285;
      69594:data<=16'd12877;
      69595:data<=16'd12971;
      69596:data<=16'd12193;
      69597:data<=16'd12041;
      69598:data<=16'd11421;
      69599:data<=16'd11435;
      69600:data<=16'd12475;
      69601:data<=16'd12815;
      69602:data<=16'd12284;
      69603:data<=16'd11552;
      69604:data<=16'd11391;
      69605:data<=16'd11524;
      69606:data<=16'd11705;
      69607:data<=16'd12674;
      69608:data<=16'd12713;
      69609:data<=16'd11855;
      69610:data<=16'd12087;
      69611:data<=16'd11439;
      69612:data<=16'd11198;
      69613:data<=16'd13113;
      69614:data<=16'd11726;
      69615:data<=16'd7482;
      69616:data<=16'd5700;
      69617:data<=16'd5228;
      69618:data<=16'd5482;
      69619:data<=16'd6689;
      69620:data<=16'd6940;
      69621:data<=16'd6887;
      69622:data<=16'd6586;
      69623:data<=16'd5990;
      69624:data<=16'd6637;
      69625:data<=16'd7280;
      69626:data<=16'd7154;
      69627:data<=16'd6995;
      69628:data<=16'd6564;
      69629:data<=16'd6402;
      69630:data<=16'd6302;
      69631:data<=16'd6446;
      69632:data<=16'd7450;
      69633:data<=16'd7571;
      69634:data<=16'd7183;
      69635:data<=16'd6986;
      69636:data<=16'd5870;
      69637:data<=16'd6123;
      69638:data<=16'd7697;
      69639:data<=16'd7653;
      69640:data<=16'd7191;
      69641:data<=16'd6531;
      69642:data<=16'd5759;
      69643:data<=16'd6681;
      69644:data<=16'd7297;
      69645:data<=16'd7168;
      69646:data<=16'd7090;
      69647:data<=16'd5623;
      69648:data<=16'd6583;
      69649:data<=16'd11361;
      69650:data<=16'd13267;
      69651:data<=16'd12148;
      69652:data<=16'd12270;
      69653:data<=16'd12013;
      69654:data<=16'd10419;
      69655:data<=16'd9685;
      69656:data<=16'd9515;
      69657:data<=16'd8718;
      69658:data<=16'd8301;
      69659:data<=16'd8172;
      69660:data<=16'd7171;
      69661:data<=16'd6579;
      69662:data<=16'd6073;
      69663:data<=16'd4190;
      69664:data<=16'd3289;
      69665:data<=16'd3480;
      69666:data<=16'd2711;
      69667:data<=16'd2334;
      69668:data<=16'd1838;
      69669:data<=16'd83;
      69670:data<=-16'd652;
      69671:data<=-16'd232;
      69672:data<=-16'd491;
      69673:data<=-16'd1324;
      69674:data<=-16'd1861;
      69675:data<=-16'd2535;
      69676:data<=-16'd3692;
      69677:data<=-16'd3644;
      69678:data<=-16'd3368;
      69679:data<=-16'd4211;
      69680:data<=-16'd3574;
      69681:data<=-16'd4717;
      69682:data<=-16'd10208;
      69683:data<=-16'd12505;
      69684:data<=-16'd11223;
      69685:data<=-16'd11358;
      69686:data<=-16'd11060;
      69687:data<=-16'd11220;
      69688:data<=-16'd12671;
      69689:data<=-16'd12422;
      69690:data<=-16'd11862;
      69691:data<=-16'd11549;
      69692:data<=-16'd10774;
      69693:data<=-16'd11436;
      69694:data<=-16'd12669;
      69695:data<=-16'd12985;
      69696:data<=-16'd12484;
      69697:data<=-16'd11702;
      69698:data<=-16'd11829;
      69699:data<=-16'd11970;
      69700:data<=-16'd12170;
      69701:data<=-16'd13026;
      69702:data<=-16'd12727;
      69703:data<=-16'd12352;
      69704:data<=-16'd12254;
      69705:data<=-16'd11145;
      69706:data<=-16'd11664;
      69707:data<=-16'd13038;
      69708:data<=-16'd12725;
      69709:data<=-16'd12449;
      69710:data<=-16'd12081;
      69711:data<=-16'd11515;
      69712:data<=-16'd11728;
      69713:data<=-16'd12457;
      69714:data<=-16'd13691;
      69715:data<=-16'd11424;
      69716:data<=-16'd5773;
      69717:data<=-16'd4716;
      69718:data<=-16'd6772;
      69719:data<=-16'd6846;
      69720:data<=-16'd7344;
      69721:data<=-16'd7679;
      69722:data<=-16'd6933;
      69723:data<=-16'd6968;
      69724:data<=-16'd6581;
      69725:data<=-16'd6780;
      69726:data<=-16'd8348;
      69727:data<=-16'd8308;
      69728:data<=-16'd7582;
      69729:data<=-16'd7389;
      69730:data<=-16'd6569;
      69731:data<=-16'd7004;
      69732:data<=-16'd8472;
      69733:data<=-16'd8150;
      69734:data<=-16'd7448;
      69735:data<=-16'd7386;
      69736:data<=-16'd6883;
      69737:data<=-16'd7385;
      69738:data<=-16'd8595;
      69739:data<=-16'd8392;
      69740:data<=-16'd7964;
      69741:data<=-16'd7871;
      69742:data<=-16'd7374;
      69743:data<=-16'd7359;
      69744:data<=-16'd7726;
      69745:data<=-16'd8285;
      69746:data<=-16'd8478;
      69747:data<=-16'd7227;
      69748:data<=-16'd7733;
      69749:data<=-16'd11335;
      69750:data<=-16'd13696;
      69751:data<=-16'd13937;
      69752:data<=-16'd13755;
      69753:data<=-16'd13144;
      69754:data<=-16'd12340;
      69755:data<=-16'd11403;
      69756:data<=-16'd10815;
      69757:data<=-16'd10548;
      69758:data<=-16'd9735;
      69759:data<=-16'd9147;
      69760:data<=-16'd8740;
      69761:data<=-16'd8156;
      69762:data<=-16'd7589;
      69763:data<=-16'd5867;
      69764:data<=-16'd4404;
      69765:data<=-16'd4444;
      69766:data<=-16'd3971;
      69767:data<=-16'd3635;
      69768:data<=-16'd3533;
      69769:data<=-16'd2088;
      69770:data<=-16'd993;
      69771:data<=-16'd773;
      69772:data<=-16'd481;
      69773:data<=-16'd334;
      69774:data<=-16'd18;
      69775:data<=16'd557;
      69776:data<=16'd1820;
      69777:data<=16'd2717;
      69778:data<=16'd2112;
      69779:data<=16'd2500;
      69780:data<=16'd2717;
      69781:data<=16'd2071;
      69782:data<=16'd5824;
      69783:data<=16'd10869;
      69784:data<=16'd11079;
      69785:data<=16'd10046;
      69786:data<=16'd10117;
      69787:data<=16'd10331;
      69788:data<=16'd11224;
      69789:data<=16'd11624;
      69790:data<=16'd11230;
      69791:data<=16'd10824;
      69792:data<=16'd10182;
      69793:data<=16'd9973;
      69794:data<=16'd10563;
      69795:data<=16'd11323;
      69796:data<=16'd11430;
      69797:data<=16'd10968;
      69798:data<=16'd10554;
      69799:data<=16'd9878;
      69800:data<=16'd10261;
      69801:data<=16'd11731;
      69802:data<=16'd11535;
      69803:data<=16'd11092;
      69804:data<=16'd11274;
      69805:data<=16'd10339;
      69806:data<=16'd10731;
      69807:data<=16'd12367;
      69808:data<=16'd12143;
      69809:data<=16'd11371;
      69810:data<=16'd11130;
      69811:data<=16'd10927;
      69812:data<=16'd10819;
      69813:data<=16'd11195;
      69814:data<=16'd12192;
      69815:data<=16'd10334;
      69816:data<=16'd5726;
      69817:data<=16'd4082;
      69818:data<=16'd4582;
      69819:data<=16'd4843;
      69820:data<=16'd5920;
      69821:data<=16'd5911;
      69822:data<=16'd5316;
      69823:data<=16'd5642;
      69824:data<=16'd5034;
      69825:data<=16'd5306;
      69826:data<=16'd6921;
      69827:data<=16'd6602;
      69828:data<=16'd5803;
      69829:data<=16'd5796;
      69830:data<=16'd5357;
      69831:data<=16'd5806;
      69832:data<=16'd6901;
      69833:data<=16'd6605;
      69834:data<=16'd5888;
      69835:data<=16'd6026;
      69836:data<=16'd5861;
      69837:data<=16'd5468;
      69838:data<=16'd6408;
      69839:data<=16'd7053;
      69840:data<=16'd6220;
      69841:data<=16'd6188;
      69842:data<=16'd6141;
      69843:data<=16'd5209;
      69844:data<=16'd5871;
      69845:data<=16'd6884;
      69846:data<=16'd6734;
      69847:data<=16'd6554;
      69848:data<=16'd5824;
      69849:data<=16'd7232;
      69850:data<=16'd11956;
      69851:data<=16'd13579;
      69852:data<=16'd11853;
      69853:data<=16'd11828;
      69854:data<=16'd11790;
      69855:data<=16'd10586;
      69856:data<=16'd10108;
      69857:data<=16'd9459;
      69858:data<=16'd8742;
      69859:data<=16'd8592;
      69860:data<=16'd7918;
      69861:data<=16'd7316;
      69862:data<=16'd6957;
      69863:data<=16'd5557;
      69864:data<=16'd4020;
      69865:data<=16'd3506;
      69866:data<=16'd3128;
      69867:data<=16'd2637;
      69868:data<=16'd2736;
      69869:data<=16'd2234;
      69870:data<=16'd364;
      69871:data<=-16'd541;
      69872:data<=-16'd287;
      69873:data<=-16'd763;
      69874:data<=-16'd852;
      69875:data<=-16'd998;
      69876:data<=-16'd2907;
      69877:data<=-16'd3745;
      69878:data<=-16'd2931;
      69879:data<=-16'd3366;
      69880:data<=-16'd3571;
      69881:data<=-16'd3172;
      69882:data<=-16'd5999;
      69883:data<=-16'd10730;
      69884:data<=-16'd12392;
      69885:data<=-16'd11447;
      69886:data<=-16'd11027;
      69887:data<=-16'd11133;
      69888:data<=-16'd11453;
      69889:data<=-16'd12278;
      69890:data<=-16'd12190;
      69891:data<=-16'd11356;
      69892:data<=-16'd11000;
      69893:data<=-16'd10510;
      69894:data<=-16'd11147;
      69895:data<=-16'd12986;
      69896:data<=-16'd12736;
      69897:data<=-16'd11721;
      69898:data<=-16'd11773;
      69899:data<=-16'd10894;
      69900:data<=-16'd10936;
      69901:data<=-16'd12560;
      69902:data<=-16'd12236;
      69903:data<=-16'd11461;
      69904:data<=-16'd11574;
      69905:data<=-16'd10749;
      69906:data<=-16'd10912;
      69907:data<=-16'd11693;
      69908:data<=-16'd10434;
      69909:data<=-16'd9668;
      69910:data<=-16'd10035;
      69911:data<=-16'd9294;
      69912:data<=-16'd8766;
      69913:data<=-16'd9235;
      69914:data<=-16'd10040;
      69915:data<=-16'd10369;
      69916:data<=-16'd8031;
      69917:data<=-16'd4698;
      69918:data<=-16'd4184;
      69919:data<=-16'd5532;
      69920:data<=-16'd6590;
      69921:data<=-16'd6819;
      69922:data<=-16'd6193;
      69923:data<=-16'd5600;
      69924:data<=-16'd5371;
      69925:data<=-16'd5776;
      69926:data<=-16'd6916;
      69927:data<=-16'd7168;
      69928:data<=-16'd6426;
      69929:data<=-16'd6015;
      69930:data<=-16'd5750;
      69931:data<=-16'd5700;
      69932:data<=-16'd6354;
      69933:data<=-16'd7006;
      69934:data<=-16'd6783;
      69935:data<=-16'd6109;
      69936:data<=-16'd5685;
      69937:data<=-16'd5319;
      69938:data<=-16'd5846;
      69939:data<=-16'd7130;
      69940:data<=-16'd6858;
      69941:data<=-16'd6097;
      69942:data<=-16'd6102;
      69943:data<=-16'd5421;
      69944:data<=-16'd5685;
      69945:data<=-16'd6977;
      69946:data<=-16'd6816;
      69947:data<=-16'd6463;
      69948:data<=-16'd6120;
      69949:data<=-16'd6291;
      69950:data<=-16'd9253;
      69951:data<=-16'd11345;
      69952:data<=-16'd10469;
      69953:data<=-16'd10046;
      69954:data<=-16'd9753;
      69955:data<=-16'd8766;
      69956:data<=-16'd8254;
      69957:data<=-16'd7718;
      69958:data<=-16'd7319;
      69959:data<=-16'd7171;
      69960:data<=-16'd6575;
      69961:data<=-16'd6147;
      69962:data<=-16'd6147;
      69963:data<=-16'd5251;
      69964:data<=-16'd3177;
      69965:data<=-16'd2218;
      69966:data<=-16'd2511;
      69967:data<=-16'd1988;
      69968:data<=-16'd1741;
      69969:data<=-16'd1281;
      69970:data<=16'd741;
      69971:data<=16'd1387;
      69972:data<=16'd1189;
      69973:data<=16'd1941;
      69974:data<=16'd1845;
      69975:data<=16'd2343;
      69976:data<=16'd3788;
      69977:data<=16'd4196;
      69978:data<=16'd4629;
      69979:data<=16'd4754;
      69980:data<=16'd4538;
      69981:data<=16'd4755;
      69982:data<=16'd5122;
      69983:data<=16'd8146;
      69984:data<=16'd11561;
      69985:data<=16'd10910;
      69986:data<=16'd9947;
      69987:data<=16'd10266;
      69988:data<=16'd10571;
      69989:data<=16'd11876;
      69990:data<=16'd11861;
      69991:data<=16'd10919;
      69992:data<=16'd11177;
      69993:data<=16'd10643;
      69994:data<=16'd10859;
      69995:data<=16'd12464;
      69996:data<=16'd12334;
      69997:data<=16'd11614;
      69998:data<=16'd11415;
      69999:data<=16'd11079;
      70000:data<=16'd11282;
      70001:data<=16'd11914;
      70002:data<=16'd12508;
      70003:data<=16'd12293;
      70004:data<=16'd11655;
      70005:data<=16'd11494;
      70006:data<=16'd10840;
      70007:data<=16'd11218;
      70008:data<=16'd12818;
      70009:data<=16'd12404;
      70010:data<=16'd11602;
      70011:data<=16'd11634;
      70012:data<=16'd10951;
      70013:data<=16'd11339;
      70014:data<=16'd12511;
      70015:data<=16'd12420;
      70016:data<=16'd10884;
      70017:data<=16'd7768;
      70018:data<=16'd5935;
      70019:data<=16'd6960;
      70020:data<=16'd7953;
      70021:data<=16'd8231;
      70022:data<=16'd8113;
      70023:data<=16'd7635;
      70024:data<=16'd7509;
      70025:data<=16'd7186;
      70026:data<=16'd7747;
      70027:data<=16'd9162;
      70028:data<=16'd8526;
      70029:data<=16'd7444;
      70030:data<=16'd7624;
      70031:data<=16'd7021;
      70032:data<=16'd7031;
      70033:data<=16'd8405;
      70034:data<=16'd8122;
      70035:data<=16'd7279;
      70036:data<=16'd7608;
      70037:data<=16'd7063;
      70038:data<=16'd6909;
      70039:data<=16'd8395;
      70040:data<=16'd8175;
      70041:data<=16'd7191;
      70042:data<=16'd7679;
      70043:data<=16'd7065;
      70044:data<=16'd6642;
      70045:data<=16'd8184;
      70046:data<=16'd8401;
      70047:data<=16'd7639;
      70048:data<=16'd7109;
      70049:data<=16'd6302;
      70050:data<=16'd8181;
      70051:data<=16'd11500;
      70052:data<=16'd11731;
      70053:data<=16'd10801;
      70054:data<=16'd10725;
      70055:data<=16'd10241;
      70056:data<=16'd9602;
      70057:data<=16'd9034;
      70058:data<=16'd8437;
      70059:data<=16'd8076;
      70060:data<=16'd7457;
      70061:data<=16'd7025;
      70062:data<=16'd7141;
      70063:data<=16'd5912;
      70064:data<=16'd3559;
      70065:data<=16'd2999;
      70066:data<=16'd3200;
      70067:data<=16'd2302;
      70068:data<=16'd2187;
      70069:data<=16'd2003;
      70070:data<=16'd312;
      70071:data<=-16'd490;
      70072:data<=-16'd667;
      70073:data<=-16'd1115;
      70074:data<=-16'd816;
      70075:data<=-16'd1187;
      70076:data<=-16'd2359;
      70077:data<=-16'd3234;
      70078:data<=-16'd3973;
      70079:data<=-16'd3668;
      70080:data<=-16'd3375;
      70081:data<=-16'd3832;
      70082:data<=-16'd3962;
      70083:data<=-16'd6141;
      70084:data<=-16'd9586;
      70085:data<=-16'd10198;
      70086:data<=-16'd9473;
      70087:data<=-16'd9338;
      70088:data<=-16'd9697;
      70089:data<=-16'd10787;
      70090:data<=-16'd11107;
      70091:data<=-16'd10643;
      70092:data<=-16'd10461;
      70093:data<=-16'd10008;
      70094:data<=-16'd9973;
      70095:data<=-16'd11062;
      70096:data<=-16'd11949;
      70097:data<=-16'd11321;
      70098:data<=-16'd10364;
      70099:data<=-16'd10504;
      70100:data<=-16'd10185;
      70101:data<=-16'd10342;
      70102:data<=-16'd12060;
      70103:data<=-16'd11597;
      70104:data<=-16'd10372;
      70105:data<=-16'd10903;
      70106:data<=-16'd10096;
      70107:data<=-16'd10126;
      70108:data<=-16'd11984;
      70109:data<=-16'd11520;
      70110:data<=-16'd10988;
      70111:data<=-16'd11226;
      70112:data<=-16'd10210;
      70113:data<=-16'd10654;
      70114:data<=-16'd11850;
      70115:data<=-16'd11825;
      70116:data<=-16'd11303;
      70117:data<=-16'd8869;
      70118:data<=-16'd6188;
      70119:data<=-16'd6076;
      70120:data<=-16'd7021;
      70121:data<=-16'd7780;
      70122:data<=-16'd7647;
      70123:data<=-16'd7197;
      70124:data<=-16'd7370;
      70125:data<=-16'd6745;
      70126:data<=-16'd6872;
      70127:data<=-16'd8504;
      70128:data<=-16'd8349;
      70129:data<=-16'd7614;
      70130:data<=-16'd7829;
      70131:data<=-16'd7238;
      70132:data<=-16'd7394;
      70133:data<=-16'd8765;
      70134:data<=-16'd8807;
      70135:data<=-16'd8222;
      70136:data<=-16'd8202;
      70137:data<=-16'd7729;
      70138:data<=-16'd7379;
      70139:data<=-16'd8354;
      70140:data<=-16'd8890;
      70141:data<=-16'd8047;
      70142:data<=-16'd7884;
      70143:data<=-16'd7887;
      70144:data<=-16'd7209;
      70145:data<=-16'd7808;
      70146:data<=-16'd8455;
      70147:data<=-16'd7815;
      70148:data<=-16'd7670;
      70149:data<=-16'd7404;
      70150:data<=-16'd7791;
      70151:data<=-16'd10698;
      70152:data<=-16'd12575;
      70153:data<=-16'd11970;
      70154:data<=-16'd11720;
      70155:data<=-16'd11489;
      70156:data<=-16'd10460;
      70157:data<=-16'd9618;
      70158:data<=-16'd9162;
      70159:data<=-16'd8805;
      70160:data<=-16'd8131;
      70161:data<=-16'd7580;
      70162:data<=-16'd7568;
      70163:data<=-16'd6746;
      70164:data<=-16'd5063;
      70165:data<=-16'd3873;
      70166:data<=-16'd3245;
      70167:data<=-16'd2961;
      70168:data<=-16'd2921;
      70169:data<=-16'd2596;
      70170:data<=-16'd1428;
      70171:data<=16'd180;
      70172:data<=16'd746;
      70173:data<=16'd499;
      70174:data<=16'd651;
      70175:data<=16'd808;
      70176:data<=16'd1551;
      70177:data<=16'd3118;
      70178:data<=16'd3422;
      70179:data<=16'd2980;
      70180:data<=16'd3316;
      70181:data<=16'd3216;
      70182:data<=16'd3196;
      70183:data<=16'd5116;
      70184:data<=16'd7908;
      70185:data<=16'd9579;
      70186:data<=16'd9635;
      70187:data<=16'd9027;
      70188:data<=16'd9071;
      70189:data<=16'd10011;
      70190:data<=16'd10948;
      70191:data<=16'd10657;
      70192:data<=16'd9717;
      70193:data<=16'd9535;
      70194:data<=16'd9491;
      70195:data<=16'd9891;
      70196:data<=16'd11166;
      70197:data<=16'd10928;
      70198:data<=16'd9926;
      70199:data<=16'd10140;
      70200:data<=16'd9570;
      70201:data<=16'd9379;
      70202:data<=16'd11033;
      70203:data<=16'd10989;
      70204:data<=16'd10149;
      70205:data<=16'd10608;
      70206:data<=16'd9752;
      70207:data<=16'd9303;
      70208:data<=16'd11094;
      70209:data<=16'd11620;
      70210:data<=16'd11039;
      70211:data<=16'd10712;
      70212:data<=16'd9805;
      70213:data<=16'd9979;
      70214:data<=16'd11121;
      70215:data<=16'd11379;
      70216:data<=16'd11253;
      70217:data<=16'd9652;
      70218:data<=16'd6487;
      70219:data<=16'd5092;
      70220:data<=16'd5856;
      70221:data<=16'd6755;
      70222:data<=16'd7004;
      70223:data<=16'd6677;
      70224:data<=16'd6270;
      70225:data<=16'd5883;
      70226:data<=16'd6122;
      70227:data<=16'd7235;
      70228:data<=16'd7542;
      70229:data<=16'd7075;
      70230:data<=16'd6775;
      70231:data<=16'd6005;
      70232:data<=16'd5944;
      70233:data<=16'd7329;
      70234:data<=16'd7850;
      70235:data<=16'd7283;
      70236:data<=16'd7115;
      70237:data<=16'd6843;
      70238:data<=16'd6317;
      70239:data<=16'd6758;
      70240:data<=16'd7573;
      70241:data<=16'd7233;
      70242:data<=16'd6690;
      70243:data<=16'd6539;
      70244:data<=16'd5791;
      70245:data<=16'd5765;
      70246:data<=16'd6819;
      70247:data<=16'd6909;
      70248:data<=16'd6457;
      70249:data<=16'd6081;
      70250:data<=16'd6225;
      70251:data<=16'd8593;
      70252:data<=16'd10941;
      70253:data<=16'd10837;
      70254:data<=16'd10238;
      70255:data<=16'd9626;
      70256:data<=16'd8853;
      70257:data<=16'd8765;
      70258:data<=16'd8153;
      70259:data<=16'd7124;
      70260:data<=16'd6875;
      70261:data<=16'd6420;
      70262:data<=16'd5858;
      70263:data<=16'd5535;
      70264:data<=16'd3941;
      70265:data<=16'd1985;
      70266:data<=16'd1683;
      70267:data<=16'd1568;
      70268:data<=16'd883;
      70269:data<=16'd951;
      70270:data<=16'd146;
      70271:data<=-16'd1835;
      70272:data<=-16'd2061;
      70273:data<=-16'd1933;
      70274:data<=-16'd2758;
      70275:data<=-16'd2390;
      70276:data<=-16'd2726;
      70277:data<=-16'd4669;
      70278:data<=-16'd5162;
      70279:data<=-16'd4892;
      70280:data<=-16'd4948;
      70281:data<=-16'd4642;
      70282:data<=-16'd4916;
      70283:data<=-16'd6296;
      70284:data<=-16'd8833;
      70285:data<=-16'd10986;
      70286:data<=-16'd10793;
      70287:data<=-16'd10355;
      70288:data<=-16'd10627;
      70289:data<=-16'd10793;
      70290:data<=-16'd11756;
      70291:data<=-16'd11991;
      70292:data<=-16'd11229;
      70293:data<=-16'd11320;
      70294:data<=-16'd10839;
      70295:data<=-16'd10693;
      70296:data<=-16'd12231;
      70297:data<=-16'd12498;
      70298:data<=-16'd11797;
      70299:data<=-16'd11455;
      70300:data<=-16'd10475;
      70301:data<=-16'd10624;
      70302:data<=-16'd12123;
      70303:data<=-16'd12446;
      70304:data<=-16'd11897;
      70305:data<=-16'd11438;
      70306:data<=-16'd10962;
      70307:data<=-16'd11027;
      70308:data<=-16'd12116;
      70309:data<=-16'd13121;
      70310:data<=-16'd12628;
      70311:data<=-16'd11893;
      70312:data<=-16'd11931;
      70313:data<=-16'd11389;
      70314:data<=-16'd11169;
      70315:data<=-16'd12531;
      70316:data<=-16'd13154;
      70317:data<=-16'd11192;
      70318:data<=-16'd7906;
      70319:data<=-16'd6018;
      70320:data<=-16'd6683;
      70321:data<=-16'd8008;
      70322:data<=-16'd8279;
      70323:data<=-16'd7747;
      70324:data<=-16'd7197;
      70325:data<=-16'd7043;
      70326:data<=-16'd7365;
      70327:data<=-16'd8278;
      70328:data<=-16'd8724;
      70329:data<=-16'd7903;
      70330:data<=-16'd7511;
      70331:data<=-16'd7673;
      70332:data<=-16'd7303;
      70333:data<=-16'd7864;
      70334:data<=-16'd8790;
      70335:data<=-16'd8194;
      70336:data<=-16'd7821;
      70337:data<=-16'd7906;
      70338:data<=-16'd7024;
      70339:data<=-16'd7071;
      70340:data<=-16'd8166;
      70341:data<=-16'd8056;
      70342:data<=-16'd7692;
      70343:data<=-16'd7454;
      70344:data<=-16'd6504;
      70345:data<=-16'd6605;
      70346:data<=-16'd7535;
      70347:data<=-16'd7344;
      70348:data<=-16'd6783;
      70349:data<=-16'd6135;
      70350:data<=-16'd6394;
      70351:data<=-16'd9250;
      70352:data<=-16'd11441;
      70353:data<=-16'd10948;
      70354:data<=-16'd10516;
      70355:data<=-16'd10198;
      70356:data<=-16'd9306;
      70357:data<=-16'd8793;
      70358:data<=-16'd8099;
      70359:data<=-16'd7479;
      70360:data<=-16'd7292;
      70361:data<=-16'd6467;
      70362:data<=-16'd5703;
      70363:data<=-16'd5418;
      70364:data<=-16'd4231;
      70365:data<=-16'd2579;
      70366:data<=-16'd1764;
      70367:data<=-16'd1175;
      70368:data<=-16'd473;
      70369:data<=-16'd522;
      70370:data<=-16'd246;
      70371:data<=16'd1474;
      70372:data<=16'd2572;
      70373:data<=16'd2419;
      70374:data<=16'd2490;
      70375:data<=16'd2502;
      70376:data<=16'd2855;
      70377:data<=16'd4305;
      70378:data<=16'd5253;
      70379:data<=16'd4965;
      70380:data<=16'd4857;
      70381:data<=16'd5294;
      70382:data<=16'd5216;
      70383:data<=16'd6109;
      70384:data<=16'd9539;
      70385:data<=16'd11617;
      70386:data<=16'd11062;
      70387:data<=16'd11185;
      70388:data<=16'd10881;
      70389:data<=16'd10611;
      70390:data<=16'd12372;
      70391:data<=16'd12551;
      70392:data<=16'd11694;
      70393:data<=16'd12182;
      70394:data<=16'd11267;
      70395:data<=16'd11051;
      70396:data<=16'd13156;
      70397:data<=16'd13295;
      70398:data<=16'd12193;
      70399:data<=16'd12023;
      70400:data<=16'd11597;
      70401:data<=16'd11468;
      70402:data<=16'd12333;
      70403:data<=16'd13233;
      70404:data<=16'd12932;
      70405:data<=16'd12069;
      70406:data<=16'd12005;
      70407:data<=16'd11570;
      70408:data<=16'd11762;
      70409:data<=16'd13679;
      70410:data<=16'd13840;
      70411:data<=16'd12759;
      70412:data<=16'd12692;
      70413:data<=16'd11903;
      70414:data<=16'd11756;
      70415:data<=16'd13470;
      70416:data<=16'd13999;
      70417:data<=16'd12007;
      70418:data<=16'd8742;
      70419:data<=16'd6959;
      70420:data<=16'd7733;
      70421:data<=16'd8805;
      70422:data<=16'd9094;
      70423:data<=16'd8519;
      70424:data<=16'd7908;
      70425:data<=16'd8190;
      70426:data<=16'd7858;
      70427:data<=16'd7961;
      70428:data<=16'd9371;
      70429:data<=16'd9244;
      70430:data<=16'd8696;
      70431:data<=16'd8652;
      70432:data<=16'd7474;
      70433:data<=16'd7959;
      70434:data<=16'd9785;
      70435:data<=16'd9385;
      70436:data<=16'd8815;
      70437:data<=16'd8693;
      70438:data<=16'd7664;
      70439:data<=16'd8028;
      70440:data<=16'd9353;
      70441:data<=16'd9148;
      70442:data<=16'd8458;
      70443:data<=16'd8122;
      70444:data<=16'd7638;
      70445:data<=16'd7495;
      70446:data<=16'd7938;
      70447:data<=16'd8429;
      70448:data<=16'd8241;
      70449:data<=16'd7404;
      70450:data<=16'd7796;
      70451:data<=16'd9937;
      70452:data<=16'd11441;
      70453:data<=16'd11838;
      70454:data<=16'd12032;
      70455:data<=16'd11159;
      70456:data<=16'd9962;
      70457:data<=16'd9694;
      70458:data<=16'd9271;
      70459:data<=16'd8763;
      70460:data<=16'd8425;
      70461:data<=16'd7374;
      70462:data<=16'd6584;
      70463:data<=16'd6476;
      70464:data<=16'd5639;
      70465:data<=16'd4021;
      70466:data<=16'd2689;
      70467:data<=16'd2218;
      70468:data<=16'd2112;
      70469:data<=16'd1730;
      70470:data<=16'd1104;
      70471:data<=-16'd126;
      70472:data<=-16'd1290;
      70473:data<=-16'd1269;
      70474:data<=-16'd1533;
      70475:data<=-16'd2337;
      70476:data<=-16'd2029;
      70477:data<=-16'd2358;
      70478:data<=-16'd4132;
      70479:data<=-16'd4397;
      70480:data<=-16'd4037;
      70481:data<=-16'd4728;
      70482:data<=-16'd4144;
      70483:data<=-16'd4554;
      70484:data<=-16'd8658;
      70485:data<=-16'd10994;
      70486:data<=-16'd10155;
      70487:data<=-16'd10040;
      70488:data<=-16'd9671;
      70489:data<=-16'd9691;
      70490:data<=-16'd11526;
      70491:data<=-16'd11822;
      70492:data<=-16'd10863;
      70493:data<=-16'd10702;
      70494:data<=-16'd10228;
      70495:data<=-16'd10298;
      70496:data<=-16'd11383;
      70497:data<=-16'd11797;
      70498:data<=-16'd11403;
      70499:data<=-16'd11071;
      70500:data<=-16'd10951;
      70501:data<=-16'd10137;
      70502:data<=-16'd9994;
      70503:data<=-16'd11843;
      70504:data<=-16'd12272;
      70505:data<=-16'd11298;
      70506:data<=-16'd11264;
      70507:data<=-16'd10285;
      70508:data<=-16'd10290;
      70509:data<=-16'd12645;
      70510:data<=-16'd12836;
      70511:data<=-16'd11496;
      70512:data<=-16'd11235;
      70513:data<=-16'd10989;
      70514:data<=-16'd11092;
      70515:data<=-16'd11896;
      70516:data<=-16'd12460;
      70517:data<=-16'd10950;
      70518:data<=-16'd7668;
      70519:data<=-16'd6567;
      70520:data<=-16'd6821;
      70521:data<=-16'd6598;
      70522:data<=-16'd7884;
      70523:data<=-16'd8341;
      70524:data<=-16'd7439;
      70525:data<=-16'd7689;
      70526:data<=-16'd6909;
      70527:data<=-16'd6727;
      70528:data<=-16'd8886;
      70529:data<=-16'd8963;
      70530:data<=-16'd7915;
      70531:data<=-16'd7884;
      70532:data<=-16'd7242;
      70533:data<=-16'd7759;
      70534:data<=-16'd9156;
      70535:data<=-16'd8830;
      70536:data<=-16'd8205;
      70537:data<=-16'd8081;
      70538:data<=-16'd7723;
      70539:data<=-16'd7618;
      70540:data<=-16'd8249;
      70541:data<=-16'd9162;
      70542:data<=-16'd9025;
      70543:data<=-16'd8153;
      70544:data<=-16'd7697;
      70545:data<=-16'd7142;
      70546:data<=-16'd7228;
      70547:data<=-16'd8567;
      70548:data<=-16'd8702;
      70549:data<=-16'd7366;
      70550:data<=-16'd7920;
      70551:data<=-16'd10478;
      70552:data<=-16'd11826;
      70553:data<=-16'd11991;
      70554:data<=-16'd12073;
      70555:data<=-16'd11109;
      70556:data<=-16'd10425;
      70557:data<=-16'd10613;
      70558:data<=-16'd9633;
      70559:data<=-16'd8822;
      70560:data<=-16'd8872;
      70561:data<=-16'd7949;
      70562:data<=-16'd7238;
      70563:data<=-16'd6998;
      70564:data<=-16'd5827;
      70565:data<=-16'd4505;
      70566:data<=-16'd3447;
      70567:data<=-16'd2757;
      70568:data<=-16'd2437;
      70569:data<=-16'd2120;
      70570:data<=-16'd2305;
      70571:data<=-16'd1535;
      70572:data<=16'd487;
      70573:data<=16'd1057;
      70574:data<=16'd1131;
      70575:data<=16'd1538;
      70576:data<=16'd840;
      70577:data<=16'd1451;
      70578:data<=16'd3521;
      70579:data<=16'd3721;
      70580:data<=16'd3482;
      70581:data<=16'd3824;
      70582:data<=16'd3265;
      70583:data<=16'd4469;
      70584:data<=16'd8382;
      70585:data<=16'd10389;
      70586:data<=16'd9693;
      70587:data<=16'd9479;
      70588:data<=16'd9547;
      70589:data<=16'd9198;
      70590:data<=16'd9838;
      70591:data<=16'd10615;
      70592:data<=16'd10358;
      70593:data<=16'd10383;
      70594:data<=16'd10266;
      70595:data<=16'd9256;
      70596:data<=16'd9579;
      70597:data<=16'd10963;
      70598:data<=16'd10837;
      70599:data<=16'd10358;
      70600:data<=16'd10219;
      70601:data<=16'd9232;
      70602:data<=16'd9589;
      70603:data<=16'd11395;
      70604:data<=16'd11303;
      70605:data<=16'd10493;
      70606:data<=16'd10390;
      70607:data<=16'd9694;
      70608:data<=16'd9837;
      70609:data<=16'd11188;
      70610:data<=16'd11629;
      70611:data<=16'd11203;
      70612:data<=16'd10687;
      70613:data<=16'd10210;
      70614:data<=16'd9602;
      70615:data<=16'd9756;
      70616:data<=16'd11268;
      70617:data<=16'd10311;
      70618:data<=16'd6673;
      70619:data<=16'd5473;
      70620:data<=16'd5568;
      70621:data<=16'd5567;
      70622:data<=16'd7300;
      70623:data<=16'd7638;
      70624:data<=16'd6511;
      70625:data<=16'd6666;
      70626:data<=16'd5984;
      70627:data<=16'd5873;
      70628:data<=16'd7703;
      70629:data<=16'd7692;
      70630:data<=16'd6945;
      70631:data<=16'd7188;
      70632:data<=16'd6464;
      70633:data<=16'd6255;
      70634:data<=16'd7507;
      70635:data<=16'd8085;
      70636:data<=16'd7639;
      70637:data<=16'd7015;
      70638:data<=16'd6546;
      70639:data<=16'd6140;
      70640:data<=16'd6451;
      70641:data<=16'd7661;
      70642:data<=16'd7677;
      70643:data<=16'd6883;
      70644:data<=16'd6953;
      70645:data<=16'd6458;
      70646:data<=16'd6279;
      70647:data<=16'd7747;
      70648:data<=16'd7674;
      70649:data<=16'd6419;
      70650:data<=16'd7738;
      70651:data<=16'd9994;
      70652:data<=16'd10507;
      70653:data<=16'd10527;
      70654:data<=16'd10748;
      70655:data<=16'd10492;
      70656:data<=16'd9991;
      70657:data<=16'd9321;
      70658:data<=16'd8526;
      70659:data<=16'd8011;
      70660:data<=16'd7544;
      70661:data<=16'd7113;
      70662:data<=16'd6604;
      70663:data<=16'd5788;
      70664:data<=16'd5523;
      70665:data<=16'd4836;
      70666:data<=16'd2716;
      70667:data<=16'd1717;
      70668:data<=16'd1858;
      70669:data<=16'd1447;
      70670:data<=16'd1633;
      70671:data<=16'd754;
      70672:data<=-16'd1859;
      70673:data<=-16'd2296;
      70674:data<=-16'd1679;
      70675:data<=-16'd2147;
      70676:data<=-16'd1851;
      70677:data<=-16'd2426;
      70678:data<=-16'd4419;
      70679:data<=-16'd4840;
      70680:data<=-16'd4772;
      70681:data<=-16'd4951;
      70682:data<=-16'd4202;
      70683:data<=-16'd5174;
      70684:data<=-16'd8828;
      70685:data<=-16'd11277;
      70686:data<=-16'd11110;
      70687:data<=-16'd10678;
      70688:data<=-16'd10455;
      70689:data<=-16'd9740;
      70690:data<=-16'd10298;
      70691:data<=-16'd11890;
      70692:data<=-16'd11932;
      70693:data<=-16'd11471;
      70694:data<=-16'd11183;
      70695:data<=-16'd10337;
      70696:data<=-16'd11016;
      70697:data<=-16'd12468;
      70698:data<=-16'd12339;
      70699:data<=-16'd12148;
      70700:data<=-16'd11840;
      70701:data<=-16'd10927;
      70702:data<=-16'd11283;
      70703:data<=-16'd12337;
      70704:data<=-16'd12772;
      70705:data<=-16'd12486;
      70706:data<=-16'd11743;
      70707:data<=-16'd11414;
      70708:data<=-16'd11022;
      70709:data<=-16'd11301;
      70710:data<=-16'd13039;
      70711:data<=-16'd13135;
      70712:data<=-16'd12149;
      70713:data<=-16'd12184;
      70714:data<=-16'd11012;
      70715:data<=-16'd10894;
      70716:data<=-16'd12907;
      70717:data<=-16'd11168;
      70718:data<=-16'd7474;
      70719:data<=-16'd6880;
      70720:data<=-16'd6754;
      70721:data<=-16'd6573;
      70722:data<=-16'd7932;
      70723:data<=-16'd8584;
      70724:data<=-16'd8210;
      70725:data<=-16'd7949;
      70726:data<=-16'd7233;
      70727:data<=-16'd6992;
      70728:data<=-16'd8208;
      70729:data<=-16'd9072;
      70730:data<=-16'd8545;
      70731:data<=-16'd7953;
      70732:data<=-16'd7492;
      70733:data<=-16'd6887;
      70734:data<=-16'd7574;
      70735:data<=-16'd8960;
      70736:data<=-16'd8754;
      70737:data<=-16'd7975;
      70738:data<=-16'd7928;
      70739:data<=-16'd7442;
      70740:data<=-16'd7285;
      70741:data<=-16'd8463;
      70742:data<=-16'd8683;
      70743:data<=-16'd7832;
      70744:data<=-16'd7903;
      70745:data<=-16'd7371;
      70746:data<=-16'd6623;
      70747:data<=-16'd8144;
      70748:data<=-16'd8671;
      70749:data<=-16'd7225;
      70750:data<=-16'd8396;
      70751:data<=-16'd10666;
      70752:data<=-16'd11060;
      70753:data<=-16'd11670;
      70754:data<=-16'd12099;
      70755:data<=-16'd11185;
      70756:data<=-16'd10473;
      70757:data<=-16'd10066;
      70758:data<=-16'd9561;
      70759:data<=-16'd8966;
      70760:data<=-16'd8196;
      70761:data<=-16'd7827;
      70762:data<=-16'd7326;
      70763:data<=-16'd6667;
      70764:data<=-16'd6626;
      70765:data<=-16'd5524;
      70766:data<=-16'd3366;
      70767:data<=-16'd2807;
      70768:data<=-16'd3055;
      70769:data<=-16'd2584;
      70770:data<=-16'd2337;
      70771:data<=-16'd1536;
      70772:data<=16'd452;
      70773:data<=16'd1313;
      70774:data<=16'd1033;
      70775:data<=16'd1340;
      70776:data<=16'd1265;
      70777:data<=16'd1224;
      70778:data<=16'd2810;
      70779:data<=16'd3985;
      70780:data<=16'd3918;
      70781:data<=16'd4067;
      70782:data<=16'd3582;
      70783:data<=16'd3971;
      70784:data<=16'd7899;
      70785:data<=16'd11256;
      70786:data<=16'd10806;
      70787:data<=16'd10152;
      70788:data<=16'd10140;
      70789:data<=16'd9374;
      70790:data<=16'd10249;
      70791:data<=16'd12061;
      70792:data<=16'd11835;
      70793:data<=16'd11447;
      70794:data<=16'd11394;
      70795:data<=16'd10292;
      70796:data<=16'd10360;
      70797:data<=16'd11697;
      70798:data<=16'd12167;
      70799:data<=16'd12201;
      70800:data<=16'd11996;
      70801:data<=16'd11383;
      70802:data<=16'd10859;
      70803:data<=16'd11317;
      70804:data<=16'd12828;
      70805:data<=16'd12728;
      70806:data<=16'd11629;
      70807:data<=16'd11819;
      70808:data<=16'd10992;
      70809:data<=16'd11018;
      70810:data<=16'd13673;
      70811:data<=16'd13521;
      70812:data<=16'd11988;
      70813:data<=16'd12383;
      70814:data<=16'd11330;
      70815:data<=16'd11163;
      70816:data<=16'd13082;
      70817:data<=16'd11637;
      70818:data<=16'd8625;
      70819:data<=16'd7958;
      70820:data<=16'd7824;
      70821:data<=16'd7843;
      70822:data<=16'd9095;
      70823:data<=16'd10014;
      70824:data<=16'd9132;
      70825:data<=16'd8539;
      70826:data<=16'd9025;
      70827:data<=16'd8498;
      70828:data<=16'd8809;
      70829:data<=16'd10396;
      70830:data<=16'd9908;
      70831:data<=16'd9247;
      70832:data<=16'd9362;
      70833:data<=16'd8349;
      70834:data<=16'd8707;
      70835:data<=16'd10122;
      70836:data<=16'd10029;
      70837:data<=16'd9767;
      70838:data<=16'd9317;
      70839:data<=16'd8443;
      70840:data<=16'd8648;
      70841:data<=16'd9749;
      70842:data<=16'd10329;
      70843:data<=16'd9480;
      70844:data<=16'd8828;
      70845:data<=16'd8936;
      70846:data<=16'd8384;
      70847:data<=16'd9233;
      70848:data<=16'd10342;
      70849:data<=16'd8780;
      70850:data<=16'd9265;
      70851:data<=16'd12169;
      70852:data<=16'd12330;
      70853:data<=16'd11991;
      70854:data<=16'd13018;
      70855:data<=16'd12871;
      70856:data<=16'd11961;
      70857:data<=16'd11311;
      70858:data<=16'd10561;
      70859:data<=16'd9630;
      70860:data<=16'd9063;
      70861:data<=16'd9118;
      70862:data<=16'd8596;
      70863:data<=16'd7729;
      70864:data<=16'd7459;
      70865:data<=16'd6593;
      70866:data<=16'd5124;
      70867:data<=16'd4190;
      70868:data<=16'd3580;
      70869:data<=16'd3177;
      70870:data<=16'd3151;
      70871:data<=16'd2883;
      70872:data<=16'd1434;
      70873:data<=-16'd111;
      70874:data<=-16'd200;
      70875:data<=-16'd328;
      70876:data<=-16'd746;
      70877:data<=-16'd355;
      70878:data<=-16'd1201;
      70879:data<=-16'd3077;
      70880:data<=-16'd3344;
      70881:data<=-16'd2966;
      70882:data<=-16'd3022;
      70883:data<=-16'd3973;
      70884:data<=-16'd7095;
      70885:data<=-16'd9805;
      70886:data<=-16'd9542;
      70887:data<=-16'd9159;
      70888:data<=-16'd9703;
      70889:data<=-16'd9013;
      70890:data<=-16'd8711;
      70891:data<=-16'd10128;
      70892:data<=-16'd10611;
      70893:data<=-16'd10205;
      70894:data<=-16'd10343;
      70895:data<=-16'd9875;
      70896:data<=-16'd9280;
      70897:data<=-16'd10096;
      70898:data<=-16'd11297;
      70899:data<=-16'd11186;
      70900:data<=-16'd10420;
      70901:data<=-16'd10648;
      70902:data<=-16'd10633;
      70903:data<=-16'd10187;
      70904:data<=-16'd11201;
      70905:data<=-16'd11380;
      70906:data<=-16'd10546;
      70907:data<=-16'd11150;
      70908:data<=-16'd10498;
      70909:data<=-16'd9746;
      70910:data<=-16'd11552;
      70911:data<=-16'd11870;
      70912:data<=-16'd11273;
      70913:data<=-16'd11606;
      70914:data<=-16'd10473;
      70915:data<=-16'd10357;
      70916:data<=-16'd11470;
      70917:data<=-16'd9834;
      70918:data<=-16'd7288;
      70919:data<=-16'd6452;
      70920:data<=-16'd6616;
      70921:data<=-16'd6446;
      70922:data<=-16'd6337;
      70923:data<=-16'd7556;
      70924:data<=-16'd7799;
      70925:data<=-16'd7157;
      70926:data<=-16'd7703;
      70927:data<=-16'd6890;
      70928:data<=-16'd6390;
      70929:data<=-16'd8202;
      70930:data<=-16'd8273;
      70931:data<=-16'd7705;
      70932:data<=-16'd7821;
      70933:data<=-16'd6701;
      70934:data<=-16'd7007;
      70935:data<=-16'd8476;
      70936:data<=-16'd8364;
      70937:data<=-16'd7908;
      70938:data<=-16'd7583;
      70939:data<=-16'd7289;
      70940:data<=-16'd7171;
      70941:data<=-16'd7732;
      70942:data<=-16'd8937;
      70943:data<=-16'd8228;
      70944:data<=-16'd7394;
      70945:data<=-16'd7918;
      70946:data<=-16'd6626;
      70947:data<=-16'd6719;
      70948:data<=-16'd8660;
      70949:data<=-16'd7488;
      70950:data<=-16'd7975;
      70951:data<=-16'd11427;
      70952:data<=-16'd11257;
      70953:data<=-16'd10198;
      70954:data<=-16'd11602;
      70955:data<=-16'd11908;
      70956:data<=-16'd10883;
      70957:data<=-16'd10420;
      70958:data<=-16'd9917;
      70959:data<=-16'd9009;
      70960:data<=-16'd8569;
      70961:data<=-16'd8263;
      70962:data<=-16'd7485;
      70963:data<=-16'd7275;
      70964:data<=-16'd7374;
      70965:data<=-16'd6774;
      70966:data<=-16'd5459;
      70967:data<=-16'd3788;
      70968:data<=-16'd3494;
      70969:data<=-16'd3694;
      70970:data<=-16'd2714;
      70971:data<=-16'd2739;
      70972:data<=-16'd2149;
      70973:data<=16'd340;
      70974:data<=16'd661;
      70975:data<=16'd146;
      70976:data<=16'd640;
      70977:data<=16'd318;
      70978:data<=16'd1066;
      70979:data<=16'd2617;
      70980:data<=16'd3098;
      70981:data<=16'd3283;
      70982:data<=16'd2582;
      70983:data<=16'd3154;
      70984:data<=16'd6610;
      70985:data<=16'd9088;
      70986:data<=16'd9556;
      70987:data<=16'd9259;
      70988:data<=16'd8812;
      70989:data<=16'd8792;
      70990:data<=16'd8288;
      70991:data<=16'd8900;
      70992:data<=16'd10731;
      70993:data<=16'd10339;
      70994:data<=16'd9687;
      70995:data<=16'd10085;
      70996:data<=16'd9191;
      70997:data<=16'd9370;
      70998:data<=16'd11122;
      70999:data<=16'd11203;
      71000:data<=16'd10611;
      71001:data<=16'd10466;
      71002:data<=16'd9785;
      71003:data<=16'd9841;
      71004:data<=16'd11171;
      71005:data<=16'd11593;
      71006:data<=16'd11030;
      71007:data<=16'd10728;
      71008:data<=16'd10038;
      71009:data<=16'd10046;
      71010:data<=16'd11543;
      71011:data<=16'd11847;
      71012:data<=16'd11326;
      71013:data<=16'd11479;
      71014:data<=16'd10919;
      71015:data<=16'd10460;
      71016:data<=16'd10420;
      71017:data<=16'd8997;
      71018:data<=16'd7283;
      71019:data<=16'd6821;
      71020:data<=16'd6857;
      71021:data<=16'd6208;
      71022:data<=16'd5906;
      71023:data<=16'd7225;
      71024:data<=16'd7639;
      71025:data<=16'd6980;
      71026:data<=16'd7218;
      71027:data<=16'd6460;
      71028:data<=16'd6006;
      71029:data<=16'd7594;
      71030:data<=16'd7718;
      71031:data<=16'd6687;
      71032:data<=16'd6378;
      71033:data<=16'd6043;
      71034:data<=16'd6352;
      71035:data<=16'd6884;
      71036:data<=16'd7065;
      71037:data<=16'd7071;
      71038:data<=16'd6605;
      71039:data<=16'd6520;
      71040:data<=16'd5938;
      71041:data<=16'd5752;
      71042:data<=16'd7630;
      71043:data<=16'd7580;
      71044:data<=16'd6375;
      71045:data<=16'd6724;
      71046:data<=16'd5655;
      71047:data<=16'd5883;
      71048:data<=16'd7667;
      71049:data<=16'd6517;
      71050:data<=16'd7492;
      71051:data<=16'd10619;
      71052:data<=16'd9940;
      71053:data<=16'd9626;
      71054:data<=16'd11250;
      71055:data<=16'd11189;
      71056:data<=16'd10613;
      71057:data<=16'd10178;
      71058:data<=16'd9649;
      71059:data<=16'd9162;
      71060:data<=16'd8328;
      71061:data<=16'd8234;
      71062:data<=16'd8149;
      71063:data<=16'd6978;
      71064:data<=16'd6642;
      71065:data<=16'd7110;
      71066:data<=16'd5841;
      71067:data<=16'd3513;
      71068:data<=16'd3068;
      71069:data<=16'd3242;
      71070:data<=16'd2223;
      71071:data<=16'd2130;
      71072:data<=16'd1845;
      71073:data<=-16'd180;
      71074:data<=-16'd1177;
      71075:data<=-16'd1225;
      71076:data<=-16'd1225;
      71077:data<=-16'd1077;
      71078:data<=-16'd2162;
      71079:data<=-16'd3380;
      71080:data<=-16'd4074;
      71081:data<=-16'd4272;
      71082:data<=-16'd3353;
      71083:data<=-16'd4578;
      71084:data<=-16'd7573;
      71085:data<=-16'd8904;
      71086:data<=-16'd9969;
      71087:data<=-16'd10222;
      71088:data<=-16'd9562;
      71089:data<=-16'd9650;
      71090:data<=-16'd8722;
      71091:data<=-16'd8925;
      71092:data<=-16'd11109;
      71093:data<=-16'd11153;
      71094:data<=-16'd10713;
      71095:data<=-16'd10848;
      71096:data<=-16'd10035;
      71097:data<=-16'd10296;
      71098:data<=-16'd11348;
      71099:data<=-16'd12032;
      71100:data<=-16'd12117;
      71101:data<=-16'd10968;
      71102:data<=-16'd10493;
      71103:data<=-16'd10986;
      71104:data<=-16'd11650;
      71105:data<=-16'd12345;
      71106:data<=-16'd11471;
      71107:data<=-16'd10906;
      71108:data<=-16'd11238;
      71109:data<=-16'd10151;
      71110:data<=-16'd10416;
      71111:data<=-16'd12082;
      71112:data<=-16'd12125;
      71113:data<=-16'd11926;
      71114:data<=-16'd11611;
      71115:data<=-16'd11091;
      71116:data<=-16'd10627;
      71117:data<=-16'd8639;
      71118:data<=-16'd7312;
      71119:data<=-16'd7884;
      71120:data<=-16'd7494;
      71121:data<=-16'd6229;
      71122:data<=-16'd6211;
      71123:data<=-16'd7764;
      71124:data<=-16'd8549;
      71125:data<=-16'd7723;
      71126:data<=-16'd7577;
      71127:data<=-16'd7326;
      71128:data<=-16'd6734;
      71129:data<=-16'd7773;
      71130:data<=-16'd8141;
      71131:data<=-16'd7209;
      71132:data<=-16'd7366;
      71133:data<=-16'd7409;
      71134:data<=-16'd6516;
      71135:data<=-16'd6775;
      71136:data<=-16'd8470;
      71137:data<=-16'd8846;
      71138:data<=-16'd8023;
      71139:data<=-16'd8346;
      71140:data<=-16'd7561;
      71141:data<=-16'd6508;
      71142:data<=-16'd8519;
      71143:data<=-16'd9224;
      71144:data<=-16'd8059;
      71145:data<=-16'd8105;
      71146:data<=-16'd6783;
      71147:data<=-16'd6375;
      71148:data<=-16'd8346;
      71149:data<=-16'd8335;
      71150:data<=-16'd9016;
      71151:data<=-16'd11582;
      71152:data<=-16'd11635;
      71153:data<=-16'd10787;
      71154:data<=-16'd11564;
      71155:data<=-16'd12610;
      71156:data<=-16'd12373;
      71157:data<=-16'd10951;
      71158:data<=-16'd10322;
      71159:data<=-16'd10420;
      71160:data<=-16'd9996;
      71161:data<=-16'd9417;
      71162:data<=-16'd8804;
      71163:data<=-16'd8216;
      71164:data<=-16'd7793;
      71165:data<=-16'd7767;
      71166:data<=-16'd6902;
      71167:data<=-16'd4102;
      71168:data<=-16'd3272;
      71169:data<=-16'd4420;
      71170:data<=-16'd3175;
      71171:data<=-16'd2311;
      71172:data<=-16'd2537;
      71173:data<=-16'd726;
      71174:data<=16'd249;
      71175:data<=16'd126;
      71176:data<=16'd1140;
      71177:data<=16'd1296;
      71178:data<=16'd625;
      71179:data<=16'd1234;
      71180:data<=16'd3181;
      71181:data<=16'd4035;
      71182:data<=16'd3251;
      71183:data<=16'd4689;
      71184:data<=16'd7228;
      71185:data<=16'd7743;
      71186:data<=16'd8883;
      71187:data<=16'd10187;
      71188:data<=16'd9884;
      71189:data<=16'd9693;
      71190:data<=16'd9289;
      71191:data<=16'd9321;
      71192:data<=16'd10630;
      71193:data<=16'd11203;
      71194:data<=16'd11059;
      71195:data<=16'd10660;
      71196:data<=16'd9809;
      71197:data<=16'd9641;
      71198:data<=16'd10549;
      71199:data<=16'd11374;
      71200:data<=16'd10633;
      71201:data<=16'd9688;
      71202:data<=16'd9752;
      71203:data<=16'd9125;
      71204:data<=16'd9536;
      71205:data<=16'd11028;
      71206:data<=16'd10270;
      71207:data<=16'd9976;
      71208:data<=16'd10393;
      71209:data<=16'd8774;
      71210:data<=16'd9025;
      71211:data<=16'd11089;
      71212:data<=16'd11277;
      71213:data<=16'd11016;
      71214:data<=16'd10437;
      71215:data<=16'd9488;
      71216:data<=16'd9088;
      71217:data<=16'd7738;
      71218:data<=16'd6633;
      71219:data<=16'd7171;
      71220:data<=16'd7263;
      71221:data<=16'd6508;
      71222:data<=16'd6181;
      71223:data<=16'd6790;
      71224:data<=16'd7618;
      71225:data<=16'd7608;
      71226:data<=16'd7110;
      71227:data<=16'd6304;
      71228:data<=16'd5460;
      71229:data<=16'd5755;
      71230:data<=16'd6863;
      71231:data<=16'd7649;
      71232:data<=16'd7676;
      71233:data<=16'd6981;
      71234:data<=16'd6317;
      71235:data<=16'd6786;
      71236:data<=16'd8299;
      71237:data<=16'd8725;
      71238:data<=16'd7739;
      71239:data<=16'd7253;
      71240:data<=16'd6811;
      71241:data<=16'd6610;
      71242:data<=16'd7568;
      71243:data<=16'd7856;
      71244:data<=16'd8009;
      71245:data<=16'd8437;
      71246:data<=16'd7098;
      71247:data<=16'd6592;
      71248:data<=16'd7997;
      71249:data<=16'd8516;
      71250:data<=16'd9882;
      71251:data<=16'd11972;
      71252:data<=16'd11708;
      71253:data<=16'd10985;
      71254:data<=16'd11327;
      71255:data<=16'd11913;
      71256:data<=16'd12442;
      71257:data<=16'd11629;
      71258:data<=16'd10493;
      71259:data<=16'd10652;
      71260:data<=16'd10329;
      71261:data<=16'd9498;
      71262:data<=16'd9124;
      71263:data<=16'd8199;
      71264:data<=16'd7514;
      71265:data<=16'd7460;
      71266:data<=16'd6528;
      71267:data<=16'd5510;
      71268:data<=16'd5248;
      71269:data<=16'd4675;
      71270:data<=16'd3683;
      71271:data<=16'd2881;
      71272:data<=16'd2663;
      71273:data<=16'd2408;
      71274:data<=16'd893;
      71275:data<=-16'd479;
      71276:data<=-16'd496;
      71277:data<=-16'd622;
      71278:data<=-16'd643;
      71279:data<=-16'd745;
      71280:data<=-16'd2428;
      71281:data<=-16'd3127;
      71282:data<=-16'd2312;
      71283:data<=-16'd4165;
      71284:data<=-16'd7103;
      71285:data<=-16'd7736;
      71286:data<=-16'd8631;
      71287:data<=-16'd9771;
      71288:data<=-16'd8498;
      71289:data<=-16'd7407;
      71290:data<=-16'd8226;
      71291:data<=-16'd8671;
      71292:data<=-16'd9266;
      71293:data<=-16'd10349;
      71294:data<=-16'd9624;
      71295:data<=-16'd8672;
      71296:data<=-16'd8960;
      71297:data<=-16'd8399;
      71298:data<=-16'd8719;
      71299:data<=-16'd10687;
      71300:data<=-16'd10536;
      71301:data<=-16'd9535;
      71302:data<=-16'd9282;
      71303:data<=-16'd8091;
      71304:data<=-16'd8890;
      71305:data<=-16'd11250;
      71306:data<=-16'd10642;
      71307:data<=-16'd9920;
      71308:data<=-16'd10528;
      71309:data<=-16'd9605;
      71310:data<=-16'd9248;
      71311:data<=-16'd10473;
      71312:data<=-16'd11285;
      71313:data<=-16'd11461;
      71314:data<=-16'd10922;
      71315:data<=-16'd10269;
      71316:data<=-16'd8795;
      71317:data<=-16'd6043;
      71318:data<=-16'd5359;
      71319:data<=-16'd6143;
      71320:data<=-16'd5771;
      71321:data<=-16'd5671;
      71322:data<=-16'd5489;
      71323:data<=-16'd5532;
      71324:data<=-16'd7043;
      71325:data<=-16'd7274;
      71326:data<=-16'd6363;
      71327:data<=-16'd5915;
      71328:data<=-16'd5053;
      71329:data<=-16'd5611;
      71330:data<=-16'd7028;
      71331:data<=-16'd6492;
      71332:data<=-16'd6281;
      71333:data<=-16'd6966;
      71334:data<=-16'd6435;
      71335:data<=-16'd6529;
      71336:data<=-16'd7736;
      71337:data<=-16'd7303;
      71338:data<=-16'd6244;
      71339:data<=-16'd6643;
      71340:data<=-16'd6206;
      71341:data<=-16'd4980;
      71342:data<=-16'd5724;
      71343:data<=-16'd6267;
      71344:data<=-16'd5958;
      71345:data<=-16'd6824;
      71346:data<=-16'd6438;
      71347:data<=-16'd5369;
      71348:data<=-16'd6196;
      71349:data<=-16'd7307;
      71350:data<=-16'd9373;
      71351:data<=-16'd11341;
      71352:data<=-16'd10182;
      71353:data<=-16'd9212;
      71354:data<=-16'd9985;
      71355:data<=-16'd10627;
      71356:data<=-16'd11332;
      71357:data<=-16'd11016;
      71358:data<=-16'd10050;
      71359:data<=-16'd9609;
      71360:data<=-16'd8766;
      71361:data<=-16'd8526;
      71362:data<=-16'd8737;
      71363:data<=-16'd8254;
      71364:data<=-16'd7908;
      71365:data<=-16'd6981;
      71366:data<=-16'd5890;
      71367:data<=-16'd5233;
      71368:data<=-16'd3316;
      71369:data<=-16'd1858;
      71370:data<=-16'd2244;
      71371:data<=-16'd2391;
      71372:data<=-16'd1933;
      71373:data<=-16'd852;
      71374:data<=16'd666;
      71375:data<=16'd1265;
      71376:data<=16'd1251;
      71377:data<=16'd1165;
      71378:data<=16'd1045;
      71379:data<=16'd1895;
      71380:data<=16'd3718;
      71381:data<=16'd4261;
      71382:data<=16'd3516;
      71383:data<=16'd5074;
      71384:data<=16'd7832;
      71385:data<=16'd8247;
      71386:data<=16'd8828;
      71387:data<=16'd10257;
      71388:data<=16'd9920;
      71389:data<=16'd9309;
      71390:data<=16'd8881;
      71391:data<=16'd8396;
      71392:data<=16'd10020;
      71393:data<=16'd11906;
      71394:data<=16'd11356;
      71395:data<=16'd10331;
      71396:data<=16'd9961;
      71397:data<=16'd9085;
      71398:data<=16'd8921;
      71399:data<=16'd10774;
      71400:data<=16'd11735;
      71401:data<=16'd10483;
      71402:data<=16'd9787;
      71403:data<=16'd10031;
      71404:data<=16'd10378;
      71405:data<=16'd10866;
      71406:data<=16'd10857;
      71407:data<=16'd10790;
      71408:data<=16'd10336;
      71409:data<=16'd8787;
      71410:data<=16'd8143;
      71411:data<=16'd9624;
      71412:data<=16'd11517;
      71413:data<=16'd11273;
      71414:data<=16'd10097;
      71415:data<=16'd10328;
      71416:data<=16'd8828;
      71417:data<=16'd6601;
      71418:data<=16'd7732;
      71419:data<=16'd7655;
      71420:data<=16'd5999;
      71421:data<=16'd7009;
      71422:data<=16'd7025;
      71423:data<=16'd5959;
      71424:data<=16'd7019;
      71425:data<=16'd7210;
      71426:data<=16'd5806;
      71427:data<=16'd5682;
      71428:data<=16'd6721;
      71429:data<=16'd6352;
      71430:data<=16'd5557;
      71431:data<=16'd7494;
      71432:data<=16'd8802;
      71433:data<=16'd7474;
      71434:data<=16'd6893;
      71435:data<=16'd6645;
      71436:data<=16'd7104;
      71437:data<=16'd8008;
      71438:data<=16'd6986;
      71439:data<=16'd6892;
      71440:data<=16'd7021;
      71441:data<=16'd6363;
      71442:data<=16'd8237;
      71443:data<=16'd8589;
      71444:data<=16'd7319;
      71445:data<=16'd8590;
      71446:data<=16'd8251;
      71447:data<=16'd7191;
      71448:data<=16'd7699;
      71449:data<=16'd7480;
      71450:data<=16'd9188;
      71451:data<=16'd11191;
      71452:data<=16'd10561;
      71453:data<=16'd9720;
      71454:data<=16'd8467;
      71455:data<=16'd9320;
      71456:data<=16'd11590;
      71457:data<=16'd9841;
      71458:data<=16'd8440;
      71459:data<=16'd9042;
      71460:data<=16'd7756;
      71461:data<=16'd7086;
      71462:data<=16'd6975;
      71463:data<=16'd6021;
      71464:data<=16'd5567;
      71465:data<=16'd5618;
      71466:data<=16'd6569;
      71467:data<=16'd5162;
      71468:data<=16'd1386;
      71469:data<=16'd1425;
      71470:data<=16'd2373;
      71471:data<=16'd1383;
      71472:data<=16'd2141;
      71473:data<=16'd1642;
      71474:data<=-16'd899;
      71475:data<=-16'd654;
      71476:data<=16'd273;
      71477:data<=-16'd804;
      71478:data<=-16'd1165;
      71479:data<=-16'd1025;
      71480:data<=-16'd3175;
      71481:data<=-16'd5019;
      71482:data<=-16'd4225;
      71483:data<=-16'd5304;
      71484:data<=-16'd8408;
      71485:data<=-16'd8696;
      71486:data<=-16'd8326;
      71487:data<=-16'd10231;
      71488:data<=-16'd11274;
      71489:data<=-16'd10014;
      71490:data<=-16'd9215;
      71491:data<=-16'd9935;
      71492:data<=-16'd10789;
      71493:data<=-16'd11897;
      71494:data<=-16'd12185;
      71495:data<=-16'd10657;
      71496:data<=-16'd10354;
      71497:data<=-16'd10185;
      71498:data<=-16'd9019;
      71499:data<=-16'd11171;
      71500:data<=-16'd13066;
      71501:data<=-16'd11285;
      71502:data<=-16'd11088;
      71503:data<=-16'd11121;
      71504:data<=-16'd9521;
      71505:data<=-16'd10207;
      71506:data<=-16'd11509;
      71507:data<=-16'd11323;
      71508:data<=-16'd10848;
      71509:data<=-16'd10345;
      71510:data<=-16'd10651;
      71511:data<=-16'd11248;
      71512:data<=-16'd11574;
      71513:data<=-16'd12037;
      71514:data<=-16'd11773;
      71515:data<=-16'd11160;
      71516:data<=-16'd9591;
      71517:data<=-16'd6840;
      71518:data<=-16'd6560;
      71519:data<=-16'd8440;
      71520:data<=-16'd8784;
      71521:data<=-16'd7453;
      71522:data<=-16'd6182;
      71523:data<=-16'd6639;
      71524:data<=-16'd8129;
      71525:data<=-16'd8621;
      71526:data<=-16'd8466;
      71527:data<=-16'd7805;
      71528:data<=-16'd6731;
      71529:data<=-16'd6852;
      71530:data<=-16'd7965;
      71531:data<=-16'd8204;
      71532:data<=-16'd7727;
      71533:data<=-16'd8402;
      71534:data<=-16'd8918;
      71535:data<=-16'd7533;
      71536:data<=-16'd7442;
      71537:data<=-16'd8752;
      71538:data<=-16'd8223;
      71539:data<=-16'd8072;
      71540:data<=-16'd8859;
      71541:data<=-16'd7908;
      71542:data<=-16'd7558;
      71543:data<=-16'd8837;
      71544:data<=-16'd8837;
      71545:data<=-16'd8006;
      71546:data<=-16'd7746;
      71547:data<=-16'd7316;
      71548:data<=-16'd7316;
      71549:data<=-16'd8789;
      71550:data<=-16'd10563;
      71551:data<=-16'd11612;
      71552:data<=-16'd11826;
      71553:data<=-16'd10942;
      71554:data<=-16'd10266;
      71555:data<=-16'd10598;
      71556:data<=-16'd10866;
      71557:data<=-16'd11294;
      71558:data<=-16'd11107;
      71559:data<=-16'd9326;
      71560:data<=-16'd8361;
      71561:data<=-16'd8231;
      71562:data<=-16'd6924;
      71563:data<=-16'd6043;
      71564:data<=-16'd6075;
      71565:data<=-16'd5465;
      71566:data<=-16'd5148;
      71567:data<=-16'd5212;
      71568:data<=-16'd3729;
      71569:data<=-16'd2343;
      71570:data<=-16'd2968;
      71571:data<=-16'd2329;
      71572:data<=-16'd698;
      71573:data<=-16'd1585;
      71574:data<=-16'd1162;
      71575:data<=16'd1492;
      71576:data<=16'd1527;
      71577:data<=16'd1386;
      71578:data<=16'd1894;
      71579:data<=16'd766;
      71580:data<=16'd2329;
      71581:data<=16'd4499;
      71582:data<=16'd2770;
      71583:data<=16'd3751;
      71584:data<=16'd7934;
      71585:data<=16'd8834;
      71586:data<=16'd8658;
      71587:data<=16'd9303;
      71588:data<=16'd8611;
      71589:data<=16'd8160;
      71590:data<=16'd8599;
      71591:data<=16'd8026;
      71592:data<=16'd7298;
      71593:data<=16'd8205;
      71594:data<=16'd9912;
      71595:data<=16'd10756;
      71596:data<=16'd10575;
      71597:data<=16'd9984;
      71598:data<=16'd9696;
      71599:data<=16'd10096;
      71600:data<=16'd10119;
      71601:data<=16'd9388;
      71602:data<=16'd9638;
      71603:data<=16'd10288;
      71604:data<=16'd9427;
      71605:data<=16'd9600;
      71606:data<=16'd11267;
      71607:data<=16'd10147;
      71608:data<=16'd8853;
      71609:data<=16'd10551;
      71610:data<=16'd10480;
      71611:data<=16'd9777;
      71612:data<=16'd11285;
      71613:data<=16'd10402;
      71614:data<=16'd9145;
      71615:data<=16'd10378;
      71616:data<=16'd8986;
      71617:data<=16'd6557;
      71618:data<=16'd6596;
      71619:data<=16'd6126;
      71620:data<=16'd5618;
      71621:data<=16'd6475;
      71622:data<=16'd6608;
      71623:data<=16'd5623;
      71624:data<=16'd5542;
      71625:data<=16'd7030;
      71626:data<=16'd7394;
      71627:data<=16'd7282;
      71628:data<=16'd8349;
      71629:data<=16'd6699;
      71630:data<=16'd5309;
      71631:data<=16'd8088;
      71632:data<=16'd8536;
      71633:data<=16'd7809;
      71634:data<=16'd8771;
      71635:data<=16'd6602;
      71636:data<=16'd6175;
      71637:data<=16'd9022;
      71638:data<=16'd7843;
      71639:data<=16'd6246;
      71640:data<=16'd6269;
      71641:data<=16'd5216;
      71642:data<=16'd6166;
      71643:data<=16'd7097;
      71644:data<=16'd6228;
      71645:data<=16'd6337;
      71646:data<=16'd5962;
      71647:data<=16'd5753;
      71648:data<=16'd6050;
      71649:data<=16'd5709;
      71650:data<=16'd8066;
      71651:data<=16'd10831;
      71652:data<=16'd10584;
      71653:data<=16'd10431;
      71654:data<=16'd10097;
      71655:data<=16'd9583;
      71656:data<=16'd10301;
      71657:data<=16'd9774;
      71658:data<=16'd8715;
      71659:data<=16'd9010;
      71660:data<=16'd9347;
      71661:data<=16'd8757;
      71662:data<=16'd7321;
      71663:data<=16'd6874;
      71664:data<=16'd7294;
      71665:data<=16'd6551;
      71666:data<=16'd5729;
      71667:data<=16'd4999;
      71668:data<=16'd3215;
      71669:data<=16'd820;
      71670:data<=-16'd180;
      71671:data<=16'd1850;
      71672:data<=16'd3048;
      71673:data<=16'd2080;
      71674:data<=16'd1572;
      71675:data<=-16'd817;
      71676:data<=-16'd1713;
      71677:data<=16'd640;
      71678:data<=-16'd790;
      71679:data<=-16'd975;
      71680:data<=16'd879;
      71681:data<=-16'd2525;
      71682:data<=-16'd3;
      71683:data<=16'd8719;
      71684:data<=16'd8921;
      71685:data<=16'd6482;
      71686:data<=16'd6998;
      71687:data<=16'd6373;
      71688:data<=16'd5594;
      71689:data<=16'd3338;
      71690:data<=16'd1789;
      71691:data<=16'd2341;
      71692:data<=16'd1105;
      71693:data<=16'd672;
      71694:data<=-16'd1759;
      71695:data<=-16'd6889;
      71696:data<=-16'd7579;
      71697:data<=-16'd12157;
      71698:data<=-16'd21105;
      71699:data<=-16'd21575;
      71700:data<=-16'd20271;
      71701:data<=-16'd21470;
      71702:data<=-16'd19863;
      71703:data<=-16'd19843;
      71704:data<=-16'd19943;
      71705:data<=-16'd16299;
      71706:data<=-16'd8769;
      71707:data<=16'd140;
      71708:data<=-16'd6032;
      71709:data<=-16'd24275;
      71710:data<=-16'd28617;
      71711:data<=-16'd23511;
      71712:data<=-16'd23914;
      71713:data<=-16'd24295;
      71714:data<=-16'd23344;
      71715:data<=-16'd22568;
      71716:data<=-16'd21549;
      71717:data<=-16'd22754;
      71718:data<=-16'd21655;
      71719:data<=-16'd18534;
      71720:data<=-16'd18252;
      71721:data<=-16'd14997;
      71722:data<=-16'd10633;
      71723:data<=-16'd14248;
      71724:data<=-16'd17687;
      71725:data<=-16'd8355;
      71726:data<=16'd7094;
      71727:data<=16'd12753;
      71728:data<=16'd8266;
      71729:data<=16'd5454;
      71730:data<=16'd7712;
      71731:data<=16'd9612;
      71732:data<=16'd6075;
      71733:data<=16'd2834;
      71734:data<=16'd9066;
      71735:data<=16'd13908;
      71736:data<=16'd8345;
      71737:data<=16'd5060;
      71738:data<=16'd9840;
      71739:data<=16'd18463;
      71740:data<=16'd23892;
      71741:data<=16'd17729;
      71742:data<=16'd7987;
      71743:data<=16'd3286;
      71744:data<=16'd2784;
      71745:data<=16'd8893;
      71746:data<=16'd13491;
      71747:data<=16'd10302;
      71748:data<=16'd5532;
      71749:data<=16'd2403;
      71750:data<=16'd7970;
      71751:data<=16'd12848;
      71752:data<=16'd4052;
      71753:data<=16'd3721;
      71754:data<=16'd11405;
      71755:data<=16'd7620;
      71756:data<=16'd8722;
      71757:data<=16'd13030;
      71758:data<=16'd6796;
      71759:data<=16'd5163;
      71760:data<=16'd9059;
      71761:data<=16'd8469;
      71762:data<=-16'd1689;
      71763:data<=-16'd17690;
      71764:data<=-16'd19907;
      71765:data<=-16'd17473;
      71766:data<=-16'd20445;
      71767:data<=-16'd13179;
      71768:data<=-16'd11079;
      71769:data<=-16'd16487;
      71770:data<=-16'd11523;
      71771:data<=-16'd12916;
      71772:data<=-16'd12440;
      71773:data<=-16'd1353;
      71774:data<=-16'd7350;
      71775:data<=-16'd16172;
      71776:data<=-16'd13242;
      71777:data<=-16'd12739;
      71778:data<=-16'd7990;
      71779:data<=-16'd6790;
      71780:data<=-16'd8874;
      71781:data<=-16'd305;
      71782:data<=-16'd5145;
      71783:data<=-16'd17728;
      71784:data<=-16'd14762;
      71785:data<=-16'd15399;
      71786:data<=-16'd16310;
      71787:data<=-16'd12404;
      71788:data<=-16'd17738;
      71789:data<=-16'd14355;
      71790:data<=-16'd5841;
      71791:data<=-16'd10111;
      71792:data<=-16'd8047;
      71793:data<=-16'd2675;
      71794:data<=-16'd8228;
      71795:data<=-16'd12123;
      71796:data<=-16'd10834;
      71797:data<=-16'd7915;
      71798:data<=-16'd8628;
      71799:data<=-16'd11209;
      71800:data<=-16'd378;
      71801:data<=16'd8549;
      71802:data<=16'd1184;
      71803:data<=16'd385;
      71804:data<=16'd6704;
      71805:data<=16'd8231;
      71806:data<=16'd10094;
      71807:data<=16'd7095;
      71808:data<=16'd2109;
      71809:data<=16'd1485;
      71810:data<=-16'd3797;
      71811:data<=-16'd5356;
      71812:data<=16'd2340;
      71813:data<=16'd5086;
      71814:data<=16'd2913;
      71815:data<=-16'd332;
      71816:data<=-16'd1134;
      71817:data<=16'd2946;
      71818:data<=16'd223;
      71819:data<=-16'd405;
      71820:data<=16'd8654;
      71821:data<=16'd4708;
      71822:data<=-16'd2118;
      71823:data<=16'd3955;
      71824:data<=16'd2127;
      71825:data<=16'd183;
      71826:data<=16'd8516;
      71827:data<=16'd7274;
      71828:data<=16'd2895;
      71829:data<=16'd3007;
      71830:data<=16'd1697;
      71831:data<=16'd8052;
      71832:data<=16'd12325;
      71833:data<=16'd6516;
      71834:data<=16'd5792;
      71835:data<=16'd6187;
      71836:data<=16'd6611;
      71837:data<=16'd8507;
      71838:data<=-16'd2604;
      71839:data<=-16'd10957;
      71840:data<=-16'd5874;
      71841:data<=-16'd9585;
      71842:data<=-16'd14049;
      71843:data<=-16'd9636;
      71844:data<=-16'd10496;
      71845:data<=-16'd9445;
      71846:data<=-16'd4905;
      71847:data<=-16'd8200;
      71848:data<=-16'd11732;
      71849:data<=-16'd12351;
      71850:data<=-16'd11705;
      71851:data<=-16'd5485;
      71852:data<=16'd114;
      71853:data<=-16'd1064;
      71854:data<=-16'd5422;
      71855:data<=-16'd5567;
      71856:data<=-16'd1240;
      71857:data<=-16'd2620;
      71858:data<=-16'd6402;
      71859:data<=-16'd6319;
      71860:data<=-16'd9400;
      71861:data<=-16'd9649;
      71862:data<=-16'd3612;
      71863:data<=-16'd3001;
      71864:data<=-16'd4353;
      71865:data<=-16'd2268;
      71866:data<=-16'd1168;
      71867:data<=-16'd2029;
      71868:data<=-16'd5157;
      71869:data<=-16'd5433;
      71870:data<=-16'd3162;
      71871:data<=-16'd5912;
      71872:data<=-16'd7644;
      71873:data<=-16'd9356;
      71874:data<=-16'd15609;
      71875:data<=-16'd10346;
      71876:data<=16'd5036;
      71877:data<=16'd8890;
      71878:data<=16'd4353;
      71879:data<=16'd6807;
      71880:data<=16'd12299;
      71881:data<=16'd11036;
      71882:data<=16'd7847;
      71883:data<=16'd3767;
      71884:data<=-16'd4279;
      71885:data<=-16'd2118;
      71886:data<=16'd6079;
      71887:data<=16'd2308;
      71888:data<=16'd993;
      71889:data<=16'd4863;
      71890:data<=16'd1354;
      71891:data<=16'd5028;
      71892:data<=16'd10592;
      71893:data<=16'd1736;
      71894:data<=-16'd2673;
      71895:data<=16'd1287;
      71896:data<=-16'd2766;
      71897:data<=-16'd5876;
      71898:data<=16'd1212;
      71899:data<=16'd3413;
      71900:data<=-16'd2508;
      71901:data<=16'd1387;
      71902:data<=16'd8147;
      71903:data<=16'd3109;
      71904:data<=16'd2097;
      71905:data<=16'd4666;
      71906:data<=16'd1374;
      71907:data<=16'd6097;
      71908:data<=16'd8184;
      71909:data<=-16'd1387;
      71910:data<=16'd384;
      71911:data<=16'd7943;
      71912:data<=16'd2787;
      71913:data<=-16'd7699;
      71914:data<=-16'd13715;
      71915:data<=-16'd14707;
      71916:data<=-16'd15044;
      71917:data<=-16'd9479;
      71918:data<=-16'd205;
      71919:data<=-16'd3694;
      71920:data<=-16'd4868;
      71921:data<=16'd3920;
      71922:data<=-16'd118;
      71923:data<=-16'd3234;
      71924:data<=16'd5802;
      71925:data<=16'd5601;
      71926:data<=-16'd619;
      71927:data<=-16'd3146;
      71928:data<=-16'd2253;
      71929:data<=16'd2146;
      71930:data<=16'd958;
      71931:data<=-16'd262;
      71932:data<=16'd5723;
      71933:data<=16'd5797;
      71934:data<=16'd406;
      71935:data<=16'd1104;
      71936:data<=16'd4887;
      71937:data<=16'd1042;
      71938:data<=-16'd3497;
      71939:data<=16'd4582;
      71940:data<=16'd5817;
      71941:data<=-16'd3556;
      71942:data<=16'd2796;
      71943:data<=16'd8164;
      71944:data<=16'd1107;
      71945:data<=16'd2643;
      71946:data<=16'd2237;
      71947:data<=-16'd361;
      71948:data<=16'd6346;
      71949:data<=16'd7192;
      71950:data<=16'd10555;
      71951:data<=16'd21983;
      71952:data<=16'd24109;
      71953:data<=16'd25297;
      71954:data<=16'd25539;
      71955:data<=16'd18022;
      71956:data<=16'd17429;
      71957:data<=16'd18298;
      71958:data<=16'd13928;
      71959:data<=16'd17252;
      71960:data<=16'd23115;
      71961:data<=16'd20219;
      71962:data<=16'd13747;
      71963:data<=16'd11074;
      71964:data<=16'd8757;
      71965:data<=16'd5291;
      71966:data<=16'd7567;
      71967:data<=16'd8545;
      71968:data<=16'd5627;
      71969:data<=16'd7874;
      71970:data<=16'd6784;
      71971:data<=16'd6616;
      71972:data<=16'd10922;
      71973:data<=16'd1105;
      71974:data<=-16'd2989;
      71975:data<=16'd8668;
      71976:data<=16'd6569;
      71977:data<=16'd4654;
      71978:data<=16'd10472;
      71979:data<=16'd5177;
      71980:data<=16'd4931;
      71981:data<=16'd6138;
      71982:data<=16'd6;
      71983:data<=16'd4067;
      71984:data<=16'd3729;
      71985:data<=16'd942;
      71986:data<=16'd11630;
      71987:data<=16'd6346;
      71988:data<=-16'd10346;
      71989:data<=-16'd11952;
      71990:data<=-16'd13426;
      71991:data<=-16'd14821;
      71992:data<=-16'd10847;
      71993:data<=-16'd11873;
      71994:data<=-16'd10138;
      71995:data<=-16'd5727;
      71996:data<=-16'd6687;
      71997:data<=-16'd5468;
      71998:data<=-16'd2651;
      71999:data<=-16'd5332;
      72000:data<=-16'd6531;
      72001:data<=16'd437;
      72002:data<=16'd1503;
      72003:data<=-16'd6443;
      72004:data<=-16'd3905;
      72005:data<=-16'd1762;
      72006:data<=-16'd7403;
      72007:data<=16'd2593;
      72008:data<=16'd9527;
      72009:data<=16'd144;
      72010:data<=16'd4256;
      72011:data<=16'd9723;
      72012:data<=16'd2221;
      72013:data<=16'd1155;
      72014:data<=16'd1105;
      72015:data<=-16'd1104;
      72016:data<=16'd170;
      72017:data<=-16'd1392;
      72018:data<=16'd2438;
      72019:data<=16'd9094;
      72020:data<=16'd4963;
      72021:data<=16'd455;
      72022:data<=16'd2040;
      72023:data<=16'd3013;
      72024:data<=16'd4347;
      72025:data<=16'd12292;
      72026:data<=16'd22571;
      72027:data<=16'd20768;
      72028:data<=16'd15206;
      72029:data<=16'd19549;
      72030:data<=16'd19746;
      72031:data<=16'd14801;
      72032:data<=16'd17744;
      72033:data<=16'd20046;
      72034:data<=16'd14410;
      72035:data<=16'd9981;
      72036:data<=16'd12616;
      72037:data<=16'd14222;
      72038:data<=16'd12046;
      72039:data<=16'd14390;
      72040:data<=16'd13728;
      72041:data<=16'd8727;
      72042:data<=16'd12725;
      72043:data<=16'd13869;
      72044:data<=16'd6407;
      72045:data<=16'd5729;
      72046:data<=16'd7840;
      72047:data<=16'd6072;
      72048:data<=16'd4109;
      72049:data<=16'd4212;
      72050:data<=16'd5588;
      72051:data<=16'd2070;
      72052:data<=-16'd372;
      72053:data<=16'd793;
      72054:data<=-16'd5009;
      72055:data<=-16'd5341;
      72056:data<=16'd3362;
      72057:data<=16'd1521;
      72058:data<=-16'd4364;
      72059:data<=-16'd3565;
      72060:data<=-16'd1647;
      72061:data<=16'd133;
      72062:data<=-16'd963;
      72063:data<=-16'd7185;
      72064:data<=-16'd14662;
      72065:data<=-16'd18072;
      72066:data<=-16'd20325;
      72067:data<=-16'd26024;
      72068:data<=-16'd20583;
      72069:data<=-16'd8423;
      72070:data<=-16'd13238;
      72071:data<=-16'd19161;
      72072:data<=-16'd13562;
      72073:data<=-16'd11247;
      72074:data<=-16'd9165;
      72075:data<=-16'd6050;
      72076:data<=-16'd6411;
      72077:data<=-16'd9241;
      72078:data<=-16'd15499;
      72079:data<=-16'd13060;
      72080:data<=-16'd5488;
      72081:data<=-16'd7823;
      72082:data<=-16'd8530;
      72083:data<=-16'd8185;
      72084:data<=-16'd10419;
      72085:data<=-16'd4455;
      72086:data<=-16'd4552;
      72087:data<=-16'd11984;
      72088:data<=-16'd7612;
      72089:data<=-16'd2196;
      72090:data<=-16'd5858;
      72091:data<=-16'd8005;
      72092:data<=-16'd4666;
      72093:data<=-16'd4557;
      72094:data<=-16'd8275;
      72095:data<=-16'd2290;
      72096:data<=16'd4546;
      72097:data<=16'd2432;
      72098:data<=16'd5985;
      72099:data<=16'd7777;
      72100:data<=16'd6693;
      72101:data<=16'd16324;
      72102:data<=16'd19385;
      72103:data<=16'd19546;
      72104:data<=16'd25543;
      72105:data<=16'd16666;
      72106:data<=16'd10743;
      72107:data<=16'd17673;
      72108:data<=16'd13364;
      72109:data<=16'd11291;
      72110:data<=16'd14625;
      72111:data<=16'd10170;
      72112:data<=16'd12439;
      72113:data<=16'd14889;
      72114:data<=16'd9777;
      72115:data<=16'd10630;
      72116:data<=16'd10803;
      72117:data<=16'd9630;
      72118:data<=16'd13123;
      72119:data<=16'd10292;
      72120:data<=16'd4487;
      72121:data<=16'd5447;
      72122:data<=16'd7024;
      72123:data<=16'd4026;
      72124:data<=16'd1791;
      72125:data<=16'd4273;
      72126:data<=16'd3448;
      72127:data<=16'd1483;
      72128:data<=16'd7097;
      72129:data<=16'd6461;
      72130:data<=-16'd65;
      72131:data<=16'd4587;
      72132:data<=16'd6031;
      72133:data<=-16'd4096;
      72134:data<=-16'd6240;
      72135:data<=-16'd1004;
      72136:data<=-16'd1025;
      72137:data<=-16'd5031;
      72138:data<=-16'd11729;
      72139:data<=-16'd20286;
      72140:data<=-16'd23739;
      72141:data<=-16'd21055;
      72142:data<=-16'd19869;
      72143:data<=-16'd21675;
      72144:data<=-16'd21978;
      72145:data<=-16'd21614;
      72146:data<=-16'd23003;
      72147:data<=-16'd24278;
      72148:data<=-16'd22005;
      72149:data<=-16'd19707;
      72150:data<=-16'd23892;
      72151:data<=-16'd24799;
      72152:data<=-16'd15506;
      72153:data<=-16'd12486;
      72154:data<=-16'd17687;
      72155:data<=-16'd16013;
      72156:data<=-16'd12856;
      72157:data<=-16'd15161;
      72158:data<=-16'd14002;
      72159:data<=-16'd10722;
      72160:data<=-16'd14455;
      72161:data<=-16'd20424;
      72162:data<=-16'd21526;
      72163:data<=-16'd20318;
      72164:data<=-16'd15549;
      72165:data<=-16'd8387;
      72166:data<=-16'd9429;
      72167:data<=-16'd14598;
      72168:data<=-16'd14662;
      72169:data<=-16'd13947;
      72170:data<=-16'd11761;
      72171:data<=-16'd8928;
      72172:data<=-16'd9620;
      72173:data<=-16'd8141;
      72174:data<=-16'd8652;
      72175:data<=-16'd10031;
      72176:data<=-16'd5;
      72177:data<=16'd6438;
      72178:data<=16'd2406;
      72179:data<=16'd5720;
      72180:data<=16'd9068;
      72181:data<=16'd4561;
      72182:data<=16'd2638;
      72183:data<=16'd2641;
      72184:data<=16'd5788;
      72185:data<=16'd12947;
      72186:data<=16'd13382;
      72187:data<=16'd7464;
      72188:data<=16'd6404;
      72189:data<=16'd12722;
      72190:data<=16'd15013;
      72191:data<=16'd11160;
      72192:data<=16'd11946;
      72193:data<=16'd8536;
      72194:data<=16'd1004;
      72195:data<=16'd6874;
      72196:data<=16'd9737;
      72197:data<=16'd1698;
      72198:data<=16'd3474;
      72199:data<=16'd7188;
      72200:data<=16'd4404;
      72201:data<=16'd3808;
      72202:data<=16'd5092;
      72203:data<=16'd8984;
      72204:data<=16'd8713;
      72205:data<=16'd3419;
      72206:data<=16'd4191;
      72207:data<=16'd4484;
      72208:data<=16'd4214;
      72209:data<=16'd2426;
      72210:data<=-16'd5571;
      72211:data<=16'd1694;
      72212:data<=16'd7206;
      72213:data<=-16'd11869;
      72214:data<=-16'd15238;
      72215:data<=-16'd8040;
      72216:data<=-16'd16801;
      72217:data<=-16'd13876;
      72218:data<=-16'd9638;
      72219:data<=-16'd16057;
      72220:data<=-16'd8992;
      72221:data<=-16'd5944;
      72222:data<=-16'd11697;
      72223:data<=-16'd9882;
      72224:data<=-16'd13756;
      72225:data<=-16'd17341;
      72226:data<=-16'd14883;
      72227:data<=-16'd14859;
      72228:data<=-16'd10878;
      72229:data<=-16'd12461;
      72230:data<=-16'd16548;
      72231:data<=-16'd12120;
      72232:data<=-16'd18369;
      72233:data<=-16'd22501;
      72234:data<=-16'd11744;
      72235:data<=-16'd12245;
      72236:data<=-16'd14392;
      72237:data<=-16'd10366;
      72238:data<=-16'd16797;
      72239:data<=-16'd18694;
      72240:data<=-16'd14092;
      72241:data<=-16'd15079;
      72242:data<=-16'd12686;
      72243:data<=-16'd10848;
      72244:data<=-16'd10008;
      72245:data<=-16'd5397;
      72246:data<=-16'd7360;
      72247:data<=-16'd8621;
      72248:data<=-16'd6511;
      72249:data<=-16'd9477;
      72250:data<=-16'd2300;
      72251:data<=16'd10762;
      72252:data<=16'd11779;
      72253:data<=16'd10906;
      72254:data<=16'd8765;
      72255:data<=16'd5063;
      72256:data<=16'd10604;
      72257:data<=16'd11429;
      72258:data<=16'd5406;
      72259:data<=16'd7427;
      72260:data<=16'd8028;
      72261:data<=16'd7759;
      72262:data<=16'd12217;
      72263:data<=16'd7456;
      72264:data<=16'd1504;
      72265:data<=16'd4660;
      72266:data<=16'd6402;
      72267:data<=16'd9054;
      72268:data<=16'd9788;
      72269:data<=16'd4561;
      72270:data<=16'd7056;
      72271:data<=16'd8208;
      72272:data<=16'd795;
      72273:data<=16'd4825;
      72274:data<=16'd12972;
      72275:data<=16'd10493;
      72276:data<=16'd10082;
      72277:data<=16'd11853;
      72278:data<=16'd6837;
      72279:data<=16'd2884;
      72280:data<=16'd7307;
      72281:data<=16'd12722;
      72282:data<=16'd9837;
      72283:data<=16'd6848;
      72284:data<=16'd9740;
      72285:data<=16'd6878;
      72286:data<=16'd2103;
      72287:data<=16'd2907;
      72288:data<=-16'd1510;
      72289:data<=-16'd5832;
      72290:data<=-16'd2833;
      72291:data<=-16'd5729;
      72292:data<=-16'd11397;
      72293:data<=-16'd11285;
      72294:data<=-16'd11890;
      72295:data<=-16'd10690;
      72296:data<=-16'd8288;
      72297:data<=-16'd9041;
      72298:data<=-16'd3036;
      72299:data<=16'd2566;
      72300:data<=-16'd4868;
      72301:data<=-16'd9461;
      72302:data<=-16'd5092;
      72303:data<=-16'd2393;
      72304:data<=-16'd2056;
      72305:data<=-16'd4974;
      72306:data<=-16'd7820;
      72307:data<=-16'd7915;
      72308:data<=-16'd9444;
      72309:data<=-16'd4021;
      72310:data<=16'd3016;
      72311:data<=-16'd3272;
      72312:data<=-16'd6673;
      72313:data<=-16'd1054;
      72314:data<=-16'd159;
      72315:data<=-16'd121;
      72316:data<=16'd291;
      72317:data<=-16'd490;
      72318:data<=-16'd1403;
      72319:data<=-16'd7488;
      72320:data<=-16'd10463;
      72321:data<=-16'd8715;
      72322:data<=-16'd9638;
      72323:data<=-16'd6687;
      72324:data<=-16'd5517;
      72325:data<=-16'd3166;
      72326:data<=16'd11929;
      72327:data<=16'd17261;
      72328:data<=16'd11122;
      72329:data<=16'd12713;
      72330:data<=16'd12733;
      72331:data<=16'd13928;
      72332:data<=16'd16610;
      72333:data<=16'd10621;
      72334:data<=16'd11767;
      72335:data<=16'd13761;
      72336:data<=16'd6945;
      72337:data<=16'd12069;
      72338:data<=16'd17708;
      72339:data<=16'd12527;
      72340:data<=16'd13086;
      72341:data<=16'd12992;
      72342:data<=16'd9919;
      72343:data<=16'd11408;
      72344:data<=16'd11075;
      72345:data<=16'd9922;
      72346:data<=16'd7774;
      72347:data<=16'd6987;
      72348:data<=16'd10836;
      72349:data<=16'd6170;
      72350:data<=16'd2770;
      72351:data<=16'd11088;
      72352:data<=16'd9163;
      72353:data<=16'd3654;
      72354:data<=16'd9060;
      72355:data<=16'd8581;
      72356:data<=16'd6166;
      72357:data<=16'd11661;
      72358:data<=16'd12642;
      72359:data<=16'd8348;
      72360:data<=16'd6176;
      72361:data<=16'd10052;
      72362:data<=16'd15802;
      72363:data<=16'd9021;
      72364:data<=-16'd687;
      72365:data<=16'd2452;
      72366:data<=16'd3198;
      72367:data<=-16'd3110;
      72368:data<=-16'd4323;
      72369:data<=-16'd4361;
      72370:data<=-16'd3941;
      72371:data<=-16'd701;
      72372:data<=16'd320;
      72373:data<=16'd2416;
      72374:data<=16'd4514;
      72375:data<=16'd3015;
      72376:data<=16'd3007;
      72377:data<=-16'd638;
      72378:data<=-16'd7764;
      72379:data<=-16'd6426;
      72380:data<=16'd597;
      72381:data<=16'd6217;
      72382:data<=16'd4884;
      72383:data<=-16'd1644;
      72384:data<=16'd925;
      72385:data<=16'd5022;
      72386:data<=16'd1903;
      72387:data<=16'd2931;
      72388:data<=16'd1421;
      72389:data<=-16'd467;
      72390:data<=16'd8002;
      72391:data<=16'd7191;
      72392:data<=16'd1113;
      72393:data<=16'd7500;
      72394:data<=16'd8781;
      72395:data<=16'd4141;
      72396:data<=16'd4948;
      72397:data<=16'd1613;
      72398:data<=-16'd3980;
      72399:data<=-16'd2234;
      72400:data<=16'd7110;
      72401:data<=16'd15940;
      72402:data<=16'd17241;
      72403:data<=16'd18921;
      72404:data<=16'd18883;
      72405:data<=16'd14328;
      72406:data<=16'd17916;
      72407:data<=16'd18406;
      72408:data<=16'd9445;
      72409:data<=16'd7729;
      72410:data<=16'd6370;
      72411:data<=16'd4067;
      72412:data<=16'd8254;
      72413:data<=16'd5715;
      72414:data<=16'd3254;
      72415:data<=16'd8225;
      72416:data<=16'd4217;
      72417:data<=-16'd1406;
      72418:data<=16'd2875;
      72419:data<=16'd6234;
      72420:data<=16'd3788;
      72421:data<=16'd364;
      72422:data<=16'd3629;
      72423:data<=16'd10354;
      72424:data<=16'd8522;
      72425:data<=16'd4599;
      72426:data<=16'd5362;
      72427:data<=16'd5550;
      72428:data<=16'd6992;
      72429:data<=16'd7116;
      72430:data<=16'd3835;
      72431:data<=16'd4645;
      72432:data<=16'd4071;
      72433:data<=-16'd390;
      72434:data<=16'd846;
      72435:data<=16'd1444;
      72436:data<=-16'd2;
      72437:data<=16'd4804;
      72438:data<=16'd1835;
      72439:data<=-16'd10599;
      72440:data<=-16'd13088;
      72441:data<=-16'd10467;
      72442:data<=-16'd9750;
      72443:data<=-16'd8672;
      72444:data<=-16'd12278;
      72445:data<=-16'd11612;
      72446:data<=-16'd8698;
      72447:data<=-16'd16421;
      72448:data<=-16'd14395;
      72449:data<=-16'd2467;
      72450:data<=-16'd5072;
      72451:data<=-16'd7253;
      72452:data<=-16'd70;
      72453:data<=16'd1961;
      72454:data<=16'd1356;
      72455:data<=16'd2135;
      72456:data<=16'd5336;
      72457:data<=16'd5153;
      72458:data<=-16'd2497;
      72459:data<=16'd343;
      72460:data<=16'd7059;
      72461:data<=16'd240;
      72462:data<=-16'd2464;
      72463:data<=16'd1240;
      72464:data<=-16'd5;
      72465:data<=-16'd214;
      72466:data<=16'd153;
      72467:data<=16'd1262;
      72468:data<=16'd1348;
      72469:data<=-16'd2769;
      72470:data<=-16'd1794;
      72471:data<=16'd588;
      72472:data<=16'd2567;
      72473:data<=16'd5934;
      72474:data<=-16'd325;
      72475:data<=16'd1676;
      72476:data<=16'd16933;
      72477:data<=16'd15526;
      72478:data<=16'd12108;
      72479:data<=16'd19440;
      72480:data<=16'd16031;
      72481:data<=16'd10398;
      72482:data<=16'd9577;
      72483:data<=16'd8511;
      72484:data<=16'd11326;
      72485:data<=16'd9896;
      72486:data<=16'd10731;
      72487:data<=16'd17285;
      72488:data<=16'd10921;
      72489:data<=16'd4811;
      72490:data<=16'd7471;
      72491:data<=16'd3192;
      72492:data<=16'd3600;
      72493:data<=16'd12343;
      72494:data<=16'd14539;
      72495:data<=16'd10760;
      72496:data<=16'd3298;
      72497:data<=-16'd616;
      72498:data<=16'd2461;
      72499:data<=16'd2998;
      72500:data<=16'd1973;
      72501:data<=-16'd1342;
      72502:data<=-16'd5607;
      72503:data<=-16'd1263;
      72504:data<=16'd852;
      72505:data<=-16'd2966;
      72506:data<=-16'd808;
      72507:data<=-16'd302;
      72508:data<=-16'd3303;
      72509:data<=-16'd4275;
      72510:data<=-16'd10132;
      72511:data<=-16'd11353;
      72512:data<=-16'd2370;
      72513:data<=-16'd4711;
      72514:data<=-16'd16678;
      72515:data<=-16'd17220;
      72516:data<=-16'd14051;
      72517:data<=-16'd17007;
      72518:data<=-16'd14357;
      72519:data<=-16'd11192;
      72520:data<=-16'd19279;
      72521:data<=-16'd21567;
      72522:data<=-16'd13050;
      72523:data<=-16'd13386;
      72524:data<=-16'd18918;
      72525:data<=-16'd18160;
      72526:data<=-16'd16830;
      72527:data<=-16'd17191;
      72528:data<=-16'd18648;
      72529:data<=-16'd19199;
      72530:data<=-16'd16433;
      72531:data<=-16'd16551;
      72532:data<=-16'd15079;
      72533:data<=-16'd7310;
      72534:data<=-16'd7473;
      72535:data<=-16'd13074;
      72536:data<=-16'd12007;
      72537:data<=-16'd12342;
      72538:data<=-16'd13135;
      72539:data<=-16'd9256;
      72540:data<=-16'd10213;
      72541:data<=-16'd8880;
      72542:data<=16'd1644;
      72543:data<=16'd3334;
      72544:data<=-16'd2719;
      72545:data<=-16'd1392;
      72546:data<=-16'd1105;
      72547:data<=-16'd4375;
      72548:data<=-16'd3266;
      72549:data<=-16'd3424;
      72550:data<=16'd21;
      72551:data<=16'd12169;
      72552:data<=16'd15675;
      72553:data<=16'd10531;
      72554:data<=16'd10060;
      72555:data<=16'd10131;
      72556:data<=16'd10693;
      72557:data<=16'd11667;
      72558:data<=16'd9758;
      72559:data<=16'd13920;
      72560:data<=16'd15499;
      72561:data<=16'd5742;
      72562:data<=16'd5372;
      72563:data<=16'd10128;
      72564:data<=16'd3063;
      72565:data<=16'd966;
      72566:data<=16'd6385;
      72567:data<=16'd5100;
      72568:data<=16'd4598;
      72569:data<=16'd7139;
      72570:data<=16'd5280;
      72571:data<=16'd3039;
      72572:data<=16'd3482;
      72573:data<=16'd2975;
      72574:data<=16'd587;
      72575:data<=-16'd118;
      72576:data<=16'd303;
      72577:data<=-16'd1394;
      72578:data<=-16'd2349;
      72579:data<=-16'd4284;
      72580:data<=-16'd6657;
      72581:data<=-16'd708;
      72582:data<=16'd4349;
      72583:data<=16'd1225;
      72584:data<=16'd1002;
      72585:data<=-16'd1202;
      72586:data<=-16'd6769;
      72587:data<=-16'd5371;
      72588:data<=-16'd11759;
      72589:data<=-16'd27445;
      72590:data<=-16'd27661;
      72591:data<=-16'd20845;
      72592:data<=-16'd24501;
      72593:data<=-16'd24215;
      72594:data<=-16'd18199;
      72595:data<=-16'd23296;
      72596:data<=-16'd27038;
      72597:data<=-16'd15834;
      72598:data<=-16'd13888;
      72599:data<=-16'd24447;
      72600:data<=-16'd21984;
      72601:data<=-16'd18964;
      72602:data<=-16'd25276;
      72603:data<=-16'd18823;
      72604:data<=-16'd10428;
      72605:data<=-16'd13961;
      72606:data<=-16'd13849;
      72607:data<=-16'd14113;
      72608:data<=-16'd14601;
      72609:data<=-16'd6419;
      72610:data<=-16'd8020;
      72611:data<=-16'd15517;
      72612:data<=-16'd10293;
      72613:data<=-16'd8220;
      72614:data<=-16'd12630;
      72615:data<=-16'd9843;
      72616:data<=-16'd5891;
      72617:data<=-16'd6858;
      72618:data<=-16'd10185;
      72619:data<=-16'd8522;
      72620:data<=-16'd4761;
      72621:data<=-16'd11620;
      72622:data<=-16'd12696;
      72623:data<=-16'd2288;
      72624:data<=-16'd4592;
      72625:data<=-16'd4960;
      72626:data<=16'd8637;
      72627:data<=16'd13571;
      72628:data<=16'd13526;
      72629:data<=16'd11831;
      72630:data<=16'd7022;
      72631:data<=16'd14178;
      72632:data<=16'd19552;
      72633:data<=16'd17638;
      72634:data<=16'd21228;
      72635:data<=16'd14728;
      72636:data<=16'd7929;
      72637:data<=16'd14498;
      72638:data<=16'd11565;
      72639:data<=16'd7098;
      72640:data<=16'd11223;
      72641:data<=16'd12422;
      72642:data<=16'd14586;
      72643:data<=16'd9700;
      72644:data<=16'd3592;
      72645:data<=16'd9677;
      72646:data<=16'd9545;
      72647:data<=16'd11204;
      72648:data<=16'd14289;
      72649:data<=16'd1497;
      72650:data<=16'd5958;
      72651:data<=16'd15338;
      72652:data<=-16'd625;
      72653:data<=16'd1676;
      72654:data<=16'd12232;
      72655:data<=16'd1895;
      72656:data<=16'd3560;
      72657:data<=16'd6373;
      72658:data<=16'd2340;
      72659:data<=16'd11765;
      72660:data<=16'd10510;
      72661:data<=16'd4323;
      72662:data<=16'd8637;
      72663:data<=16'd197;
      72664:data<=-16'd9330;
      72665:data<=-16'd11899;
      72666:data<=-16'd16463;
      72667:data<=-16'd10049;
      72668:data<=-16'd6457;
      72669:data<=-16'd10610;
      72670:data<=-16'd4661;
      72671:data<=-16'd5186;
      72672:data<=-16'd11681;
      72673:data<=-16'd7492;
      72674:data<=-16'd6968;
      72675:data<=-16'd13568;
      72676:data<=-16'd18051;
      72677:data<=-16'd17162;
      72678:data<=-16'd12701;
      72679:data<=-16'd16195;
      72680:data<=-16'd19849;
      72681:data<=-16'd13699;
      72682:data<=-16'd11086;
      72683:data<=-16'd11464;
      72684:data<=-16'd9702;
      72685:data<=-16'd10633;
      72686:data<=-16'd10947;
      72687:data<=-16'd10411;
      72688:data<=-16'd9683;
      72689:data<=-16'd9556;
      72690:data<=-16'd10743;
      72691:data<=-16'd4249;
      72692:data<=-16'd428;
      72693:data<=-16'd8008;
      72694:data<=-16'd8097;
      72695:data<=-16'd6087;
      72696:data<=-16'd8260;
      72697:data<=-16'd1586;
      72698:data<=-16'd3433;
      72699:data<=-16'd12780;
      72700:data<=-16'd3762;
      72701:data<=16'd7692;
      72702:data<=16'd11377;
      72703:data<=16'd14583;
      72704:data<=16'd9646;
      72705:data<=16'd9376;
      72706:data<=16'd16622;
      72707:data<=16'd12930;
      72708:data<=16'd10319;
      72709:data<=16'd13264;
      72710:data<=16'd10713;
      72711:data<=16'd10816;
      72712:data<=16'd11455;
      72713:data<=16'd9388;
      72714:data<=16'd9937;
      72715:data<=16'd8519;
      72716:data<=16'd11427;
      72717:data<=16'd16634;
      72718:data<=16'd12029;
      72719:data<=16'd10913;
      72720:data<=16'd14223;
      72721:data<=16'd13047;
      72722:data<=16'd16722;
      72723:data<=16'd17550;
      72724:data<=16'd13446;
      72725:data<=16'd16836;
      72726:data<=16'd16920;
      72727:data<=16'd14433;
      72728:data<=16'd16172;
      72729:data<=16'd11400;
      72730:data<=16'd11811;
      72731:data<=16'd19755;
      72732:data<=16'd14718;
      72733:data<=16'd9670;
      72734:data<=16'd13671;
      72735:data<=16'd11435;
      72736:data<=16'd12016;
      72737:data<=16'd17250;
      72738:data<=16'd7485;
      72739:data<=-16'd5513;
      72740:data<=-16'd3642;
      72741:data<=-16'd2176;
      72742:data<=-16'd7022;
      72743:data<=-16'd4249;
      72744:data<=16'd155;
      72745:data<=-16'd3748;
      72746:data<=-16'd6246;
      72747:data<=-16'd2819;
      72748:data<=-16'd961;
      72749:data<=-16'd2989;
      72750:data<=-16'd1850;
      72751:data<=16'd5285;
      72752:data<=16'd7753;
      72753:data<=16'd5090;
      72754:data<=16'd6949;
      72755:data<=16'd7138;
      72756:data<=16'd4379;
      72757:data<=16'd5836;
      72758:data<=16'd5313;
      72759:data<=16'd3102;
      72760:data<=16'd3697;
      72761:data<=16'd3262;
      72762:data<=16'd5471;
      72763:data<=16'd8222;
      72764:data<=16'd4059;
      72765:data<=-16'd244;
      72766:data<=-16'd1968;
      72767:data<=-16'd3876;
      72768:data<=-16'd3083;
      72769:data<=-16'd2546;
      72770:data<=-16'd4816;
      72771:data<=-16'd5189;
      72772:data<=-16'd2481;
      72773:data<=-16'd1281;
      72774:data<=-16'd2964;
      72775:data<=16'd1127;
      72776:data<=16'd12933;
      72777:data<=16'd19088;
      72778:data<=16'd17042;
      72779:data<=16'd15938;
      72780:data<=16'd15699;
      72781:data<=16'd14883;
      72782:data<=16'd15485;
      72783:data<=16'd14317;
      72784:data<=16'd11802;
      72785:data<=16'd12985;
      72786:data<=16'd13673;
      72787:data<=16'd11348;
      72788:data<=16'd12460;
      72789:data<=16'd13729;
      72790:data<=16'd11530;
      72791:data<=16'd12695;
      72792:data<=16'd13691;
      72793:data<=16'd9705;
      72794:data<=16'd8166;
      72795:data<=16'd9999;
      72796:data<=16'd10666;
      72797:data<=16'd9492;
      72798:data<=16'd7736;
      72799:data<=16'd8578;
      72800:data<=16'd9865;
      72801:data<=16'd8925;
      72802:data<=16'd8849;
      72803:data<=16'd8113;
      72804:data<=16'd5571;
      72805:data<=16'd5040;
      72806:data<=16'd5473;
      72807:data<=16'd4306;
      72808:data<=16'd5513;
      72809:data<=16'd12084;
      72810:data<=16'd15650;
      72811:data<=16'd13556;
      72812:data<=16'd14835;
      72813:data<=16'd11823;
      72814:data<=-16'd1145;
      72815:data<=-16'd7077;
      72816:data<=-16'd5104;
      72817:data<=-16'd4946;
      72818:data<=-16'd4020;
      72819:data<=-16'd4723;
      72820:data<=-16'd6184;
      72821:data<=-16'd4560;
      72822:data<=-16'd4874;
      72823:data<=-16'd4763;
      72824:data<=-16'd2259;
      72825:data<=-16'd2259;
      72826:data<=-16'd3040;
      72827:data<=-16'd2899;
      72828:data<=-16'd2870;
      72829:data<=-16'd4360;
      72830:data<=-16'd5859;
      72831:data<=-16'd3568;
      72832:data<=-16'd3751;
      72833:data<=-16'd7265;
      72834:data<=-16'd6479;
      72835:data<=-16'd5271;
      72836:data<=-16'd3894;
      72837:data<=-16'd1034;
      72838:data<=-16'd2153;
      72839:data<=-16'd2911;
      72840:data<=-16'd3039;
      72841:data<=-16'd4770;
      72842:data<=-16'd2748;
      72843:data<=-16'd2525;
      72844:data<=-16'd4181;
      72845:data<=-16'd1524;
      72846:data<=-16'd2000;
      72847:data<=-16'd4272;
      72848:data<=-16'd4000;
      72849:data<=-16'd4843;
      72850:data<=-16'd44;
      72851:data<=16'd10815;
      72852:data<=16'd16255;
      72853:data<=16'd13373;
      72854:data<=16'd7370;
      72855:data<=16'd4737;
      72856:data<=16'd4572;
      72857:data<=16'd3997;
      72858:data<=16'd4648;
      72859:data<=16'd3909;
      72860:data<=16'd3269;
      72861:data<=16'd5171;
      72862:data<=16'd5573;
      72863:data<=16'd5809;
      72864:data<=16'd5142;
      72865:data<=16'd3477;
      72866:data<=16'd4868;
      72867:data<=16'd3803;
      72868:data<=16'd1955;
      72869:data<=16'd3336;
      72870:data<=16'd977;
      72871:data<=16'd273;
      72872:data<=16'd3729;
      72873:data<=16'd2702;
      72874:data<=16'd1199;
      72875:data<=16'd1475;
      72876:data<=16'd2158;
      72877:data<=16'd4399;
      72878:data<=16'd3186;
      72879:data<=16'd522;
      72880:data<=-16'd230;
      72881:data<=-16'd901;
      72882:data<=16'd117;
      72883:data<=-16'd59;
      72884:data<=16'd429;
      72885:data<=16'd3222;
      72886:data<=16'd1210;
      72887:data<=16'd156;
      72888:data<=-16'd1877;
      72889:data<=-16'd13277;
      72890:data<=-16'd17887;
      72891:data<=-16'd14534;
      72892:data<=-16'd16487;
      72893:data<=-16'd15797;
      72894:data<=-16'd13311;
      72895:data<=-16'd15174;
      72896:data<=-16'd14292;
      72897:data<=-16'd11728;
      72898:data<=-16'd9444;
      72899:data<=-16'd5125;
      72900:data<=-16'd1994;
      72901:data<=-16'd1368;
      72902:data<=-16'd2259;
      72903:data<=-16'd2705;
      72904:data<=-16'd2170;
      72905:data<=-16'd2779;
      72906:data<=-16'd3015;
      72907:data<=-16'd3104;
      72908:data<=-16'd3726;
      72909:data<=-16'd3184;
      72910:data<=-16'd3284;
      72911:data<=-16'd2981;
      72912:data<=-16'd2302;
      72913:data<=-16'd4408;
      72914:data<=-16'd5291;
      72915:data<=-16'd4073;
      72916:data<=-16'd4614;
      72917:data<=-16'd6088;
      72918:data<=-16'd6769;
      72919:data<=-16'd5210;
      72920:data<=-16'd4764;
      72921:data<=-16'd6634;
      72922:data<=-16'd4361;
      72923:data<=-16'd3002;
      72924:data<=-16'd6808;
      72925:data<=-16'd4875;
      72926:data<=16'd3465;
      72927:data<=16'd9448;
      72928:data<=16'd10542;
      72929:data<=16'd8498;
      72930:data<=16'd7862;
      72931:data<=16'd8446;
      72932:data<=16'd7805;
      72933:data<=16'd7567;
      72934:data<=16'd6839;
      72935:data<=16'd5632;
      72936:data<=16'd5286;
      72937:data<=16'd4408;
      72938:data<=16'd3172;
      72939:data<=16'd1642;
      72940:data<=16'd1027;
      72941:data<=16'd1817;
      72942:data<=-16'd782;
      72943:data<=-16'd6176;
      72944:data<=-16'd8525;
      72945:data<=-16'd7404;
      72946:data<=-16'd7219;
      72947:data<=-16'd8953;
      72948:data<=-16'd7423;
      72949:data<=-16'd5882;
      72950:data<=-16'd9382;
      72951:data<=-16'd9397;
      72952:data<=-16'd6761;
      72953:data<=-16'd8337;
      72954:data<=-16'd8490;
      72955:data<=-16'd7577;
      72956:data<=-16'd7526;
      72957:data<=-16'd6692;
      72958:data<=-16'd8251;
      72959:data<=-16'd7095;
      72960:data<=-16'd4102;
      72961:data<=-16'd5726;
      72962:data<=-16'd4871;
      72963:data<=-16'd9122;
      72964:data<=-16'd23455;
      72965:data<=-16'd27150;
      72966:data<=-16'd22792;
      72967:data<=-16'd23364;
      72968:data<=-16'd22183;
      72969:data<=-16'd21346;
      72970:data<=-16'd21463;
      72971:data<=-16'd18299;
      72972:data<=-16'd18460;
      72973:data<=-16'd18779;
      72974:data<=-16'd16874;
      72975:data<=-16'd18668;
      72976:data<=-16'd17935;
      72977:data<=-16'd15030;
      72978:data<=-16'd16372;
      72979:data<=-16'd16167;
      72980:data<=-16'd14327;
      72981:data<=-16'd13664;
      72982:data<=-16'd12237;
      72983:data<=-16'd12994;
      72984:data<=-16'd13124;
      72985:data<=-16'd10026;
      72986:data<=-16'd10073;
      72987:data<=-16'd9779;
      72988:data<=-16'd5471;
      72989:data<=-16'd4331;
      72990:data<=-16'd4778;
      72991:data<=-16'd2646;
      72992:data<=-16'd2027;
      72993:data<=-16'd2643;
      72994:data<=-16'd2256;
      72995:data<=-16'd2384;
      72996:data<=-16'd2804;
      72997:data<=-16'd2638;
      72998:data<=-16'd2493;
      72999:data<=-16'd3331;
      73000:data<=-16'd1592;
      73001:data<=16'd7178;
      73002:data<=16'd14504;
      73003:data<=16'd13345;
      73004:data<=16'd12490;
      73005:data<=16'd13750;
      73006:data<=16'd11133;
      73007:data<=16'd9409;
      73008:data<=16'd11529;
      73009:data<=16'd11682;
      73010:data<=16'd9624;
      73011:data<=16'd9805;
      73012:data<=16'd10207;
      73013:data<=16'd7444;
      73014:data<=16'd5685;
      73015:data<=16'd5981;
      73016:data<=16'd5137;
      73017:data<=16'd5799;
      73018:data<=16'd6097;
      73019:data<=16'd4200;
      73020:data<=16'd5867;
      73021:data<=16'd6883;
      73022:data<=16'd4710;
      73023:data<=16'd5321;
      73024:data<=16'd4077;
      73025:data<=16'd1855;
      73026:data<=16'd3741;
      73027:data<=16'd2655;
      73028:data<=16'd1154;
      73029:data<=16'd3603;
      73030:data<=16'd3559;
      73031:data<=16'd1457;
      73032:data<=-16'd2584;
      73033:data<=-16'd5755;
      73034:data<=-16'd3057;
      73035:data<=-16'd4520;
      73036:data<=-16'd7342;
      73037:data<=-16'd2957;
      73038:data<=-16'd8034;
      73039:data<=-16'd21570;
      73040:data<=-16'd24119;
      73041:data<=-16'd21159;
      73042:data<=-16'd20168;
      73043:data<=-16'd18950;
      73044:data<=-16'd18724;
      73045:data<=-16'd16933;
      73046:data<=-16'd15646;
      73047:data<=-16'd16806;
      73048:data<=-16'd13943;
      73049:data<=-16'd11743;
      73050:data<=-16'd14607;
      73051:data<=-16'd14049;
      73052:data<=-16'd11415;
      73053:data<=-16'd11688;
      73054:data<=-16'd10749;
      73055:data<=-16'd9708;
      73056:data<=-16'd10774;
      73057:data<=-16'd10201;
      73058:data<=-16'd8536;
      73059:data<=-16'd7928;
      73060:data<=-16'd7115;
      73061:data<=-16'd6463;
      73062:data<=-16'd7453;
      73063:data<=-16'd8805;
      73064:data<=-16'd7570;
      73065:data<=-16'd5917;
      73066:data<=-16'd7639;
      73067:data<=-16'd7694;
      73068:data<=-16'd4549;
      73069:data<=-16'd4331;
      73070:data<=-16'd4460;
      73071:data<=-16'd3300;
      73072:data<=-16'd3855;
      73073:data<=-16'd3078;
      73074:data<=-16'd4077;
      73075:data<=-16'd4529;
      73076:data<=16'd8379;
      73077:data<=16'd22529;
      73078:data<=16'd22557;
      73079:data<=16'd20216;
      73080:data<=16'd20256;
      73081:data<=16'd18706;
      73082:data<=16'd19362;
      73083:data<=16'd19509;
      73084:data<=16'd17373;
      73085:data<=16'd16807;
      73086:data<=16'd16457;
      73087:data<=16'd16020;
      73088:data<=16'd15549;
      73089:data<=16'd13711;
      73090:data<=16'd13009;
      73091:data<=16'd13634;
      73092:data<=16'd13048;
      73093:data<=16'd11723;
      73094:data<=16'd11668;
      73095:data<=16'd11914;
      73096:data<=16'd10046;
      73097:data<=16'd9693;
      73098:data<=16'd11696;
      73099:data<=16'd9961;
      73100:data<=16'd7603;
      73101:data<=16'd8578;
      73102:data<=16'd8082;
      73103:data<=16'd6373;
      73104:data<=16'd5463;
      73105:data<=16'd5228;
      73106:data<=16'd6408;
      73107:data<=16'd5971;
      73108:data<=16'd5557;
      73109:data<=16'd7940;
      73110:data<=16'd7445;
      73111:data<=16'd6288;
      73112:data<=16'd8012;
      73113:data<=16'd2990;
      73114:data<=-16'd8172;
      73115:data<=-16'd12498;
      73116:data<=-16'd10470;
      73117:data<=-16'd10091;
      73118:data<=-16'd9817;
      73119:data<=-16'd7780;
      73120:data<=-16'd9271;
      73121:data<=-16'd14045;
      73122:data<=-16'd16392;
      73123:data<=-16'd16207;
      73124:data<=-16'd14210;
      73125:data<=-16'd11292;
      73126:data<=-16'd10756;
      73127:data<=-16'd10498;
      73128:data<=-16'd8849;
      73129:data<=-16'd8740;
      73130:data<=-16'd8660;
      73131:data<=-16'd7265;
      73132:data<=-16'd6839;
      73133:data<=-16'd7094;
      73134:data<=-16'd6811;
      73135:data<=-16'd6023;
      73136:data<=-16'd5454;
      73137:data<=-16'd4924;
      73138:data<=-16'd3115;
      73139:data<=-16'd1413;
      73140:data<=-16'd855;
      73141:data<=-16'd629;
      73142:data<=-16'd1360;
      73143:data<=-16'd1337;
      73144:data<=16'd276;
      73145:data<=-16'd167;
      73146:data<=-16'd2023;
      73147:data<=-16'd1639;
      73148:data<=-16'd318;
      73149:data<=-16'd529;
      73150:data<=16'd1938;
      73151:data<=16'd11617;
      73152:data<=16'd19898;
      73153:data<=16'd19707;
      73154:data<=16'd19165;
      73155:data<=16'd19858;
      73156:data<=16'd17459;
      73157:data<=16'd16381;
      73158:data<=16'd16568;
      73159:data<=16'd16131;
      73160:data<=16'd16466;
      73161:data<=16'd14481;
      73162:data<=16'd13831;
      73163:data<=16'd16553;
      73164:data<=16'd15341;
      73165:data<=16'd16134;
      73166:data<=16'd22536;
      73167:data<=16'd23787;
      73168:data<=16'd21820;
      73169:data<=16'd21414;
      73170:data<=16'd19760;
      73171:data<=16'd19660;
      73172:data<=16'd19347;
      73173:data<=16'd16430;
      73174:data<=16'd16668;
      73175:data<=16'd18352;
      73176:data<=16'd17518;
      73177:data<=16'd16947;
      73178:data<=16'd17001;
      73179:data<=16'd16122;
      73180:data<=16'd14903;
      73181:data<=16'd14449;
      73182:data<=16'd13259;
      73183:data<=16'd11568;
      73184:data<=16'd12921;
      73185:data<=16'd12756;
      73186:data<=16'd10701;
      73187:data<=16'd13910;
      73188:data<=16'd10836;
      73189:data<=-16'd2567;
      73190:data<=-16'd6519;
      73191:data<=-16'd3306;
      73192:data<=-16'd5266;
      73193:data<=-16'd5805;
      73194:data<=-16'd4992;
      73195:data<=-16'd6307;
      73196:data<=-16'd5676;
      73197:data<=-16'd4554;
      73198:data<=-16'd3797;
      73199:data<=-16'd2992;
      73200:data<=-16'd3432;
      73201:data<=-16'd2745;
      73202:data<=-16'd1847;
      73203:data<=-16'd2343;
      73204:data<=-16'd2476;
      73205:data<=-16'd2866;
      73206:data<=-16'd3033;
      73207:data<=-16'd2846;
      73208:data<=-16'd2702;
      73209:data<=-16'd2288;
      73210:data<=-16'd5970;
      73211:data<=-16'd11088;
      73212:data<=-16'd10363;
      73213:data<=-16'd8856;
      73214:data<=-16'd8731;
      73215:data<=-16'd6470;
      73216:data<=-16'd6067;
      73217:data<=-16'd7045;
      73218:data<=-16'd6266;
      73219:data<=-16'd6313;
      73220:data<=-16'd6581;
      73221:data<=-16'd6390;
      73222:data<=-16'd6197;
      73223:data<=-16'd5403;
      73224:data<=-16'd6573;
      73225:data<=-16'd4983;
      73226:data<=16'd5473;
      73227:data<=16'd14408;
      73228:data<=16'd14944;
      73229:data<=16'd14160;
      73230:data<=16'd13385;
      73231:data<=16'd11682;
      73232:data<=16'd11500;
      73233:data<=16'd11054;
      73234:data<=16'd10825;
      73235:data<=16'd11462;
      73236:data<=16'd9488;
      73237:data<=16'd8943;
      73238:data<=16'd12044;
      73239:data<=16'd11849;
      73240:data<=16'd9873;
      73241:data<=16'd10208;
      73242:data<=16'd9703;
      73243:data<=16'd8637;
      73244:data<=16'd7779;
      73245:data<=16'd6431;
      73246:data<=16'd6088;
      73247:data<=16'd5494;
      73248:data<=16'd5087;
      73249:data<=16'd5908;
      73250:data<=16'd5799;
      73251:data<=16'd6566;
      73252:data<=16'd7209;
      73253:data<=16'd5685;
      73254:data<=16'd7844;
      73255:data<=16'd12521;
      73256:data<=16'd13667;
      73257:data<=16'd12895;
      73258:data<=16'd12129;
      73259:data<=16'd12138;
      73260:data<=16'd11032;
      73261:data<=16'd9101;
      73262:data<=16'd11656;
      73263:data<=16'd8925;
      73264:data<=-16'd4091;
      73265:data<=-16'd8849;
      73266:data<=-16'd5833;
      73267:data<=-16'd7671;
      73268:data<=-16'd7236;
      73269:data<=-16'd5289;
      73270:data<=-16'd7962;
      73271:data<=-16'd8207;
      73272:data<=-16'd6748;
      73273:data<=-16'd7482;
      73274:data<=-16'd7177;
      73275:data<=-16'd6337;
      73276:data<=-16'd5260;
      73277:data<=-16'd4219;
      73278:data<=-16'd4739;
      73279:data<=-16'd4678;
      73280:data<=-16'd4937;
      73281:data<=-16'd5870;
      73282:data<=-16'd4799;
      73283:data<=-16'd4487;
      73284:data<=-16'd5418;
      73285:data<=-16'd5106;
      73286:data<=-16'd5127;
      73287:data<=-16'd4423;
      73288:data<=-16'd2529;
      73289:data<=-16'd2452;
      73290:data<=-16'd3184;
      73291:data<=-16'd3116;
      73292:data<=-16'd2716;
      73293:data<=-16'd3124;
      73294:data<=-16'd4322;
      73295:data<=-16'd3686;
      73296:data<=-16'd3682;
      73297:data<=-16'd4945;
      73298:data<=-16'd3048;
      73299:data<=-16'd5677;
      73300:data<=-16'd11896;
      73301:data<=-16'd4323;
      73302:data<=16'd8041;
      73303:data<=16'd8311;
      73304:data<=16'd6253;
      73305:data<=16'd6449;
      73306:data<=16'd5096;
      73307:data<=16'd5752;
      73308:data<=16'd5683;
      73309:data<=16'd4175;
      73310:data<=16'd4636;
      73311:data<=16'd4029;
      73312:data<=16'd3576;
      73313:data<=16'd4068;
      73314:data<=16'd2895;
      73315:data<=16'd2857;
      73316:data<=16'd2725;
      73317:data<=16'd1292;
      73318:data<=16'd1733;
      73319:data<=16'd1530;
      73320:data<=16'd525;
      73321:data<=16'd258;
      73322:data<=-16'd931;
      73323:data<=-16'd220;
      73324:data<=16'd957;
      73325:data<=-16'd1031;
      73326:data<=-16'd2079;
      73327:data<=-16'd1626;
      73328:data<=-16'd1750;
      73329:data<=-16'd2215;
      73330:data<=-16'd2943;
      73331:data<=-16'd1820;
      73332:data<=-16'd1583;
      73333:data<=-16'd3550;
      73334:data<=-16'd2426;
      73335:data<=-16'd2276;
      73336:data<=-16'd3633;
      73337:data<=-16'd881;
      73338:data<=-16'd5805;
      73339:data<=-16'd20104;
      73340:data<=-16'd24468;
      73341:data<=-16'd21235;
      73342:data<=-16'd22250;
      73343:data<=-16'd20081;
      73344:data<=-16'd13113;
      73345:data<=-16'd10184;
      73346:data<=-16'd10254;
      73347:data<=-16'd10420;
      73348:data<=-16'd10968;
      73349:data<=-16'd9953;
      73350:data<=-16'd9570;
      73351:data<=-16'd11439;
      73352:data<=-16'd11674;
      73353:data<=-16'd10950;
      73354:data<=-16'd10519;
      73355:data<=-16'd9051;
      73356:data<=-16'd8816;
      73357:data<=-16'd9175;
      73358:data<=-16'd8642;
      73359:data<=-16'd8856;
      73360:data<=-16'd8188;
      73361:data<=-16'd7909;
      73362:data<=-16'd9831;
      73363:data<=-16'd10158;
      73364:data<=-16'd9536;
      73365:data<=-16'd9458;
      73366:data<=-16'd8868;
      73367:data<=-16'd8959;
      73368:data<=-16'd8671;
      73369:data<=-16'd8454;
      73370:data<=-16'd9028;
      73371:data<=-16'd8715;
      73372:data<=-16'd9618;
      73373:data<=-16'd9338;
      73374:data<=-16'd7821;
      73375:data<=-16'd9536;
      73376:data<=-16'd4284;
      73377:data<=16'd7521;
      73378:data<=16'd10038;
      73379:data<=16'd8454;
      73380:data<=16'd8851;
      73381:data<=16'd6778;
      73382:data<=16'd6464;
      73383:data<=16'd7040;
      73384:data<=16'd6323;
      73385:data<=16'd6883;
      73386:data<=16'd5862;
      73387:data<=16'd5077;
      73388:data<=16'd3362;
      73389:data<=-16'd2892;
      73390:data<=-16'd5100;
      73391:data<=-16'd3715;
      73392:data<=-16'd4866;
      73393:data<=-16'd4438;
      73394:data<=-16'd3774;
      73395:data<=-16'd4085;
      73396:data<=-16'd3300;
      73397:data<=-16'd3906;
      73398:data<=-16'd3933;
      73399:data<=-16'd3304;
      73400:data<=-16'd4302;
      73401:data<=-16'd4681;
      73402:data<=-16'd5321;
      73403:data<=-16'd4902;
      73404:data<=-16'd3459;
      73405:data<=-16'd4757;
      73406:data<=-16'd4244;
      73407:data<=-16'd2898;
      73408:data<=-16'd4176;
      73409:data<=-16'd3018;
      73410:data<=-16'd3576;
      73411:data<=-16'd4807;
      73412:data<=-16'd325;
      73413:data<=-16'd4579;
      73414:data<=-16'd18777;
      73415:data<=-16'd23443;
      73416:data<=-16'd21184;
      73417:data<=-16'd21309;
      73418:data<=-16'd20345;
      73419:data<=-16'd18968;
      73420:data<=-16'd18685;
      73421:data<=-16'd17605;
      73422:data<=-16'd16827;
      73423:data<=-16'd16258;
      73424:data<=-16'd14634;
      73425:data<=-16'd14099;
      73426:data<=-16'd15449;
      73427:data<=-16'd15429;
      73428:data<=-16'd13923;
      73429:data<=-16'd13517;
      73430:data<=-16'd13361;
      73431:data<=-16'd12609;
      73432:data<=-16'd10884;
      73433:data<=-16'd6975;
      73434:data<=-16'd3368;
      73435:data<=-16'd2370;
      73436:data<=-16'd2291;
      73437:data<=-16'd2123;
      73438:data<=-16'd2804;
      73439:data<=-16'd4344;
      73440:data<=-16'd4687;
      73441:data<=-16'd3830;
      73442:data<=-16'd3624;
      73443:data<=-16'd3219;
      73444:data<=-16'd2403;
      73445:data<=-16'd1444;
      73446:data<=-16'd1101;
      73447:data<=-16'd2776;
      73448:data<=-16'd1905;
      73449:data<=-16'd264;
      73450:data<=-16'd3225;
      73451:data<=16'd1522;
      73452:data<=16'd14269;
      73453:data<=16'd16468;
      73454:data<=16'd13635;
      73455:data<=16'd15746;
      73456:data<=16'd15124;
      73457:data<=16'd13136;
      73458:data<=16'd13605;
      73459:data<=16'd13537;
      73460:data<=16'd13370;
      73461:data<=16'd12566;
      73462:data<=16'd11979;
      73463:data<=16'd11928;
      73464:data<=16'd9592;
      73465:data<=16'd8546;
      73466:data<=16'd9802;
      73467:data<=16'd9485;
      73468:data<=16'd8893;
      73469:data<=16'd8715;
      73470:data<=16'd8787;
      73471:data<=16'd8481;
      73472:data<=16'd6722;
      73473:data<=16'd7259;
      73474:data<=16'd8454;
      73475:data<=16'd7004;
      73476:data<=16'd6587;
      73477:data<=16'd4158;
      73478:data<=-16'd1042;
      73479:data<=-16'd1733;
      73480:data<=-16'd696;
      73481:data<=-16'd1471;
      73482:data<=-16'd1942;
      73483:data<=-16'd2179;
      73484:data<=-16'd632;
      73485:data<=-16'd35;
      73486:data<=-16'd1028;
      73487:data<=16'd1471;
      73488:data<=-16'd2405;
      73489:data<=-16'd15954;
      73490:data<=-16'd21141;
      73491:data<=-16'd18075;
      73492:data<=-16'd18066;
      73493:data<=-16'd17173;
      73494:data<=-16'd15241;
      73495:data<=-16'd15496;
      73496:data<=-16'd14560;
      73497:data<=-16'd13509;
      73498:data<=-16'd13217;
      73499:data<=-16'd11879;
      73500:data<=-16'd11606;
      73501:data<=-16'd12198;
      73502:data<=-16'd11866;
      73503:data<=-16'd11433;
      73504:data<=-16'd10845;
      73505:data<=-16'd10151;
      73506:data<=-16'd9529;
      73507:data<=-16'd8715;
      73508:data<=-16'd8141;
      73509:data<=-16'd7345;
      73510:data<=-16'd6608;
      73511:data<=-16'd6217;
      73512:data<=-16'd5192;
      73513:data<=-16'd4915;
      73514:data<=-16'd5288;
      73515:data<=-16'd4564;
      73516:data<=-16'd4493;
      73517:data<=-16'd4730;
      73518:data<=-16'd4062;
      73519:data<=-16'd3838;
      73520:data<=-16'd2822;
      73521:data<=-16'd1842;
      73522:data<=-16'd705;
      73523:data<=16'd4595;
      73524:data<=16'd6592;
      73525:data<=16'd3145;
      73526:data<=16'd10660;
      73527:data<=16'd25020;
      73528:data<=16'd27129;
      73529:data<=16'd23804;
      73530:data<=16'd24720;
      73531:data<=16'd23461;
      73532:data<=16'd21165;
      73533:data<=16'd21664;
      73534:data<=16'd21318;
      73535:data<=16'd20221;
      73536:data<=16'd19849;
      73537:data<=16'd19133;
      73538:data<=16'd18785;
      73539:data<=16'd19109;
      73540:data<=16'd19387;
      73541:data<=16'd19271;
      73542:data<=16'd18641;
      73543:data<=16'd18134;
      73544:data<=16'd17280;
      73545:data<=16'd15746;
      73546:data<=16'd15048;
      73547:data<=16'd15168;
      73548:data<=16'd14916;
      73549:data<=16'd14157;
      73550:data<=16'd13979;
      73551:data<=16'd15537;
      73552:data<=16'd16613;
      73553:data<=16'd15567;
      73554:data<=16'd14904;
      73555:data<=16'd14891;
      73556:data<=16'd14017;
      73557:data<=16'd12677;
      73558:data<=16'd11708;
      73559:data<=16'd11785;
      73560:data<=16'd10848;
      73561:data<=16'd9597;
      73562:data<=16'd11455;
      73563:data<=16'd8498;
      73564:data<=-16'd2052;
      73565:data<=-16'd6566;
      73566:data<=-16'd6549;
      73567:data<=-16'd11173;
      73568:data<=-16'd12681;
      73569:data<=-16'd10375;
      73570:data<=-16'd11270;
      73571:data<=-16'd11377;
      73572:data<=-16'd10178;
      73573:data<=-16'd10336;
      73574:data<=-16'd9721;
      73575:data<=-16'd9364;
      73576:data<=-16'd8484;
      73577:data<=-16'd6404;
      73578:data<=-16'd6866;
      73579:data<=-16'd7459;
      73580:data<=-16'd5961;
      73581:data<=-16'd5433;
      73582:data<=-16'd5189;
      73583:data<=-16'd4802;
      73584:data<=-16'd4726;
      73585:data<=-16'd3924;
      73586:data<=-16'd4197;
      73587:data<=-16'd5084;
      73588:data<=-16'd4366;
      73589:data<=-16'd2826;
      73590:data<=-16'd1259;
      73591:data<=-16'd1741;
      73592:data<=-16'd3127;
      73593:data<=-16'd1917;
      73594:data<=-16'd1450;
      73595:data<=-16'd1729;
      73596:data<=-16'd425;
      73597:data<=-16'd1163;
      73598:data<=-16'd943;
      73599:data<=16'd429;
      73600:data<=-16'd1475;
      73601:data<=16'd4552;
      73602:data<=16'd18036;
      73603:data<=16'd20648;
      73604:data<=16'd17509;
      73605:data<=16'd18906;
      73606:data<=16'd17919;
      73607:data<=16'd15731;
      73608:data<=16'd16251;
      73609:data<=16'd15458;
      73610:data<=16'd14395;
      73611:data<=16'd15575;
      73612:data<=16'd18286;
      73613:data<=16'd20817;
      73614:data<=16'd21024;
      73615:data<=16'd20395;
      73616:data<=16'd20078;
      73617:data<=16'd18847;
      73618:data<=16'd17499;
      73619:data<=16'd16501;
      73620:data<=16'd15810;
      73621:data<=16'd15377;
      73622:data<=16'd14542;
      73623:data<=16'd14017;
      73624:data<=16'd13556;
      73625:data<=16'd13144;
      73626:data<=16'd13890;
      73627:data<=16'd14125;
      73628:data<=16'd13540;
      73629:data<=16'd13118;
      73630:data<=16'd12128;
      73631:data<=16'd11723;
      73632:data<=16'd11268;
      73633:data<=16'd9662;
      73634:data<=16'd9394;
      73635:data<=16'd8833;
      73636:data<=16'd7404;
      73637:data<=16'd8370;
      73638:data<=16'd5789;
      73639:data<=-16'd3724;
      73640:data<=-16'd9791;
      73641:data<=-16'd9339;
      73642:data<=-16'd9374;
      73643:data<=-16'd10126;
      73644:data<=-16'd9568;
      73645:data<=-16'd9207;
      73646:data<=-16'd8998;
      73647:data<=-16'd9021;
      73648:data<=-16'd9185;
      73649:data<=-16'd8493;
      73650:data<=-16'd8275;
      73651:data<=-16'd7303;
      73652:data<=-16'd4655;
      73653:data<=-16'd4485;
      73654:data<=-16'd5413;
      73655:data<=-16'd5894;
      73656:data<=-16'd9539;
      73657:data<=-16'd12020;
      73658:data<=-16'd11323;
      73659:data<=-16'd12214;
      73660:data<=-16'd11530;
      73661:data<=-16'd9841;
      73662:data<=-16'd11321;
      73663:data<=-16'd10983;
      73664:data<=-16'd8880;
      73665:data<=-16'd8804;
      73666:data<=-16'd8479;
      73667:data<=-16'd7837;
      73668:data<=-16'd7800;
      73669:data<=-16'd7926;
      73670:data<=-16'd7353;
      73671:data<=-16'd6244;
      73672:data<=-16'd7309;
      73673:data<=-16'd7050;
      73674:data<=-16'd5711;
      73675:data<=-16'd8278;
      73676:data<=-16'd2608;
      73677:data<=16'd12064;
      73678:data<=16'd15215;
      73679:data<=16'd11333;
      73680:data<=16'd12889;
      73681:data<=16'd12968;
      73682:data<=16'd11159;
      73683:data<=16'd10654;
      73684:data<=16'd9465;
      73685:data<=16'd9414;
      73686:data<=16'd9555;
      73687:data<=16'd9075;
      73688:data<=16'd9579;
      73689:data<=16'd9256;
      73690:data<=16'd8812;
      73691:data<=16'd9219;
      73692:data<=16'd8774;
      73693:data<=16'd7761;
      73694:data<=16'd6637;
      73695:data<=16'd5727;
      73696:data<=16'd5151;
      73697:data<=16'd5187;
      73698:data<=16'd5679;
      73699:data<=16'd4711;
      73700:data<=16'd5796;
      73701:data<=16'd10467;
      73702:data<=16'd12020;
      73703:data<=16'd11435;
      73704:data<=16'd11593;
      73705:data<=16'd9969;
      73706:data<=16'd9139;
      73707:data<=16'd8648;
      73708:data<=16'd7116;
      73709:data<=16'd8117;
      73710:data<=16'd7618;
      73711:data<=16'd5629;
      73712:data<=16'd7203;
      73713:data<=16'd3612;
      73714:data<=-16'd7470;
      73715:data<=-16'd13655;
      73716:data<=-16'd13392;
      73717:data<=-16'd13176;
      73718:data<=-16'd13405;
      73719:data<=-16'd12625;
      73720:data<=-16'd11856;
      73721:data<=-16'd12034;
      73722:data<=-16'd11952;
      73723:data<=-16'd11195;
      73724:data<=-16'd10757;
      73725:data<=-16'd11230;
      73726:data<=-16'd12733;
      73727:data<=-16'd13571;
      73728:data<=-16'd13220;
      73729:data<=-16'd13086;
      73730:data<=-16'd12760;
      73731:data<=-16'd12407;
      73732:data<=-16'd12119;
      73733:data<=-16'd11235;
      73734:data<=-16'd10951;
      73735:data<=-16'd10871;
      73736:data<=-16'd10798;
      73737:data<=-16'd11547;
      73738:data<=-16'd11700;
      73739:data<=-16'd12199;
      73740:data<=-16'd12992;
      73741:data<=-16'd12192;
      73742:data<=-16'd12222;
      73743:data<=-16'd11923;
      73744:data<=-16'd10040;
      73745:data<=-16'd11875;
      73746:data<=-16'd16307;
      73747:data<=-16'd17688;
      73748:data<=-16'd15711;
      73749:data<=-16'd14557;
      73750:data<=-16'd16172;
      73751:data<=-16'd11449;
      73752:data<=16'd523;
      73753:data<=16'd4379;
      73754:data<=16'd1454;
      73755:data<=16'd2353;
      73756:data<=16'd2978;
      73757:data<=16'd1717;
      73758:data<=16'd1249;
      73759:data<=16'd846;
      73760:data<=16'd1682;
      73761:data<=16'd2035;
      73762:data<=16'd1472;
      73763:data<=16'd1971;
      73764:data<=16'd435;
      73765:data<=-16'd1650;
      73766:data<=-16'd819;
      73767:data<=-16'd397;
      73768:data<=-16'd846;
      73769:data<=-16'd311;
      73770:data<=-16'd177;
      73771:data<=-16'd1186;
      73772:data<=-16'd1792;
      73773:data<=-16'd679;
      73774:data<=-16'd79;
      73775:data<=-16'd544;
      73776:data<=-16'd220;
      73777:data<=-16'd1260;
      73778:data<=-16'd2262;
      73779:data<=-16'd1069;
      73780:data<=-16'd1528;
      73781:data<=-16'd2146;
      73782:data<=-16'd1666;
      73783:data<=-16'd2338;
      73784:data<=-16'd1158;
      73785:data<=-16'd846;
      73786:data<=-16'd2546;
      73787:data<=-16'd732;
      73788:data<=-16'd3855;
      73789:data<=-16'd14146;
      73790:data<=-16'd17156;
      73791:data<=-16'd14683;
      73792:data<=-16'd14786;
      73793:data<=-16'd14254;
      73794:data<=-16'd13229;
      73795:data<=-16'd12924;
      73796:data<=-16'd12502;
      73797:data<=-16'd12401;
      73798:data<=-16'd11594;
      73799:data<=-16'd11362;
      73800:data<=-16'd11596;
      73801:data<=-16'd10907;
      73802:data<=-16'd11984;
      73803:data<=-16'd12457;
      73804:data<=-16'd10557;
      73805:data<=-16'd10672;
      73806:data<=-16'd10269;
      73807:data<=-16'd8091;
      73808:data<=-16'd8583;
      73809:data<=-16'd9009;
      73810:data<=-16'd7887;
      73811:data<=-16'd8119;
      73812:data<=-16'd8146;
      73813:data<=-16'd7982;
      73814:data<=-16'd9028;
      73815:data<=-16'd9468;
      73816:data<=-16'd9150;
      73817:data<=-16'd9270;
      73818:data<=-16'd9544;
      73819:data<=-16'd8563;
      73820:data<=-16'd6828;
      73821:data<=-16'd7714;
      73822:data<=-16'd8992;
      73823:data<=-16'd6429;
      73824:data<=-16'd5871;
      73825:data<=-16'd8364;
      73826:data<=-16'd2108;
      73827:data<=16'd10157;
      73828:data<=16'd13063;
      73829:data<=16'd10301;
      73830:data<=16'd11118;
      73831:data<=16'd10266;
      73832:data<=16'd8543;
      73833:data<=16'd10254;
      73834:data<=16'd8455;
      73835:data<=16'd3956;
      73836:data<=16'd3483;
      73837:data<=16'd3582;
      73838:data<=16'd3046;
      73839:data<=16'd3309;
      73840:data<=16'd1642;
      73841:data<=-16'd35;
      73842:data<=16'd288;
      73843:data<=16'd453;
      73844:data<=16'd540;
      73845:data<=16'd745;
      73846:data<=16'd920;
      73847:data<=16'd1296;
      73848:data<=16'd1081;
      73849:data<=16'd1249;
      73850:data<=16'd2008;
      73851:data<=16'd1327;
      73852:data<=-16'd364;
      73853:data<=-16'd822;
      73854:data<=16'd200;
      73855:data<=16'd447;
      73856:data<=-16'd206;
      73857:data<=16'd212;
      73858:data<=16'd858;
      73859:data<=16'd1604;
      73860:data<=16'd2112;
      73861:data<=16'd1074;
      73862:data<=16'd1698;
      73863:data<=-16'd167;
      73864:data<=-16'd11139;
      73865:data<=-16'd19600;
      73866:data<=-16'd18744;
      73867:data<=-16'd18230;
      73868:data<=-16'd18183;
      73869:data<=-16'd15948;
      73870:data<=-16'd15611;
      73871:data<=-16'd15393;
      73872:data<=-16'd13744;
      73873:data<=-16'd13073;
      73874:data<=-16'd12848;
      73875:data<=-16'd12163;
      73876:data<=-16'd11985;
      73877:data<=-16'd13535;
      73878:data<=-16'd13076;
      73879:data<=-16'd7838;
      73880:data<=-16'd4993;
      73881:data<=-16'd5322;
      73882:data<=-16'd3068;
      73883:data<=-16'd2185;
      73884:data<=-16'd2960;
      73885:data<=-16'd1556;
      73886:data<=-16'd1724;
      73887:data<=-16'd2634;
      73888:data<=-16'd2338;
      73889:data<=-16'd3353;
      73890:data<=-16'd3398;
      73891:data<=-16'd3133;
      73892:data<=-16'd4355;
      73893:data<=-16'd3692;
      73894:data<=-16'd2722;
      73895:data<=-16'd2132;
      73896:data<=-16'd785;
      73897:data<=-16'd1557;
      73898:data<=-16'd1080;
      73899:data<=16'd143;
      73900:data<=-16'd2291;
      73901:data<=16'd2719;
      73902:data<=16'd15403;
      73903:data<=16'd18255;
      73904:data<=16'd14966;
      73905:data<=16'd16189;
      73906:data<=16'd15998;
      73907:data<=16'd14060;
      73908:data<=16'd14769;
      73909:data<=16'd14656;
      73910:data<=16'd13634;
      73911:data<=16'd14084;
      73912:data<=16'd13990;
      73913:data<=16'd13089;
      73914:data<=16'd12954;
      73915:data<=16'd13060;
      73916:data<=16'd12897;
      73917:data<=16'd12596;
      73918:data<=16'd11916;
      73919:data<=16'd11097;
      73920:data<=16'd10698;
      73921:data<=16'd11001;
      73922:data<=16'd11247;
      73923:data<=16'd8994;
      73924:data<=16'd4643;
      73925:data<=16'd2643;
      73926:data<=16'd3768;
      73927:data<=16'd5098;
      73928:data<=16'd5918;
      73929:data<=16'd6247;
      73930:data<=16'd6228;
      73931:data<=16'd6560;
      73932:data<=16'd6472;
      73933:data<=16'd6269;
      73934:data<=16'd6927;
      73935:data<=16'd6357;
      73936:data<=16'd5118;
      73937:data<=16'd6228;
      73938:data<=16'd4052;
      73939:data<=-16'd5662;
      73940:data<=-16'd12279;
      73941:data<=-16'd11062;
      73942:data<=-16'd10684;
      73943:data<=-16'd11035;
      73944:data<=-16'd9360;
      73945:data<=-16'd9407;
      73946:data<=-16'd8839;
      73947:data<=-16'd7174;
      73948:data<=-16'd7702;
      73949:data<=-16'd6949;
      73950:data<=-16'd6182;
      73951:data<=-16'd7321;
      73952:data<=-16'd5268;
      73953:data<=-16'd2811;
      73954:data<=-16'd3151;
      73955:data<=-16'd2869;
      73956:data<=-16'd2617;
      73957:data<=-16'd2006;
      73958:data<=-16'd719;
      73959:data<=-16'd980;
      73960:data<=-16'd878;
      73961:data<=-16'd694;
      73962:data<=-16'd1246;
      73963:data<=-16'd954;
      73964:data<=-16'd654;
      73965:data<=16'd1061;
      73966:data<=16'd2003;
      73967:data<=16'd563;
      73968:data<=16'd4285;
      73969:data<=16'd9086;
      73970:data<=16'd8229;
      73971:data<=16'd8100;
      73972:data<=16'd7791;
      73973:data<=16'd7066;
      73974:data<=16'd8467;
      73975:data<=16'd6626;
      73976:data<=16'd11033;
      73977:data<=16'd25062;
      73978:data<=16'd29144;
      73979:data<=16'd25799;
      73980:data<=16'd26699;
      73981:data<=16'd25485;
      73982:data<=16'd23604;
      73983:data<=16'd23933;
      73984:data<=16'd22365;
      73985:data<=16'd21476;
      73986:data<=16'd21535;
      73987:data<=16'd20879;
      73988:data<=16'd20378;
      73989:data<=16'd19144;
      73990:data<=16'd19176;
      73991:data<=16'd19752;
      73992:data<=16'd18184;
      73993:data<=16'd17365;
      73994:data<=16'd16777;
      73995:data<=16'd15156;
      73996:data<=16'd14707;
      73997:data<=16'd14273;
      73998:data<=16'd13753;
      73999:data<=16'd13690;
      74000:data<=16'd12948;
      74001:data<=16'd12888;
      74002:data<=16'd13417;
      74003:data<=16'd13599;
      74004:data<=16'd13647;
      74005:data<=16'd12857;
      74006:data<=16'd12087;
      74007:data<=16'd11230;
      74008:data<=16'd10419;
      74009:data<=16'd11186;
      74010:data<=16'd10426;
      74011:data<=16'd8669;
      74012:data<=16'd8349;
      74013:data<=16'd2188;
      74014:data<=-16'd9617;
      74015:data<=-16'd15658;
      74016:data<=-16'd15423;
      74017:data<=-16'd14968;
      74018:data<=-16'd14609;
      74019:data<=-16'd13916;
      74020:data<=-16'd13609;
      74021:data<=-16'd13232;
      74022:data<=-16'd12460;
      74023:data<=-16'd11982;
      74024:data<=-16'd11690;
      74025:data<=-16'd11315;
      74026:data<=-16'd11600;
      74027:data<=-16'd11119;
      74028:data<=-16'd8813;
      74029:data<=-16'd7559;
      74030:data<=-16'd8023;
      74031:data<=-16'd7830;
      74032:data<=-16'd7031;
      74033:data<=-16'd6808;
      74034:data<=-16'd6824;
      74035:data<=-16'd6504;
      74036:data<=-16'd6187;
      74037:data<=-16'd6047;
      74038:data<=-16'd6079;
      74039:data<=-16'd5683;
      74040:data<=-16'd3771;
      74041:data<=-16'd2817;
      74042:data<=-16'd3668;
      74043:data<=-16'd2335;
      74044:data<=-16'd916;
      74045:data<=-16'd1851;
      74046:data<=-16'd1788;
      74047:data<=-16'd1876;
      74048:data<=-16'd1654;
      74049:data<=-16'd743;
      74050:data<=-16'd2755;
      74051:data<=16'd1535;
      74052:data<=16'd13861;
      74053:data<=16'd17593;
      74054:data<=16'd15547;
      74055:data<=16'd16409;
      74056:data<=16'd14345;
      74057:data<=16'd14803;
      74058:data<=16'd20237;
      74059:data<=16'd20315;
      74060:data<=16'd18061;
      74061:data<=16'd17943;
      74062:data<=16'd16750;
      74063:data<=16'd16028;
      74064:data<=16'd15879;
      74065:data<=16'd15969;
      74066:data<=16'd16677;
      74067:data<=16'd15044;
      74068:data<=16'd13159;
      74069:data<=16'd13054;
      74070:data<=16'd12026;
      74071:data<=16'd11063;
      74072:data<=16'd10475;
      74073:data<=16'd9476;
      74074:data<=16'd9712;
      74075:data<=16'd9512;
      74076:data<=16'd7952;
      74077:data<=16'd7823;
      74078:data<=16'd9066;
      74079:data<=16'd9219;
      74080:data<=16'd7764;
      74081:data<=16'd7103;
      74082:data<=16'd7371;
      74083:data<=16'd6326;
      74084:data<=16'd6023;
      74085:data<=16'd6138;
      74086:data<=16'd4155;
      74087:data<=16'd4134;
      74088:data<=16'd3468;
      74089:data<=-16'd4487;
      74090:data<=-16'd11160;
      74091:data<=-16'd10731;
      74092:data<=-16'd10681;
      74093:data<=-16'd11160;
      74094:data<=-16'd9624;
      74095:data<=-16'd10137;
      74096:data<=-16'd11356;
      74097:data<=-16'd10366;
      74098:data<=-16'd10307;
      74099:data<=-16'd10883;
      74100:data<=-16'd9835;
      74101:data<=-16'd10621;
      74102:data<=-16'd13841;
      74103:data<=-16'd14595;
      74104:data<=-16'd13432;
      74105:data<=-16'd13396;
      74106:data<=-16'd12592;
      74107:data<=-16'd11358;
      74108:data<=-16'd11966;
      74109:data<=-16'd12236;
      74110:data<=-16'd11700;
      74111:data<=-16'd11825;
      74112:data<=-16'd11147;
      74113:data<=-16'd10369;
      74114:data<=-16'd10780;
      74115:data<=-16'd10751;
      74116:data<=-16'd10637;
      74117:data<=-16'd10628;
      74118:data<=-16'd9911;
      74119:data<=-16'd9899;
      74120:data<=-16'd9906;
      74121:data<=-16'd9643;
      74122:data<=-16'd10402;
      74123:data<=-16'd9292;
      74124:data<=-16'd8182;
      74125:data<=-16'd9777;
      74126:data<=-16'd4616;
      74127:data<=16'd6040;
      74128:data<=16'd7696;
      74129:data<=16'd4570;
      74130:data<=16'd5347;
      74131:data<=16'd4913;
      74132:data<=16'd3955;
      74133:data<=16'd4400;
      74134:data<=16'd3058;
      74135:data<=16'd3198;
      74136:data<=16'd4264;
      74137:data<=16'd3051;
      74138:data<=16'd3230;
      74139:data<=16'd2843;
      74140:data<=16'd411;
      74141:data<=16'd441;
      74142:data<=16'd277;
      74143:data<=-16'd948;
      74144:data<=-16'd834;
      74145:data<=-16'd1947;
      74146:data<=-16'd675;
      74147:data<=16'd4485;
      74148:data<=16'd5927;
      74149:data<=16'd4532;
      74150:data<=16'd4232;
      74151:data<=16'd3451;
      74152:data<=16'd2504;
      74153:data<=16'd1365;
      74154:data<=16'd710;
      74155:data<=16'd1410;
      74156:data<=16'd1045;
      74157:data<=16'd641;
      74158:data<=16'd895;
      74159:data<=16'd161;
      74160:data<=16'd132;
      74161:data<=-16'd123;
      74162:data<=-16'd755;
      74163:data<=-16'd1303;
      74164:data<=-16'd8169;
      74165:data<=-16'd17520;
      74166:data<=-16'd18880;
      74167:data<=-16'd17534;
      74168:data<=-16'd18375;
      74169:data<=-16'd17450;
      74170:data<=-16'd16393;
      74171:data<=-16'd16651;
      74172:data<=-16'd16407;
      74173:data<=-16'd16028;
      74174:data<=-16'd15534;
      74175:data<=-16'd14986;
      74176:data<=-16'd14301;
      74177:data<=-16'd13866;
      74178:data<=-16'd14853;
      74179:data<=-16'd14889;
      74180:data<=-16'd13388;
      74181:data<=-16'd13159;
      74182:data<=-16'd12851;
      74183:data<=-16'd11618;
      74184:data<=-16'd11570;
      74185:data<=-16'd11862;
      74186:data<=-16'd11224;
      74187:data<=-16'd10809;
      74188:data<=-16'd11016;
      74189:data<=-16'd10328;
      74190:data<=-16'd10325;
      74191:data<=-16'd14495;
      74192:data<=-16'd18252;
      74193:data<=-16'd17276;
      74194:data<=-16'd16319;
      74195:data<=-16'd15917;
      74196:data<=-16'd14662;
      74197:data<=-16'd14916;
      74198:data<=-16'd13729;
      74199:data<=-16'd12492;
      74200:data<=-16'd14295;
      74201:data<=-16'd9274;
      74202:data<=16'd1691;
      74203:data<=16'd4443;
      74204:data<=16'd2103;
      74205:data<=16'd2673;
      74206:data<=16'd2881;
      74207:data<=16'd2463;
      74208:data<=16'd2781;
      74209:data<=16'd2441;
      74210:data<=16'd2713;
      74211:data<=16'd3360;
      74212:data<=16'd2999;
      74213:data<=16'd2943;
      74214:data<=16'd2825;
      74215:data<=16'd1378;
      74216:data<=16'd0;
      74217:data<=-16'd253;
      74218:data<=-16'd264;
      74219:data<=-16'd346;
      74220:data<=-16'd141;
      74221:data<=-16'd288;
      74222:data<=-16'd569;
      74223:data<=16'd152;
      74224:data<=16'd484;
      74225:data<=-16'd540;
      74226:data<=-16'd775;
      74227:data<=-16'd688;
      74228:data<=-16'd2079;
      74229:data<=-16'd2469;
      74230:data<=-16'd1222;
      74231:data<=-16'd1060;
      74232:data<=-16'd1030;
      74233:data<=-16'd704;
      74234:data<=-16'd1201;
      74235:data<=16'd397;
      74236:data<=16'd3914;
      74237:data<=16'd5814;
      74238:data<=16'd5238;
      74239:data<=-16'd1019;
      74240:data<=-16'd10551;
      74241:data<=-16'd13400;
      74242:data<=-16'd11606;
      74243:data<=-16'd11665;
      74244:data<=-16'd11091;
      74245:data<=-16'd10141;
      74246:data<=-16'd10163;
      74247:data<=-16'd9383;
      74248:data<=-16'd9257;
      74249:data<=-16'd9441;
      74250:data<=-16'd8448;
      74251:data<=-16'd7808;
      74252:data<=-16'd7756;
      74253:data<=-16'd8258;
      74254:data<=-16'd8589;
      74255:data<=-16'd7814;
      74256:data<=-16'd7253;
      74257:data<=-16'd6364;
      74258:data<=-16'd5638;
      74259:data<=-16'd6401;
      74260:data<=-16'd6067;
      74261:data<=-16'd5018;
      74262:data<=-16'd4996;
      74263:data<=-16'd4858;
      74264:data<=-16'd4916;
      74265:data<=-16'd4775;
      74266:data<=-16'd4993;
      74267:data<=-16'd5893;
      74268:data<=-16'd4877;
      74269:data<=-16'd4581;
      74270:data<=-16'd5500;
      74271:data<=-16'd4287;
      74272:data<=-16'd4043;
      74273:data<=-16'd3451;
      74274:data<=-16'd2355;
      74275:data<=-16'd4670;
      74276:data<=-16'd27;
      74277:data<=16'd11312;
      74278:data<=16'd13315;
      74279:data<=16'd10396;
      74280:data<=16'd8934;
      74281:data<=16'd4742;
      74282:data<=16'd3371;
      74283:data<=16'd4992;
      74284:data<=16'd4329;
      74285:data<=16'd4695;
      74286:data<=16'd5357;
      74287:data<=16'd4751;
      74288:data<=16'd5106;
      74289:data<=16'd4946;
      74290:data<=16'd3953;
      74291:data<=16'd2689;
      74292:data<=16'd1538;
      74293:data<=16'd1965;
      74294:data<=16'd2087;
      74295:data<=16'd1827;
      74296:data<=16'd2629;
      74297:data<=16'd2607;
      74298:data<=16'd2513;
      74299:data<=16'd2836;
      74300:data<=16'd1992;
      74301:data<=16'd2167;
      74302:data<=16'd3294;
      74303:data<=16'd2287;
      74304:data<=16'd834;
      74305:data<=16'd1384;
      74306:data<=16'd2129;
      74307:data<=16'd1685;
      74308:data<=16'd1660;
      74309:data<=16'd2440;
      74310:data<=16'd2120;
      74311:data<=16'd795;
      74312:data<=16'd1530;
      74313:data<=16'd2981;
      74314:data<=-16'd2470;
      74315:data<=-16'd11928;
      74316:data<=-16'd13947;
      74317:data<=-16'd12098;
      74318:data<=-16'd12440;
      74319:data<=-16'd10836;
      74320:data<=-16'd9784;
      74321:data<=-16'd10258;
      74322:data<=-16'd8909;
      74323:data<=-16'd9561;
      74324:data<=-16'd8360;
      74325:data<=-16'd2138;
      74326:data<=16'd77;
      74327:data<=-16'd211;
      74328:data<=16'd1751;
      74329:data<=16'd2083;
      74330:data<=16'd1764;
      74331:data<=16'd2237;
      74332:data<=16'd2807;
      74333:data<=16'd3714;
      74334:data<=16'd3295;
      74335:data<=16'd3066;
      74336:data<=16'd3879;
      74337:data<=16'd4214;
      74338:data<=16'd4692;
      74339:data<=16'd4247;
      74340:data<=16'd4413;
      74341:data<=16'd6008;
      74342:data<=16'd5800;
      74343:data<=16'd6091;
      74344:data<=16'd6396;
      74345:data<=16'd5147;
      74346:data<=16'd6466;
      74347:data<=16'd7235;
      74348:data<=16'd6833;
      74349:data<=16'd7598;
      74350:data<=16'd5348;
      74351:data<=16'd8373;
      74352:data<=16'd19748;
      74353:data<=16'd24095;
      74354:data<=16'd22747;
      74355:data<=16'd23306;
      74356:data<=16'd22177;
      74357:data<=16'd21162;
      74358:data<=16'd20663;
      74359:data<=16'd19650;
      74360:data<=16'd20360;
      74361:data<=16'd19602;
      74362:data<=16'd18319;
      74363:data<=16'd18733;
      74364:data<=16'd17596;
      74365:data<=16'd17212;
      74366:data<=16'd18057;
      74367:data<=16'd17449;
      74368:data<=16'd17094;
      74369:data<=16'd14463;
      74370:data<=16'd9291;
      74371:data<=16'd7655;
      74372:data<=16'd8711;
      74373:data<=16'd8754;
      74374:data<=16'd8011;
      74375:data<=16'd7474;
      74376:data<=16'd7627;
      74377:data<=16'd7180;
      74378:data<=16'd6739;
      74379:data<=16'd8200;
      74380:data<=16'd8675;
      74381:data<=16'd7341;
      74382:data<=16'd7420;
      74383:data<=16'd7227;
      74384:data<=16'd6150;
      74385:data<=16'd6989;
      74386:data<=16'd6614;
      74387:data<=16'd5583;
      74388:data<=16'd7062;
      74389:data<=16'd1841;
      74390:data<=-16'd8834;
      74391:data<=-16'd9879;
      74392:data<=-16'd6742;
      74393:data<=-16'd8232;
      74394:data<=-16'd7680;
      74395:data<=-16'd6504;
      74396:data<=-16'd7436;
      74397:data<=-16'd6592;
      74398:data<=-16'd6217;
      74399:data<=-16'd6721;
      74400:data<=-16'd6317;
      74401:data<=-16'd6156;
      74402:data<=-16'd5268;
      74403:data<=-16'd4311;
      74404:data<=-16'd3436;
      74405:data<=-16'd2059;
      74406:data<=-16'd2447;
      74407:data<=-16'd2682;
      74408:data<=-16'd1591;
      74409:data<=-16'd1160;
      74410:data<=-16'd581;
      74411:data<=-16'd1069;
      74412:data<=-16'd2026;
      74413:data<=-16'd341;
      74414:data<=16'd2922;
      74415:data<=16'd6319;
      74416:data<=16'd7371;
      74417:data<=16'd6818;
      74418:data<=16'd7876;
      74419:data<=16'd6881;
      74420:data<=16'd5824;
      74421:data<=16'd7890;
      74422:data<=16'd7163;
      74423:data<=16'd6537;
      74424:data<=16'd7045;
      74425:data<=16'd3987;
      74426:data<=16'd7427;
      74427:data<=16'd18072;
      74428:data<=16'd22545;
      74429:data<=16'd22431;
      74430:data<=16'd22134;
      74431:data<=16'd20500;
      74432:data<=16'd19617;
      74433:data<=16'd19164;
      74434:data<=16'd18589;
      74435:data<=16'd18060;
      74436:data<=16'd16678;
      74437:data<=16'd16149;
      74438:data<=16'd16061;
      74439:data<=16'd15009;
      74440:data<=16'd14442;
      74441:data<=16'd14562;
      74442:data<=16'd14718;
      74443:data<=16'd14129;
      74444:data<=16'd12938;
      74445:data<=16'd12342;
      74446:data<=16'd11345;
      74447:data<=16'd10390;
      74448:data<=16'd10549;
      74449:data<=16'd9483;
      74450:data<=16'd7753;
      74451:data<=16'd7941;
      74452:data<=16'd7934;
      74453:data<=16'd7056;
      74454:data<=16'd8069;
      74455:data<=16'd8360;
      74456:data<=16'd6667;
      74457:data<=16'd7617;
      74458:data<=16'd6347;
      74459:data<=-16'd61;
      74460:data<=-16'd1641;
      74461:data<=-16'd949;
      74462:data<=-16'd2299;
      74463:data<=16'd130;
      74464:data<=-16'd3739;
      74465:data<=-16'd15420;
      74466:data<=-16'd17211;
      74467:data<=-16'd13882;
      74468:data<=-16'd14728;
      74469:data<=-16'd14223;
      74470:data<=-16'd13944;
      74471:data<=-16'd14463;
      74472:data<=-16'd13987;
      74473:data<=-16'd14422;
      74474:data<=-16'd13450;
      74475:data<=-16'd12769;
      74476:data<=-16'd13644;
      74477:data<=-16'd12549;
      74478:data<=-16'd11345;
      74479:data<=-16'd10047;
      74480:data<=-16'd8886;
      74481:data<=-16'd9615;
      74482:data<=-16'd8404;
      74483:data<=-16'd7203;
      74484:data<=-16'd7906;
      74485:data<=-16'd6784;
      74486:data<=-16'd6334;
      74487:data<=-16'd6482;
      74488:data<=-16'd5768;
      74489:data<=-16'd6877;
      74490:data<=-16'd7036;
      74491:data<=-16'd5858;
      74492:data<=-16'd5106;
      74493:data<=-16'd3726;
      74494:data<=-16'd4106;
      74495:data<=-16'd4073;
      74496:data<=-16'd2628;
      74497:data<=-16'd3924;
      74498:data<=-16'd3698;
      74499:data<=-16'd2701;
      74500:data<=-16'd5042;
      74501:data<=-16'd1723;
      74502:data<=16'd8487;
      74503:data<=16'd16164;
      74504:data<=16'd19884;
      74505:data<=16'd20727;
      74506:data<=16'd19170;
      74507:data<=16'd17867;
      74508:data<=16'd17625;
      74509:data<=16'd17067;
      74510:data<=16'd16045;
      74511:data<=16'd15890;
      74512:data<=16'd15338;
      74513:data<=16'd13996;
      74514:data<=16'd13722;
      74515:data<=16'd12464;
      74516:data<=16'd10672;
      74517:data<=16'd10975;
      74518:data<=16'd10586;
      74519:data<=16'd9215;
      74520:data<=16'd8721;
      74521:data<=16'd8031;
      74522:data<=16'd7301;
      74523:data<=16'd6907;
      74524:data<=16'd6570;
      74525:data<=16'd5463;
      74526:data<=16'd4355;
      74527:data<=16'd5007;
      74528:data<=16'd3891;
      74529:data<=16'd1657;
      74530:data<=16'd2027;
      74531:data<=16'd1034;
      74532:data<=-16'd33;
      74533:data<=16'd634;
      74534:data<=-16'd519;
      74535:data<=16'd105;
      74536:data<=16'd412;
      74537:data<=-16'd1389;
      74538:data<=16'd693;
      74539:data<=-16'd3325;
      74540:data<=-16'd15211;
      74541:data<=-16'd18953;
      74542:data<=-16'd18262;
      74543:data<=-16'd19324;
      74544:data<=-16'd18302;
      74545:data<=-16'd18008;
      74546:data<=-16'd17465;
      74547:data<=-16'd18022;
      74548:data<=-16'd22563;
      74549:data<=-16'd23608;
      74550:data<=-16'd22266;
      74551:data<=-16'd22480;
      74552:data<=-16'd20797;
      74553:data<=-16'd20340;
      74554:data<=-16'd21617;
      74555:data<=-16'd21229;
      74556:data<=-16'd20336;
      74557:data<=-16'd18679;
      74558:data<=-16'd18045;
      74559:data<=-16'd18419;
      74560:data<=-16'd16954;
      74561:data<=-16'd16460;
      74562:data<=-16'd16245;
      74563:data<=-16'd15036;
      74564:data<=-16'd15300;
      74565:data<=-16'd14659;
      74566:data<=-16'd14687;
      74567:data<=-16'd16622;
      74568:data<=-16'd15494;
      74569:data<=-16'd14451;
      74570:data<=-16'd14798;
      74571:data<=-16'd12966;
      74572:data<=-16'd12828;
      74573:data<=-16'd12774;
      74574:data<=-16'd10754;
      74575:data<=-16'd12082;
      74576:data<=-16'd9559;
      74577:data<=16'd1356;
      74578:data<=16'd6297;
      74579:data<=16'd3036;
      74580:data<=16'd2834;
      74581:data<=16'd4052;
      74582:data<=16'd2726;
      74583:data<=16'd2743;
      74584:data<=16'd3548;
      74585:data<=16'd3134;
      74586:data<=16'd3331;
      74587:data<=16'd3474;
      74588:data<=16'd2826;
      74589:data<=16'd2560;
      74590:data<=16'd1780;
      74591:data<=16'd613;
      74592:data<=16'd1712;
      74593:data<=16'd4969;
      74594:data<=16'd6222;
      74595:data<=16'd4919;
      74596:data<=16'd5065;
      74597:data<=16'd5153;
      74598:data<=16'd3629;
      74599:data<=16'd4055;
      74600:data<=16'd4191;
      74601:data<=16'd2927;
      74602:data<=16'd3685;
      74603:data<=16'd3336;
      74604:data<=16'd1856;
      74605:data<=16'd1764;
      74606:data<=16'd446;
      74607:data<=16'd226;
      74608:data<=16'd872;
      74609:data<=-16'd182;
      74610:data<=16'd1028;
      74611:data<=16'd779;
      74612:data<=-16'd989;
      74613:data<=16'd1718;
      74614:data<=-16'd2657;
      74615:data<=-16'd14499;
      74616:data<=-16'd17206;
      74617:data<=-16'd16301;
      74618:data<=-16'd18600;
      74619:data<=-16'd17599;
      74620:data<=-16'd16334;
      74621:data<=-16'd16205;
      74622:data<=-16'd14698;
      74623:data<=-16'd14607;
      74624:data<=-16'd14287;
      74625:data<=-16'd13230;
      74626:data<=-16'd13324;
      74627:data<=-16'd12484;
      74628:data<=-16'd12073;
      74629:data<=-16'd12789;
      74630:data<=-16'd12625;
      74631:data<=-16'd12511;
      74632:data<=-16'd11632;
      74633:data<=-16'd10339;
      74634:data<=-16'd10082;
      74635:data<=-16'd9048;
      74636:data<=-16'd9327;
      74637:data<=-16'd12443;
      74638:data<=-16'd14637;
      74639:data<=-16'd14692;
      74640:data<=-16'd13418;
      74641:data<=-16'd13247;
      74642:data<=-16'd14800;
      74643:data<=-16'd14123;
      74644:data<=-16'd12863;
      74645:data<=-16'd12649;
      74646:data<=-16'd10862;
      74647:data<=-16'd10642;
      74648:data<=-16'd10762;
      74649:data<=-16'd8639;
      74650:data<=-16'd9815;
      74651:data<=-16'd7674;
      74652:data<=16'd3480;
      74653:data<=16'd8865;
      74654:data<=16'd6084;
      74655:data<=16'd6216;
      74656:data<=16'd7060;
      74657:data<=16'd6256;
      74658:data<=16'd6683;
      74659:data<=16'd6886;
      74660:data<=16'd6696;
      74661:data<=16'd6658;
      74662:data<=16'd6445;
      74663:data<=16'd6740;
      74664:data<=16'd6542;
      74665:data<=16'd5786;
      74666:data<=16'd4899;
      74667:data<=16'd3347;
      74668:data<=16'd2843;
      74669:data<=16'd3219;
      74670:data<=16'd2772;
      74671:data<=16'd2528;
      74672:data<=16'd2590;
      74673:data<=16'd2951;
      74674:data<=16'd3698;
      74675:data<=16'd3189;
      74676:data<=16'd2488;
      74677:data<=16'd2840;
      74678:data<=16'd2930;
      74679:data<=16'd2332;
      74680:data<=16'd1030;
      74681:data<=16'd2171;
      74682:data<=16'd6884;
      74683:data<=16'd7965;
      74684:data<=16'd6240;
      74685:data<=16'd7667;
      74686:data<=16'd7037;
      74687:data<=16'd5838;
      74688:data<=16'd8746;
      74689:data<=16'd4011;
      74690:data<=-16'd7733;
      74691:data<=-16'd10903;
      74692:data<=-16'd9542;
      74693:data<=-16'd10880;
      74694:data<=-16'd10307;
      74695:data<=-16'd9492;
      74696:data<=-16'd9709;
      74697:data<=-16'd8467;
      74698:data<=-16'd8141;
      74699:data<=-16'd8116;
      74700:data<=-16'd7529;
      74701:data<=-16'd8211;
      74702:data<=-16'd7526;
      74703:data<=-16'd5674;
      74704:data<=-16'd5868;
      74705:data<=-16'd6620;
      74706:data<=-16'd6595;
      74707:data<=-16'd6032;
      74708:data<=-16'd5483;
      74709:data<=-16'd5592;
      74710:data<=-16'd5162;
      74711:data<=-16'd4261;
      74712:data<=-16'd3488;
      74713:data<=-16'd2834;
      74714:data<=-16'd3286;
      74715:data<=-16'd3203;
      74716:data<=-16'd2083;
      74717:data<=-16'd2074;
      74718:data<=-16'd1827;
      74719:data<=-16'd1407;
      74720:data<=-16'd1466;
      74721:data<=-16'd247;
      74722:data<=-16'd9;
      74723:data<=-16'd167;
      74724:data<=16'd1269;
      74725:data<=-16'd657;
      74726:data<=-16'd1833;
      74727:data<=16'd5065;
      74728:data<=16'd10721;
      74729:data<=16'd10319;
      74730:data<=16'd11365;
      74731:data<=16'd12701;
      74732:data<=16'd11561;
      74733:data<=16'd11394;
      74734:data<=16'd11512;
      74735:data<=16'd11019;
      74736:data<=16'd11241;
      74737:data<=16'd10840;
      74738:data<=16'd10417;
      74739:data<=16'd10787;
      74740:data<=16'd10190;
      74741:data<=16'd10006;
      74742:data<=16'd11126;
      74743:data<=16'd11388;
      74744:data<=16'd10927;
      74745:data<=16'd10592;
      74746:data<=16'd10528;
      74747:data<=16'd10464;
      74748:data<=16'd9761;
      74749:data<=16'd9547;
      74750:data<=16'd9539;
      74751:data<=16'd9113;
      74752:data<=16'd9289;
      74753:data<=16'd8705;
      74754:data<=16'd8837;
      74755:data<=16'd10924;
      74756:data<=16'd10496;
      74757:data<=16'd9216;
      74758:data<=16'd9436;
      74759:data<=16'd8671;
      74760:data<=16'd8883;
      74761:data<=16'd8152;
      74762:data<=16'd6798;
      74763:data<=16'd9711;
      74764:data<=16'd5859;
      74765:data<=-16'd6416;
      74766:data<=-16'd9201;
      74767:data<=-16'd5280;
      74768:data<=-16'd5846;
      74769:data<=-16'd6467;
      74770:data<=-16'd3650;
      74771:data<=16'd1090;
      74772:data<=16'd3303;
      74773:data<=16'd1748;
      74774:data<=16'd2118;
      74775:data<=16'd2845;
      74776:data<=16'd1961;
      74777:data<=16'd2713;
      74778:data<=16'd2919;
      74779:data<=16'd3137;
      74780:data<=16'd4726;
      74781:data<=16'd4355;
      74782:data<=16'd3980;
      74783:data<=16'd4708;
      74784:data<=16'd4390;
      74785:data<=16'd4041;
      74786:data<=16'd3914;
      74787:data<=16'd4434;
      74788:data<=16'd4846;
      74789:data<=16'd3902;
      74790:data<=16'd4084;
      74791:data<=16'd4532;
      74792:data<=16'd4643;
      74793:data<=16'd6209;
      74794:data<=16'd6229;
      74795:data<=16'd5604;
      74796:data<=16'd6243;
      74797:data<=16'd4915;
      74798:data<=16'd4880;
      74799:data<=16'd6504;
      74800:data<=16'd4040;
      74801:data<=16'd5310;
      74802:data<=16'd15778;
      74803:data<=16'd21854;
      74804:data<=16'd19647;
      74805:data<=16'd20204;
      74806:data<=16'd21920;
      74807:data<=16'd19717;
      74808:data<=16'd19077;
      74809:data<=16'd19074;
      74810:data<=16'd17203;
      74811:data<=16'd17244;
      74812:data<=16'd16587;
      74813:data<=16'd15582;
      74814:data<=16'd16489;
      74815:data<=16'd12609;
      74816:data<=16'd7315;
      74817:data<=16'd7871;
      74818:data<=16'd9195;
      74819:data<=16'd9391;
      74820:data<=16'd9045;
      74821:data<=16'd7462;
      74822:data<=16'd7400;
      74823:data<=16'd7256;
      74824:data<=16'd6035;
      74825:data<=16'd5752;
      74826:data<=16'd5589;
      74827:data<=16'd5645;
      74828:data<=16'd4798;
      74829:data<=16'd4511;
      74830:data<=16'd6786;
      74831:data<=16'd6755;
      74832:data<=16'd6109;
      74833:data<=16'd6596;
      74834:data<=16'd4725;
      74835:data<=16'd5121;
      74836:data<=16'd5247;
      74837:data<=16'd2986;
      74838:data<=16'd5651;
      74839:data<=16'd1876;
      74840:data<=-16'd11000;
      74841:data<=-16'd13396;
      74842:data<=-16'd9459;
      74843:data<=-16'd9773;
      74844:data<=-16'd9347;
      74845:data<=-16'd9130;
      74846:data<=-16'd9253;
      74847:data<=-16'd8382;
      74848:data<=-16'd8851;
      74849:data<=-16'd8449;
      74850:data<=-16'd8005;
      74851:data<=-16'd8416;
      74852:data<=-16'd7805;
      74853:data<=-16'd7911;
      74854:data<=-16'd6874;
      74855:data<=-16'd4872;
      74856:data<=-16'd5134;
      74857:data<=-16'd5009;
      74858:data<=-16'd4742;
      74859:data<=-16'd3715;
      74860:data<=16'd619;
      74861:data<=16'd2952;
      74862:data<=16'd2511;
      74863:data<=16'd2537;
      74864:data<=16'd1666;
      74865:data<=16'd1515;
      74866:data<=16'd2105;
      74867:data<=16'd2096;
      74868:data<=16'd3253;
      74869:data<=16'd3357;
      74870:data<=16'd2441;
      74871:data<=16'd2801;
      74872:data<=16'd2093;
      74873:data<=16'd2106;
      74874:data<=16'd3200;
      74875:data<=16'd1157;
      74876:data<=16'd2428;
      74877:data<=16'd11497;
      74878:data<=16'd17493;
      74879:data<=16'd16880;
      74880:data<=16'd17224;
      74881:data<=16'd17567;
      74882:data<=16'd15590;
      74883:data<=16'd15121;
      74884:data<=16'd14938;
      74885:data<=16'd13593;
      74886:data<=16'd13214;
      74887:data<=16'd12320;
      74888:data<=16'd11668;
      74889:data<=16'd12219;
      74890:data<=16'd10975;
      74891:data<=16'd9882;
      74892:data<=16'd10298;
      74893:data<=16'd10346;
      74894:data<=16'd11130;
      74895:data<=16'd10748;
      74896:data<=16'd8587;
      74897:data<=16'd7926;
      74898:data<=16'd7514;
      74899:data<=16'd6953;
      74900:data<=16'd6552;
      74901:data<=16'd5092;
      74902:data<=16'd5162;
      74903:data<=16'd5797;
      74904:data<=16'd3733;
      74905:data<=16'd817;
      74906:data<=-16'd1061;
      74907:data<=-16'd926;
      74908:data<=-16'd729;
      74909:data<=-16'd1855;
      74910:data<=-16'd1328;
      74911:data<=-16'd2228;
      74912:data<=-16'd3654;
      74913:data<=-16'd629;
      74914:data<=-16'd4425;
      74915:data<=-16'd16307;
      74916:data<=-16'd19329;
      74917:data<=-16'd16387;
      74918:data<=-16'd17068;
      74919:data<=-16'd17205;
      74920:data<=-16'd16616;
      74921:data<=-16'd16548;
      74922:data<=-16'd15570;
      74923:data<=-16'd15405;
      74924:data<=-16'd15023;
      74925:data<=-16'd14096;
      74926:data<=-16'd14468;
      74927:data<=-16'd14242;
      74928:data<=-16'd12983;
      74929:data<=-16'd12495;
      74930:data<=-16'd13336;
      74931:data<=-16'd14695;
      74932:data<=-16'd14146;
      74933:data<=-16'd12665;
      74934:data<=-16'd12624;
      74935:data<=-16'd12443;
      74936:data<=-16'd11996;
      74937:data<=-16'd11732;
      74938:data<=-16'd10895;
      74939:data<=-16'd11192;
      74940:data<=-16'd11547;
      74941:data<=-16'd10351;
      74942:data<=-16'd10716;
      74943:data<=-16'd12187;
      74944:data<=-16'd12622;
      74945:data<=-16'd12589;
      74946:data<=-16'd11245;
      74947:data<=-16'd10422;
      74948:data<=-16'd9964;
      74949:data<=-16'd6031;
      74950:data<=-16'd3764;
      74951:data<=-16'd3193;
      74952:data<=16'd5043;
      74953:data<=16'd13133;
      74954:data<=16'd11361;
      74955:data<=16'd8675;
      74956:data<=16'd8980;
      74957:data<=16'd8285;
      74958:data<=16'd7611;
      74959:data<=16'd6934;
      74960:data<=16'd6173;
      74961:data<=16'd6091;
      74962:data<=16'd5598;
      74963:data<=16'd5297;
      74964:data<=16'd5150;
      74965:data<=16'd4861;
      74966:data<=16'd4877;
      74967:data<=16'd3519;
      74968:data<=16'd1971;
      74969:data<=16'd1999;
      74970:data<=16'd1744;
      74971:data<=16'd1425;
      74972:data<=16'd986;
      74973:data<=-16'd102;
      74974:data<=16'd83;
      74975:data<=16'd417;
      74976:data<=16'd23;
      74977:data<=16'd288;
      74978:data<=16'd156;
      74979:data<=-16'd170;
      74980:data<=-16'd757;
      74981:data<=-16'd2373;
      74982:data<=-16'd2623;
      74983:data<=-16'd2584;
      74984:data<=-16'd3174;
      74985:data<=-16'd2038;
      74986:data<=-16'd2779;
      74987:data<=-16'd4208;
      74988:data<=-16'd1055;
      74989:data<=-16'd3424;
      74990:data<=-16'd14781;
      74991:data<=-16'd18821;
      74992:data<=-16'd15549;
      74993:data<=-16'd18924;
      74994:data<=-16'd24562;
      74995:data<=-16'd24294;
      74996:data<=-16'd23037;
      74997:data<=-16'd22983;
      74998:data<=-16'd21638;
      74999:data<=-16'd20404;
      75000:data<=-16'd19784;
      75001:data<=-16'd18647;
      75002:data<=-16'd17843;
      75003:data<=-16'd17371;
      75004:data<=-16'd16481;
      75005:data<=-16'd16413;
      75006:data<=-16'd17614;
      75007:data<=-16'd17691;
      75008:data<=-16'd15984;
      75009:data<=-16'd14859;
      75010:data<=-16'd14692;
      75011:data<=-16'd14411;
      75012:data<=-16'd13670;
      75013:data<=-16'd11963;
      75014:data<=-16'd11056;
      75015:data<=-16'd11808;
      75016:data<=-16'd11405;
      75017:data<=-16'd10806;
      75018:data<=-16'd11864;
      75019:data<=-16'd12217;
      75020:data<=-16'd11709;
      75021:data<=-16'd11203;
      75022:data<=-16'd10313;
      75023:data<=-16'd9458;
      75024:data<=-16'd8451;
      75025:data<=-16'd8981;
      75026:data<=-16'd8605;
      75027:data<=-16'd384;
      75028:data<=16'd8481;
      75029:data<=16'd8116;
      75030:data<=16'd5444;
      75031:data<=16'd5509;
      75032:data<=16'd5304;
      75033:data<=16'd5042;
      75034:data<=16'd4969;
      75035:data<=16'd5228;
      75036:data<=16'd5118;
      75037:data<=16'd4541;
      75038:data<=16'd7821;
      75039:data<=16'd11744;
      75040:data<=16'd10783;
      75041:data<=16'd9950;
      75042:data<=16'd10019;
      75043:data<=16'd8158;
      75044:data<=16'd7783;
      75045:data<=16'd8005;
      75046:data<=16'd7047;
      75047:data<=16'd7191;
      75048:data<=16'd7154;
      75049:data<=16'd6473;
      75050:data<=16'd6402;
      75051:data<=16'd6037;
      75052:data<=16'd5829;
      75053:data<=16'd6285;
      75054:data<=16'd6381;
      75055:data<=16'd4827;
      75056:data<=16'd3025;
      75057:data<=16'd4065;
      75058:data<=16'd4429;
      75059:data<=16'd2658;
      75060:data<=16'd3535;
      75061:data<=16'd3356;
      75062:data<=16'd1786;
      75063:data<=16'd4314;
      75064:data<=16'd1048;
      75065:data<=-16'd10246;
      75066:data<=-16'd13802;
      75067:data<=-16'd11430;
      75068:data<=-16'd13118;
      75069:data<=-16'd13885;
      75070:data<=-16'd12005;
      75071:data<=-16'd11714;
      75072:data<=-16'd11251;
      75073:data<=-16'd9682;
      75074:data<=-16'd9191;
      75075:data<=-16'd9344;
      75076:data<=-16'd8971;
      75077:data<=-16'd8319;
      75078:data<=-16'd7400;
      75079:data<=-16'd6872;
      75080:data<=-16'd7454;
      75081:data<=-16'd7950;
      75082:data<=-16'd9380;
      75083:data<=-16'd12789;
      75084:data<=-16'd13864;
      75085:data<=-16'd12182;
      75086:data<=-16'd12034;
      75087:data<=-16'd11720;
      75088:data<=-16'd9858;
      75089:data<=-16'd9647;
      75090:data<=-16'd10110;
      75091:data<=-16'd9206;
      75092:data<=-16'd9091;
      75093:data<=-16'd10061;
      75094:data<=-16'd9964;
      75095:data<=-16'd9254;
      75096:data<=-16'd8834;
      75097:data<=-16'd8138;
      75098:data<=-16'd7318;
      75099:data<=-16'd6502;
      75100:data<=-16'd6613;
      75101:data<=-16'd6234;
      75102:data<=16'd884;
      75103:data<=16'd10611;
      75104:data<=16'd11643;
      75105:data<=16'd8451;
      75106:data<=16'd8343;
      75107:data<=16'd7759;
      75108:data<=16'd7100;
      75109:data<=16'd7891;
      75110:data<=16'd7746;
      75111:data<=16'd7332;
      75112:data<=16'd6942;
      75113:data<=16'd6748;
      75114:data<=16'd7122;
      75115:data<=16'd6578;
      75116:data<=16'd6166;
      75117:data<=16'd5780;
      75118:data<=16'd5233;
      75119:data<=16'd6473;
      75120:data<=16'd6461;
      75121:data<=16'd5075;
      75122:data<=16'd5412;
      75123:data<=16'd5021;
      75124:data<=16'd5175;
      75125:data<=16'd6028;
      75126:data<=16'd4440;
      75127:data<=16'd6355;
      75128:data<=16'd11477;
      75129:data<=16'd12019;
      75130:data<=16'd11476;
      75131:data<=16'd12800;
      75132:data<=16'd12985;
      75133:data<=16'd12420;
      75134:data<=16'd12087;
      75135:data<=16'd12311;
      75136:data<=16'd11262;
      75137:data<=16'd9976;
      75138:data<=16'd12081;
      75139:data<=16'd8986;
      75140:data<=-16'd2388;
      75141:data<=-16'd7166;
      75142:data<=-16'd3745;
      75143:data<=-16'd2290;
      75144:data<=-16'd1962;
      75145:data<=-16'd1078;
      75146:data<=-16'd1130;
      75147:data<=-16'd810;
      75148:data<=-16'd476;
      75149:data<=-16'd714;
      75150:data<=-16'd631;
      75151:data<=-16'd470;
      75152:data<=-16'd284;
      75153:data<=-16'd14;
      75154:data<=16'd109;
      75155:data<=16'd883;
      75156:data<=16'd2311;
      75157:data<=16'd2796;
      75158:data<=16'd2666;
      75159:data<=16'd3269;
      75160:data<=16'd3301;
      75161:data<=16'd2681;
      75162:data<=16'd3295;
      75163:data<=16'd3977;
      75164:data<=16'd3465;
      75165:data<=16'd2629;
      75166:data<=16'd2181;
      75167:data<=16'd3256;
      75168:data<=16'd4928;
      75169:data<=16'd5069;
      75170:data<=16'd4952;
      75171:data<=16'd4366;
      75172:data<=16'd917;
      75173:data<=-16'd2003;
      75174:data<=-16'd1080;
      75175:data<=-16'd1293;
      75176:data<=-16'd2317;
      75177:data<=16'd4708;
      75178:data<=16'd14202;
      75179:data<=16'd14246;
      75180:data<=16'd12258;
      75181:data<=16'd14891;
      75182:data<=16'd14889;
      75183:data<=16'd13203;
      75184:data<=16'd13731;
      75185:data<=16'd12989;
      75186:data<=16'd11887;
      75187:data<=16'd12105;
      75188:data<=16'd11394;
      75189:data<=16'd10411;
      75190:data<=16'd10126;
      75191:data<=16'd9671;
      75192:data<=16'd9523;
      75193:data<=16'd10608;
      75194:data<=16'd11571;
      75195:data<=16'd10725;
      75196:data<=16'd9931;
      75197:data<=16'd9817;
      75198:data<=16'd8851;
      75199:data<=16'd8704;
      75200:data<=16'd9086;
      75201:data<=16'd8419;
      75202:data<=16'd8272;
      75203:data<=16'd7697;
      75204:data<=16'd7106;
      75205:data<=16'd8624;
      75206:data<=16'd9342;
      75207:data<=16'd9027;
      75208:data<=16'd9080;
      75209:data<=16'd8251;
      75210:data<=16'd8326;
      75211:data<=16'd7777;
      75212:data<=16'd6119;
      75213:data<=16'd7981;
      75214:data<=16'd5059;
      75215:data<=-16'd6343;
      75216:data<=-16'd8716;
      75217:data<=-16'd1234;
      75218:data<=16'd578;
      75219:data<=-16'd409;
      75220:data<=16'd1415;
      75221:data<=16'd1331;
      75222:data<=16'd221;
      75223:data<=16'd396;
      75224:data<=16'd472;
      75225:data<=16'd722;
      75226:data<=16'd523;
      75227:data<=-16'd11;
      75228:data<=16'd519;
      75229:data<=16'd889;
      75230:data<=16'd1290;
      75231:data<=16'd2364;
      75232:data<=16'd2516;
      75233:data<=16'd2675;
      75234:data<=16'd3333;
      75235:data<=16'd2801;
      75236:data<=16'd2127;
      75237:data<=16'd1903;
      75238:data<=16'd1249;
      75239:data<=16'd1055;
      75240:data<=16'd1306;
      75241:data<=16'd1155;
      75242:data<=16'd1318;
      75243:data<=16'd2591;
      75244:data<=16'd3600;
      75245:data<=16'd2796;
      75246:data<=16'd2288;
      75247:data<=16'd2652;
      75248:data<=16'd2165;
      75249:data<=16'd2886;
      75250:data<=16'd2886;
      75251:data<=16'd848;
      75252:data<=16'd6229;
      75253:data<=16'd16305;
      75254:data<=16'd17253;
      75255:data<=16'd14454;
      75256:data<=16'd16471;
      75257:data<=16'd16944;
      75258:data<=16'd14771;
      75259:data<=16'd14624;
      75260:data<=16'd13894;
      75261:data<=16'd10111;
      75262:data<=16'd6869;
      75263:data<=16'd6250;
      75264:data<=16'd5717;
      75265:data<=16'd4915;
      75266:data<=16'd4868;
      75267:data<=16'd4302;
      75268:data<=16'd4813;
      75269:data<=16'd6561;
      75270:data<=16'd5823;
      75271:data<=16'd4642;
      75272:data<=16'd5065;
      75273:data<=16'd4528;
      75274:data<=16'd4014;
      75275:data<=16'd4211;
      75276:data<=16'd3982;
      75277:data<=16'd4056;
      75278:data<=16'd3629;
      75279:data<=16'd2995;
      75280:data<=16'd3284;
      75281:data<=16'd3635;
      75282:data<=16'd4831;
      75283:data<=16'd5318;
      75284:data<=16'd3770;
      75285:data<=16'd3673;
      75286:data<=16'd3266;
      75287:data<=16'd2196;
      75288:data<=16'd4194;
      75289:data<=16'd717;
      75290:data<=-16'd10234;
      75291:data<=-16'd13949;
      75292:data<=-16'd11449;
      75293:data<=-16'd11893;
      75294:data<=-16'd10998;
      75295:data<=-16'd9221;
      75296:data<=-16'd9835;
      75297:data<=-16'd9047;
      75298:data<=-16'd8715;
      75299:data<=-16'd9785;
      75300:data<=-16'd8890;
      75301:data<=-16'd8601;
      75302:data<=-16'd8436;
      75303:data<=-16'd7077;
      75304:data<=-16'd7938;
      75305:data<=-16'd6425;
      75306:data<=-16'd370;
      75307:data<=16'd2003;
      75308:data<=16'd819;
      75309:data<=16'd936;
      75310:data<=16'd1152;
      75311:data<=16'd860;
      75312:data<=16'd341;
      75313:data<=-16'd164;
      75314:data<=-16'd230;
      75315:data<=-16'd553;
      75316:data<=-16'd450;
      75317:data<=-16'd560;
      75318:data<=-16'd1419;
      75319:data<=-16'd1237;
      75320:data<=-16'd1456;
      75321:data<=-16'd1676;
      75322:data<=-16'd723;
      75323:data<=-16'd1821;
      75324:data<=-16'd1989;
      75325:data<=-16'd682;
      75326:data<=-16'd2792;
      75327:data<=16'd895;
      75328:data<=16'd11932;
      75329:data<=16'd14254;
      75330:data<=16'd10404;
      75331:data<=16'd10091;
      75332:data<=16'd8490;
      75333:data<=16'd6734;
      75334:data<=16'd7674;
      75335:data<=16'd6896;
      75336:data<=16'd5964;
      75337:data<=16'd6158;
      75338:data<=16'd5016;
      75339:data<=16'd4488;
      75340:data<=16'd4748;
      75341:data<=16'd3641;
      75342:data<=16'd2441;
      75343:data<=16'd1783;
      75344:data<=16'd464;
      75345:data<=-16'd378;
      75346:data<=16'd179;
      75347:data<=-16'd622;
      75348:data<=-16'd1900;
      75349:data<=-16'd640;
      75350:data<=-16'd2015;
      75351:data<=-16'd7080;
      75352:data<=-16'd8307;
      75353:data<=-16'd7068;
      75354:data<=-16'd7078;
      75355:data<=-16'd7154;
      75356:data<=-16'd8737;
      75357:data<=-16'd9611;
      75358:data<=-16'd8420;
      75359:data<=-16'd8907;
      75360:data<=-16'd8815;
      75361:data<=-16'd8410;
      75362:data<=-16'd9379;
      75363:data<=-16'd7289;
      75364:data<=-16'd9091;
      75365:data<=-16'd19297;
      75366:data<=-16'd23916;
      75367:data<=-16'd21517;
      75368:data<=-16'd22043;
      75369:data<=-16'd22950;
      75370:data<=-16'd22001;
      75371:data<=-16'd21723;
      75372:data<=-16'd21061;
      75373:data<=-16'd19925;
      75374:data<=-16'd19021;
      75375:data<=-16'd18477;
      75376:data<=-16'd18246;
      75377:data<=-16'd17262;
      75378:data<=-16'd16233;
      75379:data<=-16'd15603;
      75380:data<=-16'd14980;
      75381:data<=-16'd15650;
      75382:data<=-16'd16280;
      75383:data<=-16'd15346;
      75384:data<=-16'd14930;
      75385:data<=-16'd14678;
      75386:data<=-16'd13614;
      75387:data<=-16'd12988;
      75388:data<=-16'd12128;
      75389:data<=-16'd11659;
      75390:data<=-16'd12392;
      75391:data<=-16'd11236;
      75392:data<=-16'd9715;
      75393:data<=-16'd11062;
      75394:data<=-16'd10948;
      75395:data<=-16'd7843;
      75396:data<=-16'd5492;
      75397:data<=-16'd4551;
      75398:data<=-16'd4557;
      75399:data<=-16'd3821;
      75400:data<=-16'd3413;
      75401:data<=-16'd5486;
      75402:data<=-16'd792;
      75403:data<=16'd10980;
      75404:data<=16'd13653;
      75405:data<=16'd9621;
      75406:data<=16'd9450;
      75407:data<=16'd8463;
      75408:data<=16'd7019;
      75409:data<=16'd7749;
      75410:data<=16'd6884;
      75411:data<=16'd6728;
      75412:data<=16'd7362;
      75413:data<=16'd6244;
      75414:data<=16'd6234;
      75415:data<=16'd6284;
      75416:data<=16'd5341;
      75417:data<=16'd5260;
      75418:data<=16'd4194;
      75419:data<=16'd2441;
      75420:data<=16'd1862;
      75421:data<=16'd1839;
      75422:data<=16'd1955;
      75423:data<=16'd1730;
      75424:data<=16'd1626;
      75425:data<=16'd1343;
      75426:data<=16'd647;
      75427:data<=16'd1175;
      75428:data<=16'd1296;
      75429:data<=16'd854;
      75430:data<=16'd1245;
      75431:data<=16'd124;
      75432:data<=-16'd684;
      75433:data<=-16'd593;
      75434:data<=-16'd1811;
      75435:data<=-16'd801;
      75436:data<=-16'd459;
      75437:data<=-16'd2009;
      75438:data<=16'd890;
      75439:data<=-16'd2306;
      75440:data<=-16'd16032;
      75441:data<=-16'd21494;
      75442:data<=-16'd18116;
      75443:data<=-16'd18747;
      75444:data<=-16'd20400;
      75445:data<=-16'd19268;
      75446:data<=-16'd17908;
      75447:data<=-16'd17176;
      75448:data<=-16'd16653;
      75449:data<=-16'd15597;
      75450:data<=-16'd14818;
      75451:data<=-16'd14340;
      75452:data<=-16'd13386;
      75453:data<=-16'd13194;
      75454:data<=-16'd12716;
      75455:data<=-16'd11338;
      75456:data<=-16'd11658;
      75457:data<=-16'd12825;
      75458:data<=-16'd12466;
      75459:data<=-16'd11207;
      75460:data<=-16'd9920;
      75461:data<=-16'd8995;
      75462:data<=-16'd8668;
      75463:data<=-16'd8326;
      75464:data<=-16'd7797;
      75465:data<=-16'd7467;
      75466:data<=-16'd7098;
      75467:data<=-16'd6995;
      75468:data<=-16'd7357;
      75469:data<=-16'd7380;
      75470:data<=-16'd7656;
      75471:data<=-16'd7418;
      75472:data<=-16'd5979;
      75473:data<=-16'd6206;
      75474:data<=-16'd5761;
      75475:data<=-16'd4255;
      75476:data<=-16'd6413;
      75477:data<=-16'd2361;
      75478:data<=16'd10023;
      75479:data<=16'd12774;
      75480:data<=16'd9568;
      75481:data<=16'd10995;
      75482:data<=16'd8895;
      75483:data<=16'd7175;
      75484:data<=16'd11257;
      75485:data<=16'd12185;
      75486:data<=16'd11165;
      75487:data<=16'd11521;
      75488:data<=16'd10804;
      75489:data<=16'd10983;
      75490:data<=16'd11042;
      75491:data<=16'd10100;
      75492:data<=16'd10046;
      75493:data<=16'd9527;
      75494:data<=16'd8595;
      75495:data<=16'd7257;
      75496:data<=16'd6129;
      75497:data<=16'd6778;
      75498:data<=16'd6402;
      75499:data<=16'd5483;
      75500:data<=16'd5849;
      75501:data<=16'd5426;
      75502:data<=16'd5520;
      75503:data<=16'd5868;
      75504:data<=16'd5353;
      75505:data<=16'd5894;
      75506:data<=16'd4996;
      75507:data<=16'd3153;
      75508:data<=16'd3392;
      75509:data<=16'd3024;
      75510:data<=16'd2604;
      75511:data<=16'd2641;
      75512:data<=16'd2432;
      75513:data<=16'd4529;
      75514:data<=16'd1991;
      75515:data<=-16'd8434;
      75516:data<=-16'd13597;
      75517:data<=-16'd11292;
      75518:data<=-16'd10448;
      75519:data<=-16'd10807;
      75520:data<=-16'd10272;
      75521:data<=-16'd9585;
      75522:data<=-16'd8658;
      75523:data<=-16'd7818;
      75524:data<=-16'd7031;
      75525:data<=-16'd6858;
      75526:data<=-16'd6825;
      75527:data<=-16'd5498;
      75528:data<=-16'd5940;
      75529:data<=-16'd9297;
      75530:data<=-16'd10308;
      75531:data<=-16'd8032;
      75532:data<=-16'd6282;
      75533:data<=-16'd5579;
      75534:data<=-16'd5115;
      75535:data<=-16'd4585;
      75536:data<=-16'd3659;
      75537:data<=-16'd3178;
      75538:data<=-16'd3024;
      75539:data<=-16'd2670;
      75540:data<=-16'd2322;
      75541:data<=-16'd1504;
      75542:data<=-16'd1339;
      75543:data<=-16'd1419;
      75544:data<=16'd274;
      75545:data<=16'd905;
      75546:data<=16'd661;
      75547:data<=16'd1868;
      75548:data<=16'd1245;
      75549:data<=16'd1234;
      75550:data<=16'd2590;
      75551:data<=16'd349;
      75552:data<=16'd4225;
      75553:data<=16'd15932;
      75554:data<=16'd18218;
      75555:data<=16'd14577;
      75556:data<=16'd16322;
      75557:data<=16'd16995;
      75558:data<=16'd15932;
      75559:data<=16'd16774;
      75560:data<=16'd16274;
      75561:data<=16'd15488;
      75562:data<=16'd15324;
      75563:data<=16'd14316;
      75564:data<=16'd13925;
      75565:data<=16'd13723;
      75566:data<=16'd12950;
      75567:data<=16'd12181;
      75568:data<=16'd11444;
      75569:data<=16'd12069;
      75570:data<=16'd13459;
      75571:data<=16'd12998;
      75572:data<=16'd11753;
      75573:data<=16'd12511;
      75574:data<=16'd14292;
      75575:data<=16'd14208;
      75576:data<=16'd13123;
      75577:data<=16'd12739;
      75578:data<=16'd12076;
      75579:data<=16'd11694;
      75580:data<=16'd11812;
      75581:data<=16'd11603;
      75582:data<=16'd12666;
      75583:data<=16'd13403;
      75584:data<=16'd12088;
      75585:data<=16'd12007;
      75586:data<=16'd11615;
      75587:data<=16'd9638;
      75588:data<=16'd10395;
      75589:data<=16'd8431;
      75590:data<=-16'd1107;
      75591:data<=-16'd7141;
      75592:data<=-16'd6032;
      75593:data<=-16'd5761;
      75594:data<=-16'd5201;
      75595:data<=-16'd3106;
      75596:data<=-16'd3432;
      75597:data<=-16'd3639;
      75598:data<=-16'd2544;
      75599:data<=-16'd2664;
      75600:data<=-16'd2594;
      75601:data<=-16'd2796;
      75602:data<=-16'd3548;
      75603:data<=-16'd2732;
      75604:data<=-16'd2466;
      75605:data<=-16'd3131;
      75606:data<=-16'd2315;
      75607:data<=-16'd1060;
      75608:data<=-16'd165;
      75609:data<=16'd177;
      75610:data<=16'd124;
      75611:data<=16'd487;
      75612:data<=16'd403;
      75613:data<=16'd741;
      75614:data<=16'd1130;
      75615:data<=16'd343;
      75616:data<=16'd1118;
      75617:data<=16'd506;
      75618:data<=-16'd3168;
      75619:data<=-16'd3034;
      75620:data<=-16'd1406;
      75621:data<=-16'd1767;
      75622:data<=-16'd731;
      75623:data<=-16'd1010;
      75624:data<=-16'd1251;
      75625:data<=-16'd306;
      75626:data<=-16'd2928;
      75627:data<=16'd870;
      75628:data<=16'd12754;
      75629:data<=16'd15173;
      75630:data<=16'd11611;
      75631:data<=16'd13073;
      75632:data<=16'd13985;
      75633:data<=16'd13571;
      75634:data<=16'd13697;
      75635:data<=16'd12273;
      75636:data<=16'd11594;
      75637:data<=16'd11497;
      75638:data<=16'd10821;
      75639:data<=16'd10840;
      75640:data<=16'd10339;
      75641:data<=16'd9737;
      75642:data<=16'd9429;
      75643:data<=16'd8345;
      75644:data<=16'd8493;
      75645:data<=16'd9611;
      75646:data<=16'd9421;
      75647:data<=16'd8672;
      75648:data<=16'd7921;
      75649:data<=16'd7051;
      75650:data<=16'd6426;
      75651:data<=16'd6404;
      75652:data<=16'd6464;
      75653:data<=16'd5416;
      75654:data<=16'd4579;
      75655:data<=16'd4751;
      75656:data<=16'd5080;
      75657:data<=16'd6355;
      75658:data<=16'd6619;
      75659:data<=16'd5398;
      75660:data<=16'd5917;
      75661:data<=16'd5306;
      75662:data<=16'd4707;
      75663:data<=16'd8919;
      75664:data<=16'd7626;
      75665:data<=-16'd3148;
      75666:data<=-16'd8530;
      75667:data<=-16'd6977;
      75668:data<=-16'd7436;
      75669:data<=-16'd7263;
      75670:data<=-16'd5053;
      75671:data<=-16'd4748;
      75672:data<=-16'd5002;
      75673:data<=-16'd4632;
      75674:data<=-16'd4689;
      75675:data<=-16'd4400;
      75676:data<=-16'd4284;
      75677:data<=-16'd4825;
      75678:data<=-16'd4540;
      75679:data<=-16'd3997;
      75680:data<=-16'd4070;
      75681:data<=-16'd3613;
      75682:data<=-16'd2626;
      75683:data<=-16'd1967;
      75684:data<=-16'd1792;
      75685:data<=-16'd1528;
      75686:data<=-16'd875;
      75687:data<=-16'd1064;
      75688:data<=-16'd1507;
      75689:data<=-16'd1033;
      75690:data<=-16'd1054;
      75691:data<=-16'd922;
      75692:data<=-16'd684;
      75693:data<=-16'd1789;
      75694:data<=-16'd1222;
      75695:data<=16'd305;
      75696:data<=-16'd115;
      75697:data<=-16'd29;
      75698:data<=16'd2;
      75699:data<=16'd305;
      75700:data<=16'd1001;
      75701:data<=-16'd1688;
      75702:data<=16'd1768;
      75703:data<=16'd13725;
      75704:data<=16'd16472;
      75705:data<=16'd13016;
      75706:data<=16'd13723;
      75707:data<=16'd11267;
      75708:data<=16'd8950;
      75709:data<=16'd10433;
      75710:data<=16'd8912;
      75711:data<=16'd8153;
      75712:data<=16'd8718;
      75713:data<=16'd6922;
      75714:data<=16'd6942;
      75715:data<=16'd7056;
      75716:data<=16'd5551;
      75717:data<=16'd5183;
      75718:data<=16'd4631;
      75719:data<=16'd4522;
      75720:data<=16'd4282;
      75721:data<=16'd2837;
      75722:data<=16'd2763;
      75723:data<=16'd2466;
      75724:data<=16'd1838;
      75725:data<=16'd1870;
      75726:data<=16'd572;
      75727:data<=16'd443;
      75728:data<=16'd593;
      75729:data<=-16'd711;
      75730:data<=16'd199;
      75731:data<=16'd82;
      75732:data<=-16'd2011;
      75733:data<=-16'd2144;
      75734:data<=-16'd2776;
      75735:data<=-16'd2951;
      75736:data<=-16'd2787;
      75737:data<=-16'd4223;
      75738:data<=-16'd2508;
      75739:data<=-16'd3891;
      75740:data<=-16'd13894;
      75741:data<=-16'd19761;
      75742:data<=-16'd18155;
      75743:data<=-16'd16929;
      75744:data<=-16'd17258;
      75745:data<=-16'd18228;
      75746:data<=-16'd18333;
      75747:data<=-16'd17617;
      75748:data<=-16'd17091;
      75749:data<=-16'd16072;
      75750:data<=-16'd16446;
      75751:data<=-16'd15729;
      75752:data<=-16'd11282;
      75753:data<=-16'd9336;
      75754:data<=-16'd10069;
      75755:data<=-16'd9304;
      75756:data<=-16'd9412;
      75757:data<=-16'd10226;
      75758:data<=-16'd10088;
      75759:data<=-16'd9891;
      75760:data<=-16'd9160;
      75761:data<=-16'd8523;
      75762:data<=-16'd8291;
      75763:data<=-16'd7595;
      75764:data<=-16'd7503;
      75765:data<=-16'd7488;
      75766:data<=-16'd6576;
      75767:data<=-16'd6325;
      75768:data<=-16'd6419;
      75769:data<=-16'd6448;
      75770:data<=-16'd8037;
      75771:data<=-16'd8746;
      75772:data<=-16'd7277;
      75773:data<=-16'd7595;
      75774:data<=-16'd7507;
      75775:data<=-16'd6190;
      75776:data<=-16'd8047;
      75777:data<=-16'd3988;
      75778:data<=16'd7877;
      75779:data<=16'd10601;
      75780:data<=16'd7321;
      75781:data<=16'd8715;
      75782:data<=16'd7533;
      75783:data<=16'd5207;
      75784:data<=16'd6037;
      75785:data<=16'd4819;
      75786:data<=16'd4137;
      75787:data<=16'd5002;
      75788:data<=16'd4282;
      75789:data<=16'd4296;
      75790:data<=16'd4111;
      75791:data<=16'd3436;
      75792:data<=16'd3494;
      75793:data<=16'd2582;
      75794:data<=16'd2540;
      75795:data<=16'd2149;
      75796:data<=-16'd1154;
      75797:data<=-16'd3536;
      75798:data<=-16'd4314;
      75799:data<=-16'd4563;
      75800:data<=-16'd4144;
      75801:data<=-16'd4209;
      75802:data<=-16'd3591;
      75803:data<=-16'd3585;
      75804:data<=-16'd4848;
      75805:data<=-16'd4034;
      75806:data<=-16'd3386;
      75807:data<=-16'd4631;
      75808:data<=-16'd5935;
      75809:data<=-16'd6787;
      75810:data<=-16'd5348;
      75811:data<=-16'd5093;
      75812:data<=-16'd7181;
      75813:data<=-16'd4943;
      75814:data<=-16'd4977;
      75815:data<=-16'd13734;
      75816:data<=-16'd19766;
      75817:data<=-16'd19115;
      75818:data<=-16'd18116;
      75819:data<=-16'd17851;
      75820:data<=-16'd18290;
      75821:data<=-16'd18575;
      75822:data<=-16'd17667;
      75823:data<=-16'd17106;
      75824:data<=-16'd16539;
      75825:data<=-16'd15386;
      75826:data<=-16'd14600;
      75827:data<=-16'd14116;
      75828:data<=-16'd13559;
      75829:data<=-16'd12812;
      75830:data<=-16'd12126;
      75831:data<=-16'd11768;
      75832:data<=-16'd11805;
      75833:data<=-16'd12334;
      75834:data<=-16'd11997;
      75835:data<=-16'd10495;
      75836:data<=-16'd9865;
      75837:data<=-16'd9505;
      75838:data<=-16'd8455;
      75839:data<=-16'd8449;
      75840:data<=-16'd7594;
      75841:data<=-16'd4046;
      75842:data<=-16'd2449;
      75843:data<=-16'd3146;
      75844:data<=-16'd2594;
      75845:data<=-16'd3398;
      75846:data<=-16'd4522;
      75847:data<=-16'd3206;
      75848:data<=-16'd3298;
      75849:data<=-16'd2552;
      75850:data<=-16'd902;
      75851:data<=-16'd3554;
      75852:data<=16'd185;
      75853:data<=16'd12196;
      75854:data<=16'd14973;
      75855:data<=16'd11808;
      75856:data<=16'd12989;
      75857:data<=16'd12190;
      75858:data<=16'd10069;
      75859:data<=16'd10279;
      75860:data<=16'd9464;
      75861:data<=16'd9016;
      75862:data<=16'd9473;
      75863:data<=16'd8933;
      75864:data<=16'd8496;
      75865:data<=16'd8072;
      75866:data<=16'd7797;
      75867:data<=16'd7870;
      75868:data<=16'd7579;
      75869:data<=16'd7228;
      75870:data<=16'd5918;
      75871:data<=16'd4563;
      75872:data<=16'd4955;
      75873:data<=16'd4928;
      75874:data<=16'd4000;
      75875:data<=16'd3676;
      75876:data<=16'd3563;
      75877:data<=16'd3701;
      75878:data<=16'd3475;
      75879:data<=16'd2372;
      75880:data<=16'd2182;
      75881:data<=16'd3011;
      75882:data<=16'd2620;
      75883:data<=16'd1090;
      75884:data<=16'd737;
      75885:data<=16'd314;
      75886:data<=-16'd2717;
      75887:data<=-16'd4332;
      75888:data<=-16'd2184;
      75889:data<=-16'd3761;
      75890:data<=-16'd11943;
      75891:data<=-16'd17816;
      75892:data<=-16'd17111;
      75893:data<=-16'd15832;
      75894:data<=-16'd16442;
      75895:data<=-16'd16407;
      75896:data<=-16'd16161;
      75897:data<=-16'd15925;
      75898:data<=-16'd15038;
      75899:data<=-16'd14375;
      75900:data<=-16'd13488;
      75901:data<=-16'd12692;
      75902:data<=-16'd12295;
      75903:data<=-16'd11122;
      75904:data<=-16'd10683;
      75905:data<=-16'd10710;
      75906:data<=-16'd9621;
      75907:data<=-16'd9838;
      75908:data<=-16'd10983;
      75909:data<=-16'd10725;
      75910:data<=-16'd9539;
      75911:data<=-16'd7955;
      75912:data<=-16'd7398;
      75913:data<=-16'd7338;
      75914:data<=-16'd6300;
      75915:data<=-16'd5708;
      75916:data<=-16'd4814;
      75917:data<=-16'd4090;
      75918:data<=-16'd4720;
      75919:data<=-16'd4047;
      75920:data<=-16'd3471;
      75921:data<=-16'd3503;
      75922:data<=-16'd2525;
      75923:data<=-16'd3104;
      75924:data<=-16'd2049;
      75925:data<=-16'd338;
      75926:data<=-16'd3090;
      75927:data<=16'd1092;
      75928:data<=16'd12854;
      75929:data<=16'd16771;
      75930:data<=16'd16856;
      75931:data<=16'd18810;
      75932:data<=16'd18240;
      75933:data<=16'd18647;
      75934:data<=16'd19664;
      75935:data<=16'd18471;
      75936:data<=16'd18333;
      75937:data<=16'd17893;
      75938:data<=16'd16756;
      75939:data<=16'd16798;
      75940:data<=16'd16404;
      75941:data<=16'd16267;
      75942:data<=16'd16066;
      75943:data<=16'd14815;
      75944:data<=16'd14839;
      75945:data<=16'd15685;
      75946:data<=16'd15934;
      75947:data<=16'd15494;
      75948:data<=16'd14336;
      75949:data<=16'd13858;
      75950:data<=16'd13371;
      75951:data<=16'd12240;
      75952:data<=16'd11931;
      75953:data<=16'd11621;
      75954:data<=16'd11148;
      75955:data<=16'd10681;
      75956:data<=16'd9547;
      75957:data<=16'd10029;
      75958:data<=16'd11667;
      75959:data<=16'd11561;
      75960:data<=16'd11129;
      75961:data<=16'd10627;
      75962:data<=16'd9459;
      75963:data<=16'd10078;
      75964:data<=16'd9186;
      75965:data<=16'd1309;
      75966:data<=-16'd6657;
      75967:data<=-16'd6801;
      75968:data<=-16'd5174;
      75969:data<=-16'd5905;
      75970:data<=-16'd4616;
      75971:data<=-16'd2981;
      75972:data<=-16'd3219;
      75973:data<=-16'd2601;
      75974:data<=-16'd3168;
      75975:data<=-16'd6137;
      75976:data<=-16'd7474;
      75977:data<=-16'd6675;
      75978:data<=-16'd6072;
      75979:data<=-16'd6203;
      75980:data<=-16'd6228;
      75981:data<=-16'd5932;
      75982:data<=-16'd5347;
      75983:data<=-16'd3541;
      75984:data<=-16'd2103;
      75985:data<=-16'd2120;
      75986:data<=-16'd1374;
      75987:data<=-16'd925;
      75988:data<=-16'd1300;
      75989:data<=-16'd723;
      75990:data<=-16'd802;
      75991:data<=-16'd952;
      75992:data<=-16'd12;
      75993:data<=-16'd3;
      75994:data<=-16'd70;
      75995:data<=16'd544;
      75996:data<=16'd1697;
      75997:data<=16'd2654;
      75998:data<=16'd1339;
      75999:data<=16'd1741;
      76000:data<=16'd3113;
      76001:data<=16'd578;
      76002:data<=16'd4393;
      76003:data<=16'd15450;
      76004:data<=16'd18257;
      76005:data<=16'd15835;
      76006:data<=16'd16045;
      76007:data<=16'd15632;
      76008:data<=16'd16380;
      76009:data<=16'd17239;
      76010:data<=16'd15359;
      76011:data<=16'd15086;
      76012:data<=16'd15488;
      76013:data<=16'd14371;
      76014:data<=16'd13675;
      76015:data<=16'd12939;
      76016:data<=16'd12669;
      76017:data<=16'd12242;
      76018:data<=16'd11235;
      76019:data<=16'd13027;
      76020:data<=16'd15594;
      76021:data<=16'd16057;
      76022:data<=16'd15901;
      76023:data<=16'd14560;
      76024:data<=16'd13479;
      76025:data<=16'd13647;
      76026:data<=16'd12521;
      76027:data<=16'd11658;
      76028:data<=16'd11477;
      76029:data<=16'd10340;
      76030:data<=16'd10037;
      76031:data<=16'd9861;
      76032:data<=16'd9589;
      76033:data<=16'd10602;
      76034:data<=16'd10451;
      76035:data<=16'd9938;
      76036:data<=16'd9887;
      76037:data<=16'd7768;
      76038:data<=16'd7360;
      76039:data<=16'd7450;
      76040:data<=-16'd262;
      76041:data<=-16'd9138;
      76042:data<=-16'd9414;
      76043:data<=-16'd7459;
      76044:data<=-16'd8182;
      76045:data<=-16'd7473;
      76046:data<=-16'd5553;
      76047:data<=-16'd5198;
      76048:data<=-16'd5454;
      76049:data<=-16'd5582;
      76050:data<=-16'd5964;
      76051:data<=-16'd5952;
      76052:data<=-16'd5582;
      76053:data<=-16'd5557;
      76054:data<=-16'd5547;
      76055:data<=-16'd5266;
      76056:data<=-16'd4940;
      76057:data<=-16'd4622;
      76058:data<=-16'd3903;
      76059:data<=-16'd2538;
      76060:data<=-16'd1932;
      76061:data<=-16'd2541;
      76062:data<=-16'd2590;
      76063:data<=-16'd3054;
      76064:data<=-16'd5424;
      76065:data<=-16'd6995;
      76066:data<=-16'd6734;
      76067:data<=-16'd6560;
      76068:data<=-16'd6156;
      76069:data<=-16'd5503;
      76070:data<=-16'd5234;
      76071:data<=-16'd4034;
      76072:data<=-16'd3339;
      76073:data<=-16'd4469;
      76074:data<=-16'd3523;
      76075:data<=-16'd2469;
      76076:data<=-16'd4958;
      76077:data<=-16'd1441;
      76078:data<=16'd9632;
      76079:data<=16'd13490;
      76080:data<=16'd10563;
      76081:data<=16'd10633;
      76082:data<=16'd10863;
      76083:data<=16'd10513;
      76084:data<=16'd11588;
      76085:data<=16'd10780;
      76086:data<=16'd9815;
      76087:data<=16'd9850;
      76088:data<=16'd8655;
      76089:data<=16'd8719;
      76090:data<=16'd9145;
      76091:data<=16'd7686;
      76092:data<=16'd7107;
      76093:data<=16'd6892;
      76094:data<=16'd6128;
      76095:data<=16'd6343;
      76096:data<=16'd6748;
      76097:data<=16'd7045;
      76098:data<=16'd6702;
      76099:data<=16'd5529;
      76100:data<=16'd5109;
      76101:data<=16'd4491;
      76102:data<=16'd3897;
      76103:data<=16'd4027;
      76104:data<=16'd3274;
      76105:data<=16'd3151;
      76106:data<=16'd2974;
      76107:data<=16'd1888;
      76108:data<=16'd4572;
      76109:data<=16'd8096;
      76110:data<=16'd7993;
      76111:data<=16'd7659;
      76112:data<=16'd6304;
      76113:data<=16'd5236;
      76114:data<=16'd5742;
      76115:data<=-16'd943;
      76116:data<=-16'd10420;
      76117:data<=-16'd10915;
      76118:data<=-16'd9209;
      76119:data<=-16'd10357;
      76120:data<=-16'd9655;
      76121:data<=-16'd8777;
      76122:data<=-16'd8995;
      76123:data<=-16'd8937;
      76124:data<=-16'd9247;
      76125:data<=-16'd9338;
      76126:data<=-16'd9392;
      76127:data<=-16'd9351;
      76128:data<=-16'd8771;
      76129:data<=-16'd9006;
      76130:data<=-16'd9019;
      76131:data<=-16'd8190;
      76132:data<=-16'd8106;
      76133:data<=-16'd8577;
      76134:data<=-16'd9454;
      76135:data<=-16'd9491;
      76136:data<=-16'd8325;
      76137:data<=-16'd8552;
      76138:data<=-16'd8727;
      76139:data<=-16'd7982;
      76140:data<=-16'd8338;
      76141:data<=-16'd8026;
      76142:data<=-16'd7759;
      76143:data<=-16'd8290;
      76144:data<=-16'd6983;
      76145:data<=-16'd7013;
      76146:data<=-16'd8664;
      76147:data<=-16'd8270;
      76148:data<=-16'd8560;
      76149:data<=-16'd8373;
      76150:data<=-16'd7028;
      76151:data<=-16'd8395;
      76152:data<=-16'd5492;
      76153:data<=16'd2754;
      76154:data<=16'd4702;
      76155:data<=16'd2758;
      76156:data<=16'd3600;
      76157:data<=16'd3475;
      76158:data<=16'd1988;
      76159:data<=16'd931;
      76160:data<=16'd227;
      76161:data<=16'd614;
      76162:data<=16'd484;
      76163:data<=-16'd103;
      76164:data<=16'd256;
      76165:data<=16'd42;
      76166:data<=-16'd346;
      76167:data<=-16'd379;
      76168:data<=-16'd887;
      76169:data<=-16'd423;
      76170:data<=-16'd8;
      76171:data<=-16'd1551;
      76172:data<=-16'd2513;
      76173:data<=-16'd2229;
      76174:data<=-16'd2564;
      76175:data<=-16'd2943;
      76176:data<=-16'd3036;
      76177:data<=-16'd3154;
      76178:data<=-16'd2917;
      76179:data<=-16'd2877;
      76180:data<=-16'd3063;
      76181:data<=-16'd3078;
      76182:data<=-16'd3348;
      76183:data<=-16'd3812;
      76184:data<=-16'd4763;
      76185:data<=-16'd5450;
      76186:data<=-16'd5150;
      76187:data<=-16'd5958;
      76188:data<=-16'd5494;
      76189:data<=-16'd3488;
      76190:data<=-16'd9347;
      76191:data<=-16'd18885;
      76192:data<=-16'd19578;
      76193:data<=-16'd17531;
      76194:data<=-16'd18004;
      76195:data<=-16'd17268;
      76196:data<=-16'd18001;
      76197:data<=-16'd17411;
      76198:data<=-16'd13124;
      76199:data<=-16'd12063;
      76200:data<=-16'd12151;
      76201:data<=-16'd10715;
      76202:data<=-16'd11253;
      76203:data<=-16'd10863;
      76204:data<=-16'd9562;
      76205:data<=-16'd9935;
      76206:data<=-16'd9477;
      76207:data<=-16'd8778;
      76208:data<=-16'd8837;
      76209:data<=-16'd9274;
      76210:data<=-16'd10002;
      76211:data<=-16'd9119;
      76212:data<=-16'd8443;
      76213:data<=-16'd8520;
      76214:data<=-16'd7191;
      76215:data<=-16'd7047;
      76216:data<=-16'd7228;
      76217:data<=-16'd6249;
      76218:data<=-16'd6361;
      76219:data<=-16'd5444;
      76220:data<=-16'd4833;
      76221:data<=-16'd6388;
      76222:data<=-16'd6475;
      76223:data<=-16'd6546;
      76224:data<=-16'd5896;
      76225:data<=-16'd4272;
      76226:data<=-16'd6482;
      76227:data<=-16'd3506;
      76228:data<=16'd8019;
      76229:data<=16'd12528;
      76230:data<=16'd10107;
      76231:data<=16'd10302;
      76232:data<=16'd10566;
      76233:data<=16'd9370;
      76234:data<=16'd7896;
      76235:data<=16'd6748;
      76236:data<=16'd7321;
      76237:data<=16'd7624;
      76238:data<=16'd7072;
      76239:data<=16'd7078;
      76240:data<=16'd7045;
      76241:data<=16'd6369;
      76242:data<=16'd4046;
      76243:data<=16'd1842;
      76244:data<=16'd2276;
      76245:data<=16'd2177;
      76246:data<=16'd450;
      76247:data<=-16'd17;
      76248:data<=16'd221;
      76249:data<=16'd132;
      76250:data<=16'd212;
      76251:data<=16'd176;
      76252:data<=16'd39;
      76253:data<=16'd23;
      76254:data<=-16'd126;
      76255:data<=-16'd370;
      76256:data<=-16'd426;
      76257:data<=-16'd464;
      76258:data<=-16'd1116;
      76259:data<=-16'd2408;
      76260:data<=-16'd2766;
      76261:data<=-16'd1806;
      76262:data<=-16'd2167;
      76263:data<=-16'd2450;
      76264:data<=-16'd1098;
      76265:data<=-16'd5938;
      76266:data<=-16'd15499;
      76267:data<=-16'd17044;
      76268:data<=-16'd14509;
      76269:data<=-16'd15421;
      76270:data<=-16'd14900;
      76271:data<=-16'd14219;
      76272:data<=-16'd15080;
      76273:data<=-16'd14035;
      76274:data<=-16'd13784;
      76275:data<=-16'd13923;
      76276:data<=-16'd12502;
      76277:data<=-16'd12339;
      76278:data<=-16'd11539;
      76279:data<=-16'd9700;
      76280:data<=-16'd9582;
      76281:data<=-16'd9506;
      76282:data<=-16'd9379;
      76283:data<=-16'd9632;
      76284:data<=-16'd9777;
      76285:data<=-16'd10393;
      76286:data<=-16'd8639;
      76287:data<=-16'd4901;
      76288:data<=-16'd3554;
      76289:data<=-16'd3421;
      76290:data<=-16'd2535;
      76291:data<=-16'd1597;
      76292:data<=-16'd1295;
      76293:data<=-16'd1604;
      76294:data<=-16'd1095;
      76295:data<=-16'd726;
      76296:data<=-16'd1500;
      76297:data<=-16'd1949;
      76298:data<=-16'd2033;
      76299:data<=-16'd590;
      76300:data<=16'd259;
      76301:data<=-16'd2341;
      76302:data<=16'd984;
      76303:data<=16'd12116;
      76304:data<=16'd16581;
      76305:data<=16'd13787;
      76306:data<=16'd13511;
      76307:data<=16'd14231;
      76308:data<=16'd13071;
      76309:data<=16'd11775;
      76310:data<=16'd10784;
      76311:data<=16'd10363;
      76312:data<=16'd10460;
      76313:data<=16'd10586;
      76314:data<=16'd10655;
      76315:data<=16'd10187;
      76316:data<=16'd9717;
      76317:data<=16'd9909;
      76318:data<=16'd9832;
      76319:data<=16'd9442;
      76320:data<=16'd9298;
      76321:data<=16'd9051;
      76322:data<=16'd9144;
      76323:data<=16'd9309;
      76324:data<=16'd8452;
      76325:data<=16'd7664;
      76326:data<=16'd7626;
      76327:data<=16'd7735;
      76328:data<=16'd7906;
      76329:data<=16'd7523;
      76330:data<=16'd6804;
      76331:data<=16'd5057;
      76332:data<=16'd1994;
      76333:data<=16'd2012;
      76334:data<=16'd3990;
      76335:data<=16'd3582;
      76336:data<=16'd3755;
      76337:data<=16'd3565;
      76338:data<=16'd2978;
      76339:data<=16'd5379;
      76340:data<=16'd745;
      76341:data<=-16'd10322;
      76342:data<=-16'd11591;
      76343:data<=-16'd8878;
      76344:data<=-16'd11004;
      76345:data<=-16'd10437;
      76346:data<=-16'd8100;
      76347:data<=-16'd7110;
      76348:data<=-16'd5874;
      76349:data<=-16'd6234;
      76350:data<=-16'd6099;
      76351:data<=-16'd4931;
      76352:data<=-16'd5051;
      76353:data<=-16'd4454;
      76354:data<=-16'd4135;
      76355:data<=-16'd4441;
      76356:data<=-16'd3803;
      76357:data<=-16'd4158;
      76358:data<=-16'd3703;
      76359:data<=-16'd1691;
      76360:data<=-16'd1168;
      76361:data<=-16'd907;
      76362:data<=-16'd537;
      76363:data<=-16'd417;
      76364:data<=16'd76;
      76365:data<=-16'd271;
      76366:data<=16'd196;
      76367:data<=16'd1186;
      76368:data<=16'd749;
      76369:data<=16'd1278;
      76370:data<=16'd1433;
      76371:data<=16'd1365;
      76372:data<=16'd3720;
      76373:data<=16'd3632;
      76374:data<=16'd2635;
      76375:data<=16'd4968;
      76376:data<=16'd5680;
      76377:data<=16'd9523;
      76378:data<=16'd19681;
      76379:data<=16'd23238;
      76380:data<=16'd20613;
      76381:data<=16'd21038;
      76382:data<=16'd20588;
      76383:data<=16'd19141;
      76384:data<=16'd20510;
      76385:data<=16'd20492;
      76386:data<=16'd19062;
      76387:data<=16'd19144;
      76388:data<=16'd18553;
      76389:data<=16'd17358;
      76390:data<=16'd16797;
      76391:data<=16'd15960;
      76392:data<=16'd15303;
      76393:data<=16'd14810;
      76394:data<=16'd14128;
      76395:data<=16'd13800;
      76396:data<=16'd13878;
      76397:data<=16'd14600;
      76398:data<=16'd14587;
      76399:data<=16'd13367;
      76400:data<=16'd13154;
      76401:data<=16'd12737;
      76402:data<=16'd11799;
      76403:data<=16'd11940;
      76404:data<=16'd10675;
      76405:data<=16'd9257;
      76406:data<=16'd9438;
      76407:data<=16'd8331;
      76408:data<=16'd8288;
      76409:data<=16'd9468;
      76410:data<=16'd9239;
      76411:data<=16'd10011;
      76412:data<=16'd8708;
      76413:data<=16'd6966;
      76414:data<=16'd9674;
      76415:data<=16'd4723;
      76416:data<=-16'd7244;
      76417:data<=-16'd9359;
      76418:data<=-16'd6680;
      76419:data<=-16'd7662;
      76420:data<=-16'd9163;
      76421:data<=-16'd11229;
      76422:data<=-16'd10393;
      76423:data<=-16'd7413;
      76424:data<=-16'd8211;
      76425:data<=-16'd8448;
      76426:data<=-16'd7250;
      76427:data<=-16'd7783;
      76428:data<=-16'd7321;
      76429:data<=-16'd7012;
      76430:data<=-16'd7124;
      76431:data<=-16'd6200;
      76432:data<=-16'd6880;
      76433:data<=-16'd6902;
      76434:data<=-16'd4881;
      76435:data<=-16'd4253;
      76436:data<=-16'd4152;
      76437:data<=-16'd3882;
      76438:data<=-16'd3876;
      76439:data<=-16'd3610;
      76440:data<=-16'd3961;
      76441:data<=-16'd3842;
      76442:data<=-16'd3403;
      76443:data<=-16'd3627;
      76444:data<=-16'd2895;
      76445:data<=-16'd2939;
      76446:data<=-16'd3183;
      76447:data<=-16'd990;
      76448:data<=-16'd487;
      76449:data<=-16'd948;
      76450:data<=16'd59;
      76451:data<=-16'd1580;
      76452:data<=16'd497;
      76453:data<=16'd10470;
      76454:data<=16'd14974;
      76455:data<=16'd12534;
      76456:data<=16'd12657;
      76457:data<=16'd12393;
      76458:data<=16'd11209;
      76459:data<=16'd12957;
      76460:data<=16'd13019;
      76461:data<=16'd11274;
      76462:data<=16'd11209;
      76463:data<=16'd10146;
      76464:data<=16'd9491;
      76465:data<=16'd11797;
      76466:data<=16'd13282;
      76467:data<=16'd12783;
      76468:data<=16'd11999;
      76469:data<=16'd11198;
      76470:data<=16'd10945;
      76471:data<=16'd11470;
      76472:data<=16'd12257;
      76473:data<=16'd11770;
      76474:data<=16'd10129;
      76475:data<=16'd9717;
      76476:data<=16'd9635;
      76477:data<=16'd9292;
      76478:data<=16'd9154;
      76479:data<=16'd7321;
      76480:data<=16'd6244;
      76481:data<=16'd6830;
      76482:data<=16'd5483;
      76483:data<=16'd5121;
      76484:data<=16'd6176;
      76485:data<=16'd5982;
      76486:data<=16'd6761;
      76487:data<=16'd5289;
      76488:data<=16'd3331;
      76489:data<=16'd6156;
      76490:data<=16'd1782;
      76491:data<=-16'd9835;
      76492:data<=-16'd11940;
      76493:data<=-16'd9620;
      76494:data<=-16'd11192;
      76495:data<=-16'd10660;
      76496:data<=-16'd8900;
      76497:data<=-16'd8146;
      76498:data<=-16'd7315;
      76499:data<=-16'd7691;
      76500:data<=-16'd7582;
      76501:data<=-16'd6895;
      76502:data<=-16'd6921;
      76503:data<=-16'd6619;
      76504:data<=-16'd7062;
      76505:data<=-16'd7403;
      76506:data<=-16'd6874;
      76507:data<=-16'd7033;
      76508:data<=-16'd6319;
      76509:data<=-16'd6435;
      76510:data<=-16'd8956;
      76511:data<=-16'd9421;
      76512:data<=-16'd8577;
      76513:data<=-16'd8740;
      76514:data<=-16'd8287;
      76515:data<=-16'd8140;
      76516:data<=-16'd8204;
      76517:data<=-16'd7970;
      76518:data<=-16'd8055;
      76519:data<=-16'd6959;
      76520:data<=-16'd6440;
      76521:data<=-16'd7213;
      76522:data<=-16'd6725;
      76523:data<=-16'd6775;
      76524:data<=-16'd6340;
      76525:data<=-16'd4992;
      76526:data<=-16'd7127;
      76527:data<=-16'd5400;
      76528:data<=16'd4643;
      76529:data<=16'd9687;
      76530:data<=16'd7365;
      76531:data<=16'd6890;
      76532:data<=16'd7288;
      76533:data<=16'd6623;
      76534:data<=16'd5706;
      76535:data<=16'd3386;
      76536:data<=16'd2308;
      76537:data<=16'd3125;
      76538:data<=16'd2664;
      76539:data<=16'd2137;
      76540:data<=16'd2193;
      76541:data<=16'd1504;
      76542:data<=16'd1375;
      76543:data<=16'd1492;
      76544:data<=16'd1357;
      76545:data<=16'd1986;
      76546:data<=16'd1307;
      76547:data<=-16'd836;
      76548:data<=-16'd1445;
      76549:data<=-16'd1412;
      76550:data<=-16'd2012;
      76551:data<=-16'd2056;
      76552:data<=-16'd1732;
      76553:data<=-16'd1450;
      76554:data<=-16'd329;
      76555:data<=16'd1635;
      76556:data<=16'd2143;
      76557:data<=16'd1130;
      76558:data<=16'd1606;
      76559:data<=16'd1254;
      76560:data<=-16'd1199;
      76561:data<=-16'd1122;
      76562:data<=-16'd1202;
      76563:data<=-16'd2165;
      76564:data<=16'd106;
      76565:data<=-16'd4214;
      76566:data<=-16'd15414;
      76567:data<=-16'd17164;
      76568:data<=-16'd14296;
      76569:data<=-16'd15963;
      76570:data<=-16'd15092;
      76571:data<=-16'd13963;
      76572:data<=-16'd15855;
      76573:data<=-16'd15318;
      76574:data<=-16'd14439;
      76575:data<=-16'd14522;
      76576:data<=-16'd13411;
      76577:data<=-16'd12950;
      76578:data<=-16'd12621;
      76579:data<=-16'd12066;
      76580:data<=-16'd11856;
      76581:data<=-16'd11059;
      76582:data<=-16'd10710;
      76583:data<=-16'd10199;
      76584:data<=-16'd10196;
      76585:data<=-16'd12234;
      76586:data<=-16'd12196;
      76587:data<=-16'd10569;
      76588:data<=-16'd10766;
      76589:data<=-16'd10686;
      76590:data<=-16'd10522;
      76591:data<=-16'd10005;
      76592:data<=-16'd8316;
      76593:data<=-16'd8125;
      76594:data<=-16'd7632;
      76595:data<=-16'd6748;
      76596:data<=-16'd7529;
      76597:data<=-16'd7201;
      76598:data<=-16'd8564;
      76599:data<=-16'd11905;
      76600:data<=-16'd11726;
      76601:data<=-16'd11926;
      76602:data<=-16'd10117;
      76603:data<=-16'd643;
      76604:data<=16'd5010;
      76605:data<=16'd3751;
      76606:data<=16'd4478;
      76607:data<=16'd4887;
      76608:data<=16'd4005;
      76609:data<=16'd3958;
      76610:data<=16'd1908;
      76611:data<=16'd549;
      76612:data<=16'd1513;
      76613:data<=16'd1451;
      76614:data<=16'd1387;
      76615:data<=16'd1433;
      76616:data<=16'd1051;
      76617:data<=16'd1809;
      76618:data<=16'd1861;
      76619:data<=16'd1216;
      76620:data<=16'd1962;
      76621:data<=16'd2020;
      76622:data<=16'd576;
      76623:data<=-16'd787;
      76624:data<=-16'd1438;
      76625:data<=-16'd1134;
      76626:data<=-16'd902;
      76627:data<=-16'd760;
      76628:data<=-16'd423;
      76629:data<=-16'd1019;
      76630:data<=-16'd1084;
      76631:data<=-16'd632;
      76632:data<=-16'd1287;
      76633:data<=-16'd687;
      76634:data<=-16'd226;
      76635:data<=-16'd1906;
      76636:data<=-16'd2077;
      76637:data<=-16'd2440;
      76638:data<=-16'd2940;
      76639:data<=-16'd105;
      76640:data<=-16'd3560;
      76641:data<=-16'd14730;
      76642:data<=-16'd17749;
      76643:data<=-16'd12969;
      76644:data<=-16'd10420;
      76645:data<=-16'd9060;
      76646:data<=-16'd8681;
      76647:data<=-16'd9626;
      76648:data<=-16'd9320;
      76649:data<=-16'd8893;
      76650:data<=-16'd8584;
      76651:data<=-16'd7881;
      76652:data<=-16'd7656;
      76653:data<=-16'd7036;
      76654:data<=-16'd6432;
      76655:data<=-16'd6270;
      76656:data<=-16'd5888;
      76657:data<=-16'd5779;
      76658:data<=-16'd5006;
      76659:data<=-16'd4681;
      76660:data<=-16'd6487;
      76661:data<=-16'd6916;
      76662:data<=-16'd5623;
      76663:data<=-16'd5285;
      76664:data<=-16'd4952;
      76665:data<=-16'd4576;
      76666:data<=-16'd4096;
      76667:data<=-16'd3166;
      76668:data<=-16'd2958;
      76669:data<=-16'd2065;
      76670:data<=-16'd1221;
      76671:data<=-16'd2417;
      76672:data<=-16'd3054;
      76673:data<=-16'd3313;
      76674:data<=-16'd3574;
      76675:data<=-16'd2563;
      76676:data<=-16'd3391;
      76677:data<=-16'd1495;
      76678:data<=16'd8046;
      76679:data<=16'd13793;
      76680:data<=16'd12000;
      76681:data<=16'd11741;
      76682:data<=16'd12452;
      76683:data<=16'd12020;
      76684:data<=16'd11354;
      76685:data<=16'd9009;
      76686:data<=16'd8034;
      76687:data<=16'd8040;
      76688:data<=16'd5134;
      76689:data<=16'd3582;
      76690:data<=16'd4164;
      76691:data<=16'd3368;
      76692:data<=16'd3594;
      76693:data<=16'd4479;
      76694:data<=16'd4056;
      76695:data<=16'd4144;
      76696:data<=16'd4266;
      76697:data<=16'd3465;
      76698:data<=16'd1974;
      76699:data<=16'd669;
      76700:data<=16'd1169;
      76701:data<=16'd1659;
      76702:data<=16'd1571;
      76703:data<=16'd2196;
      76704:data<=16'd1651;
      76705:data<=16'd1448;
      76706:data<=16'd2391;
      76707:data<=16'd1814;
      76708:data<=16'd2391;
      76709:data<=16'd2992;
      76710:data<=16'd687;
      76711:data<=16'd331;
      76712:data<=16'd535;
      76713:data<=16'd105;
      76714:data<=16'd2655;
      76715:data<=-16'd1230;
      76716:data<=-16'd12236;
      76717:data<=-16'd14651;
      76718:data<=-16'd11499;
      76719:data<=-16'd11950;
      76720:data<=-16'd11159;
      76721:data<=-16'd9755;
      76722:data<=-16'd10390;
      76723:data<=-16'd9345;
      76724:data<=-16'd7639;
      76725:data<=-16'd6953;
      76726:data<=-16'd5999;
      76727:data<=-16'd5556;
      76728:data<=-16'd5477;
      76729:data<=-16'd4893;
      76730:data<=-16'd4663;
      76731:data<=-16'd4595;
      76732:data<=-16'd2742;
      76733:data<=16'd658;
      76734:data<=16'd2303;
      76735:data<=16'd2591;
      76736:data<=16'd4091;
      76737:data<=16'd4696;
      76738:data<=16'd4291;
      76739:data<=16'd5028;
      76740:data<=16'd4833;
      76741:data<=16'd4258;
      76742:data<=16'd5037;
      76743:data<=16'd5147;
      76744:data<=16'd5430;
      76745:data<=16'd5667;
      76746:data<=16'd4269;
      76747:data<=16'd4939;
      76748:data<=16'd7069;
      76749:data<=16'd7339;
      76750:data<=16'd7488;
      76751:data<=16'd6598;
      76752:data<=16'd7632;
      76753:data<=16'd15805;
      76754:data<=16'd21890;
      76755:data<=16'd20497;
      76756:data<=16'd19878;
      76757:data<=16'd19940;
      76758:data<=16'd18164;
      76759:data<=16'd18412;
      76760:data<=16'd19355;
      76761:data<=16'd18988;
      76762:data<=16'd18242;
      76763:data<=16'd16845;
      76764:data<=16'd16378;
      76765:data<=16'd16460;
      76766:data<=16'd15271;
      76767:data<=16'd14552;
      76768:data<=16'd14213;
      76769:data<=16'd13641;
      76770:data<=16'd13402;
      76771:data<=16'd12351;
      76772:data<=16'd12337;
      76773:data<=16'd13737;
      76774:data<=16'd13080;
      76775:data<=16'd12242;
      76776:data<=16'd12038;
      76777:data<=16'd9696;
      76778:data<=16'd7588;
      76779:data<=16'd6884;
      76780:data<=16'd6128;
      76781:data<=16'd5934;
      76782:data<=16'd5439;
      76783:data<=16'd5285;
      76784:data<=16'd6299;
      76785:data<=16'd6707;
      76786:data<=16'd7189;
      76787:data<=16'd6623;
      76788:data<=16'd5752;
      76789:data<=16'd7806;
      76790:data<=16'd4008;
      76791:data<=-16'd7074;
      76792:data<=-16'd10513;
      76793:data<=-16'd8138;
      76794:data<=-16'd8740;
      76795:data<=-16'd7967;
      76796:data<=-16'd6987;
      76797:data<=-16'd7397;
      76798:data<=-16'd4969;
      76799:data<=-16'd2842;
      76800:data<=-16'd2438;
      76801:data<=-16'd1662;
      76802:data<=-16'd1868;
      76803:data<=-16'd1829;
      76804:data<=-16'd1642;
      76805:data<=-16'd2402;
      76806:data<=-16'd2018;
      76807:data<=-16'd1603;
      76808:data<=-16'd1794;
      76809:data<=-16'd1485;
      76810:data<=-16'd1277;
      76811:data<=-16'd6;
      76812:data<=16'd1124;
      76813:data<=16'd593;
      76814:data<=16'd661;
      76815:data<=16'd581;
      76816:data<=16'd246;
      76817:data<=16'd629;
      76818:data<=16'd244;
      76819:data<=16'd406;
      76820:data<=16'd258;
      76821:data<=-16'd238;
      76822:data<=16'd3463;
      76823:data<=16'd6796;
      76824:data<=16'd6337;
      76825:data<=16'd6704;
      76826:data<=16'd5623;
      76827:data<=16'd5796;
      76828:data<=16'd13050;
      76829:data<=16'd18040;
      76830:data<=16'd16698;
      76831:data<=16'd16125;
      76832:data<=16'd15667;
      76833:data<=16'd14025;
      76834:data<=16'd13652;
      76835:data<=16'd13987;
      76836:data<=16'd14063;
      76837:data<=16'd13177;
      76838:data<=16'd11855;
      76839:data<=16'd11494;
      76840:data<=16'd10956;
      76841:data<=16'd10135;
      76842:data<=16'd9817;
      76843:data<=16'd8984;
      76844:data<=16'd8200;
      76845:data<=16'd8096;
      76846:data<=16'd7736;
      76847:data<=16'd7809;
      76848:data<=16'd8375;
      76849:data<=16'd8084;
      76850:data<=16'd7551;
      76851:data<=16'd7242;
      76852:data<=16'd6758;
      76853:data<=16'd6382;
      76854:data<=16'd5416;
      76855:data<=16'd4546;
      76856:data<=16'd4839;
      76857:data<=16'd4226;
      76858:data<=16'd3515;
      76859:data<=16'd4297;
      76860:data<=16'd4576;
      76861:data<=16'd5007;
      76862:data<=16'd4584;
      76863:data<=16'd2963;
      76864:data<=16'd4673;
      76865:data<=16'd2164;
      76866:data<=-16'd9794;
      76867:data<=-16'd16231;
      76868:data<=-16'd14295;
      76869:data<=-16'd14098;
      76870:data<=-16'd13816;
      76871:data<=-16'd12678;
      76872:data<=-16'd12427;
      76873:data<=-16'd10707;
      76874:data<=-16'd9594;
      76875:data<=-16'd9353;
      76876:data<=-16'd8643;
      76877:data<=-16'd9182;
      76878:data<=-16'd9436;
      76879:data<=-16'd9071;
      76880:data<=-16'd9060;
      76881:data<=-16'd8631;
      76882:data<=-16'd8742;
      76883:data<=-16'd8440;
      76884:data<=-16'd8003;
      76885:data<=-16'd8388;
      76886:data<=-16'd6488;
      76887:data<=-16'd4949;
      76888:data<=-16'd6017;
      76889:data<=-16'd5718;
      76890:data<=-16'd5789;
      76891:data<=-16'd6405;
      76892:data<=-16'd5239;
      76893:data<=-16'd5310;
      76894:data<=-16'd5466;
      76895:data<=-16'd5049;
      76896:data<=-16'd6117;
      76897:data<=-16'd5268;
      76898:data<=-16'd3538;
      76899:data<=-16'd3278;
      76900:data<=-16'd2581;
      76901:data<=-16'd3753;
      76902:data<=-16'd3568;
      76903:data<=16'd3341;
      76904:data<=16'd9342;
      76905:data<=16'd9301;
      76906:data<=16'd7937;
      76907:data<=16'd7674;
      76908:data<=16'd7438;
      76909:data<=16'd6228;
      76910:data<=16'd6548;
      76911:data<=16'd9749;
      76912:data<=16'd11000;
      76913:data<=16'd9806;
      76914:data<=16'd9500;
      76915:data<=16'd8734;
      76916:data<=16'd7899;
      76917:data<=16'd8307;
      76918:data<=16'd7495;
      76919:data<=16'd6125;
      76920:data<=16'd6234;
      76921:data<=16'd6323;
      76922:data<=16'd5870;
      76923:data<=16'd5133;
      76924:data<=16'd3993;
      76925:data<=16'd3454;
      76926:data<=16'd3154;
      76927:data<=16'd2899;
      76928:data<=16'd3034;
      76929:data<=16'd2003;
      76930:data<=16'd1140;
      76931:data<=16'd1597;
      76932:data<=16'd785;
      76933:data<=16'd403;
      76934:data<=16'd796;
      76935:data<=-16'd1121;
      76936:data<=-16'd2231;
      76937:data<=-16'd2375;
      76938:data<=-16'd3268;
      76939:data<=-16'd1847;
      76940:data<=-16'd4657;
      76941:data<=-16'd13981;
      76942:data<=-16'd16888;
      76943:data<=-16'd14565;
      76944:data<=-16'd15362;
      76945:data<=-16'd14775;
      76946:data<=-16'd13045;
      76947:data<=-16'd13858;
      76948:data<=-16'd14425;
      76949:data<=-16'd14647;
      76950:data<=-16'd14562;
      76951:data<=-16'd13380;
      76952:data<=-16'd13336;
      76953:data<=-16'd13414;
      76954:data<=-16'd12433;
      76955:data<=-16'd13130;
      76956:data<=-16'd15177;
      76957:data<=-16'd15725;
      76958:data<=-16'd14985;
      76959:data<=-16'd14728;
      76960:data<=-16'd15010;
      76961:data<=-16'd15167;
      76962:data<=-16'd15114;
      76963:data<=-16'd14593;
      76964:data<=-16'd14117;
      76965:data<=-16'd14195;
      76966:data<=-16'd13670;
      76967:data<=-16'd12507;
      76968:data<=-16'd11761;
      76969:data<=-16'd11329;
      76970:data<=-16'd11171;
      76971:data<=-16'd10922;
      76972:data<=-16'd10419;
      76973:data<=-16'd11153;
      76974:data<=-16'd12067;
      76975:data<=-16'd11045;
      76976:data<=-16'd10897;
      76977:data<=-16'd10763;
      76978:data<=-16'd4484;
      76979:data<=16'd2969;
      76980:data<=16'd3604;
      76981:data<=16'd2526;
      76982:data<=16'd3040;
      76983:data<=16'd2478;
      76984:data<=16'd2488;
      76985:data<=16'd2138;
      76986:data<=16'd174;
      76987:data<=-16'd314;
      76988:data<=-16'd132;
      76989:data<=-16'd419;
      76990:data<=-16'd388;
      76991:data<=-16'd506;
      76992:data<=16'd61;
      76993:data<=16'd180;
      76994:data<=-16'd702;
      76995:data<=-16'd255;
      76996:data<=16'd332;
      76997:data<=16'd190;
      76998:data<=-16'd594;
      76999:data<=-16'd1575;
      77000:data<=16'd538;
      77001:data<=16'd2737;
      77002:data<=16'd2423;
      77003:data<=16'd3356;
      77004:data<=16'd2993;
      77005:data<=16'd1651;
      77006:data<=16'd2851;
      77007:data<=16'd2276;
      77008:data<=16'd1729;
      77009:data<=16'd3002;
      77010:data<=16'd1421;
      77011:data<=16'd496;
      77012:data<=16'd417;
      77013:data<=-16'd657;
      77014:data<=16'd1313;
      77015:data<=-16'd1345;
      77016:data<=-16'd10574;
      77017:data<=-16'd13212;
      77018:data<=-16'd11361;
      77019:data<=-16'd11802;
      77020:data<=-16'd10853;
      77021:data<=-16'd9536;
      77022:data<=-16'd9506;
      77023:data<=-16'd9503;
      77024:data<=-16'd10285;
      77025:data<=-16'd10222;
      77026:data<=-16'd9089;
      77027:data<=-16'd9047;
      77028:data<=-16'd8940;
      77029:data<=-16'd8160;
      77030:data<=-16'd7841;
      77031:data<=-16'd7413;
      77032:data<=-16'd6466;
      77033:data<=-16'd5923;
      77034:data<=-16'd5736;
      77035:data<=-16'd5785;
      77036:data<=-16'd6745;
      77037:data<=-16'd7021;
      77038:data<=-16'd5943;
      77039:data<=-16'd5930;
      77040:data<=-16'd6338;
      77041:data<=-16'd5818;
      77042:data<=-16'd5216;
      77043:data<=-16'd4200;
      77044:data<=-16'd4619;
      77045:data<=-16'd7571;
      77046:data<=-16'd8636;
      77047:data<=-16'd7163;
      77048:data<=-16'd7483;
      77049:data<=-16'd8948;
      77050:data<=-16'd8270;
      77051:data<=-16'd7614;
      77052:data<=-16'd7441;
      77053:data<=-16'd1844;
      77054:data<=16'd5867;
      77055:data<=16'd7113;
      77056:data<=16'd6106;
      77057:data<=16'd6601;
      77058:data<=16'd5871;
      77059:data<=16'd5880;
      77060:data<=16'd5620;
      77061:data<=16'd3495;
      77062:data<=16'd3196;
      77063:data<=16'd3642;
      77064:data<=16'd3333;
      77065:data<=16'd3445;
      77066:data<=16'd3266;
      77067:data<=16'd3880;
      77068:data<=16'd4514;
      77069:data<=16'd3733;
      77070:data<=16'd3418;
      77071:data<=16'd3245;
      77072:data<=16'd3471;
      77073:data<=16'd3551;
      77074:data<=16'd1736;
      77075:data<=16'd1677;
      77076:data<=16'd2681;
      77077:data<=16'd1962;
      77078:data<=16'd2494;
      77079:data<=16'd2614;
      77080:data<=16'd2223;
      77081:data<=16'd3513;
      77082:data<=16'd2549;
      77083:data<=16'd1864;
      77084:data<=16'd3204;
      77085:data<=16'd2143;
      77086:data<=16'd1809;
      77087:data<=16'd1125;
      77088:data<=-16'd338;
      77089:data<=16'd4200;
      77090:data<=16'd4702;
      77091:data<=-16'd4262;
      77092:data<=-16'd7699;
      77093:data<=-16'd5839;
      77094:data<=-16'd6169;
      77095:data<=-16'd5506;
      77096:data<=-16'd5080;
      77097:data<=-16'd4978;
      77098:data<=-16'd3880;
      77099:data<=-16'd5251;
      77100:data<=-16'd6035;
      77101:data<=-16'd4498;
      77102:data<=-16'd4637;
      77103:data<=-16'd4337;
      77104:data<=-16'd2946;
      77105:data<=-16'd3054;
      77106:data<=-16'd2663;
      77107:data<=-16'd1956;
      77108:data<=-16'd2460;
      77109:data<=-16'd2205;
      77110:data<=-16'd1812;
      77111:data<=-16'd2971;
      77112:data<=-16'd3874;
      77113:data<=-16'd3442;
      77114:data<=-16'd2786;
      77115:data<=-16'd2510;
      77116:data<=-16'd2513;
      77117:data<=-16'd2485;
      77118:data<=-16'd1821;
      77119:data<=-16'd628;
      77120:data<=-16'd438;
      77121:data<=-16'd1331;
      77122:data<=-16'd1081;
      77123:data<=-16'd241;
      77124:data<=-16'd335;
      77125:data<=16'd440;
      77126:data<=16'd655;
      77127:data<=-16'd541;
      77128:data<=16'd4200;
      77129:data<=16'd13041;
      77130:data<=16'd14565;
      77131:data<=16'd12138;
      77132:data<=16'd12809;
      77133:data<=16'd11561;
      77134:data<=16'd8169;
      77135:data<=16'd7427;
      77136:data<=16'd7877;
      77137:data<=16'd8269;
      77138:data<=16'd8848;
      77139:data<=16'd8795;
      77140:data<=16'd8449;
      77141:data<=16'd8066;
      77142:data<=16'd7947;
      77143:data<=16'd7953;
      77144:data<=16'd7420;
      77145:data<=16'd7233;
      77146:data<=16'd6881;
      77147:data<=16'd6065;
      77148:data<=16'd7185;
      77149:data<=16'd9248;
      77150:data<=16'd9426;
      77151:data<=16'd8584;
      77152:data<=16'd8498;
      77153:data<=16'd9018;
      77154:data<=16'd8758;
      77155:data<=16'd7953;
      77156:data<=16'd7733;
      77157:data<=16'd7451;
      77158:data<=16'd7356;
      77159:data<=16'd7166;
      77160:data<=16'd6573;
      77161:data<=16'd7926;
      77162:data<=16'd8648;
      77163:data<=16'd7509;
      77164:data<=16'd9248;
      77165:data<=16'd7354;
      77166:data<=-16'd2112;
      77167:data<=-16'd6144;
      77168:data<=-16'd3973;
      77169:data<=-16'd4514;
      77170:data<=-16'd4664;
      77171:data<=-16'd3715;
      77172:data<=-16'd3773;
      77173:data<=-16'd2311;
      77174:data<=-16'd1225;
      77175:data<=-16'd898;
      77176:data<=-16'd86;
      77177:data<=-16'd889;
      77178:data<=16'd193;
      77179:data<=16'd3850;
      77180:data<=16'd4463;
      77181:data<=16'd3962;
      77182:data<=16'd4454;
      77183:data<=16'd3717;
      77184:data<=16'd3218;
      77185:data<=16'd3450;
      77186:data<=16'd4003;
      77187:data<=16'd5324;
      77188:data<=16'd5421;
      77189:data<=16'd4883;
      77190:data<=16'd5060;
      77191:data<=16'd4558;
      77192:data<=16'd4170;
      77193:data<=16'd4114;
      77194:data<=16'd3805;
      77195:data<=16'd4243;
      77196:data<=16'd3976;
      77197:data<=16'd3318;
      77198:data<=16'd4164;
      77199:data<=16'd4676;
      77200:data<=16'd5278;
      77201:data<=16'd5466;
      77202:data<=16'd3568;
      77203:data<=16'd7000;
      77204:data<=16'd15835;
      77205:data<=16'd17807;
      77206:data<=16'd14792;
      77207:data<=16'd14753;
      77208:data<=16'd14189;
      77209:data<=16'd12649;
      77210:data<=16'd12812;
      77211:data<=16'd12792;
      77212:data<=16'd12866;
      77213:data<=16'd12977;
      77214:data<=16'd12193;
      77215:data<=16'd11788;
      77216:data<=16'd10919;
      77217:data<=16'd10006;
      77218:data<=16'd10202;
      77219:data<=16'd9303;
      77220:data<=16'd8425;
      77221:data<=16'd8702;
      77222:data<=16'd7212;
      77223:data<=16'd5160;
      77224:data<=16'd5019;
      77225:data<=16'd5238;
      77226:data<=16'd4734;
      77227:data<=16'd4341;
      77228:data<=16'd4485;
      77229:data<=16'd4115;
      77230:data<=16'd3623;
      77231:data<=16'd3832;
      77232:data<=16'd2826;
      77233:data<=16'd1885;
      77234:data<=16'd2499;
      77235:data<=16'd2021;
      77236:data<=16'd2138;
      77237:data<=16'd3339;
      77238:data<=16'd3341;
      77239:data<=16'd4573;
      77240:data<=16'd2234;
      77241:data<=-16'd6816;
      77242:data<=-16'd10683;
      77243:data<=-16'd8404;
      77244:data<=-16'd8746;
      77245:data<=-16'd9066;
      77246:data<=-16'd8372;
      77247:data<=-16'd8671;
      77248:data<=-16'd7423;
      77249:data<=-16'd5962;
      77250:data<=-16'd5260;
      77251:data<=-16'd4546;
      77252:data<=-16'd5409;
      77253:data<=-16'd5703;
      77254:data<=-16'd4620;
      77255:data<=-16'd4824;
      77256:data<=-16'd5010;
      77257:data<=-16'd4764;
      77258:data<=-16'd4868;
      77259:data<=-16'd4414;
      77260:data<=-16'd4517;
      77261:data<=-16'd4017;
      77262:data<=-16'd2002;
      77263:data<=-16'd2035;
      77264:data<=-16'd2673;
      77265:data<=-16'd2120;
      77266:data<=-16'd2972;
      77267:data<=-16'd1968;
      77268:data<=16'd1465;
      77269:data<=16'd1688;
      77270:data<=16'd776;
      77271:data<=16'd1108;
      77272:data<=16'd1058;
      77273:data<=16'd1823;
      77274:data<=16'd2065;
      77275:data<=16'd2226;
      77276:data<=16'd2949;
      77277:data<=16'd779;
      77278:data<=16'd3516;
      77279:data<=16'd13277;
      77280:data<=16'd14989;
      77281:data<=16'd11223;
      77282:data<=16'd11717;
      77283:data<=16'd11042;
      77284:data<=16'd9922;
      77285:data<=16'd10160;
      77286:data<=16'd9256;
      77287:data<=16'd10690;
      77288:data<=16'd11197;
      77289:data<=16'd8775;
      77290:data<=16'd8690;
      77291:data<=16'd8132;
      77292:data<=16'd7000;
      77293:data<=16'd7336;
      77294:data<=16'd5618;
      77295:data<=16'd4839;
      77296:data<=16'd5700;
      77297:data<=16'd4908;
      77298:data<=16'd5280;
      77299:data<=16'd6067;
      77300:data<=16'd5914;
      77301:data<=16'd6015;
      77302:data<=16'd5004;
      77303:data<=16'd4469;
      77304:data<=16'd4300;
      77305:data<=16'd3391;
      77306:data<=16'd3568;
      77307:data<=16'd2714;
      77308:data<=16'd1895;
      77309:data<=16'd2608;
      77310:data<=16'd1886;
      77311:data<=16'd2218;
      77312:data<=16'd1577;
      77313:data<=-16'd1647;
      77314:data<=-16'd517;
      77315:data<=-16'd2220;
      77316:data<=-16'd11398;
      77317:data<=-16'd14945;
      77318:data<=-16'd13418;
      77319:data<=-16'd13976;
      77320:data<=-16'd13474;
      77321:data<=-16'd12536;
      77322:data<=-16'd12542;
      77323:data<=-16'd12217;
      77324:data<=-16'd12051;
      77325:data<=-16'd11453;
      77326:data<=-16'd11303;
      77327:data<=-16'd11909;
      77328:data<=-16'd11564;
      77329:data<=-16'd10986;
      77330:data<=-16'd10555;
      77331:data<=-16'd9976;
      77332:data<=-16'd9715;
      77333:data<=-16'd9759;
      77334:data<=-16'd9721;
      77335:data<=-16'd8992;
      77336:data<=-16'd9110;
      77337:data<=-16'd10733;
      77338:data<=-16'd11256;
      77339:data<=-16'd10856;
      77340:data<=-16'd10692;
      77341:data<=-16'd10431;
      77342:data<=-16'd10414;
      77343:data<=-16'd10031;
      77344:data<=-16'd9373;
      77345:data<=-16'd9224;
      77346:data<=-16'd9150;
      77347:data<=-16'd8658;
      77348:data<=-16'd8287;
      77349:data<=-16'd9761;
      77350:data<=-16'd10193;
      77351:data<=-16'd8860;
      77352:data<=-16'd11077;
      77353:data<=-16'd8414;
      77354:data<=16'd2497;
      77355:data<=16'd4825;
      77356:data<=16'd2306;
      77357:data<=16'd6247;
      77358:data<=16'd7087;
      77359:data<=16'd5574;
      77360:data<=16'd6466;
      77361:data<=16'd4560;
      77362:data<=16'd3265;
      77363:data<=16'd3190;
      77364:data<=16'd1895;
      77365:data<=16'd2358;
      77366:data<=16'd1858;
      77367:data<=16'd1096;
      77368:data<=16'd2055;
      77369:data<=16'd1128;
      77370:data<=16'd866;
      77371:data<=16'd1372;
      77372:data<=16'd462;
      77373:data<=16'd629;
      77374:data<=-16'd523;
      77375:data<=-16'd2259;
      77376:data<=-16'd1776;
      77377:data<=-16'd2171;
      77378:data<=-16'd2130;
      77379:data<=-16'd1535;
      77380:data<=-16'd2331;
      77381:data<=-16'd2000;
      77382:data<=-16'd1829;
      77383:data<=-16'd2105;
      77384:data<=-16'd1670;
      77385:data<=-16'd2258;
      77386:data<=-16'd2240;
      77387:data<=-16'd3139;
      77388:data<=-16'd4695;
      77389:data<=-16'd2669;
      77390:data<=-16'd4901;
      77391:data<=-16'd13452;
      77392:data<=-16'd16850;
      77393:data<=-16'd15435;
      77394:data<=-16'd14956;
      77395:data<=-16'd14798;
      77396:data<=-16'd14366;
      77397:data<=-16'd13388;
      77398:data<=-16'd13015;
      77399:data<=-16'd13333;
      77400:data<=-16'd13162;
      77401:data<=-16'd14474;
      77402:data<=-16'd16642;
      77403:data<=-16'd16789;
      77404:data<=-16'd15386;
      77405:data<=-16'd14111;
      77406:data<=-16'd13584;
      77407:data<=-16'd13192;
      77408:data<=-16'd13129;
      77409:data<=-16'd12871;
      77410:data<=-16'd11353;
      77411:data<=-16'd11229;
      77412:data<=-16'd12296;
      77413:data<=-16'd11947;
      77414:data<=-16'd11837;
      77415:data<=-16'd11552;
      77416:data<=-16'd10360;
      77417:data<=-16'd9894;
      77418:data<=-16'd9385;
      77419:data<=-16'd9053;
      77420:data<=-16'd8987;
      77421:data<=-16'd8370;
      77422:data<=-16'd7691;
      77423:data<=-16'd6789;
      77424:data<=-16'd7647;
      77425:data<=-16'd8825;
      77426:data<=-16'd7812;
      77427:data<=-16'd8634;
      77428:data<=-16'd5401;
      77429:data<=16'd5095;
      77430:data<=16'd8152;
      77431:data<=16'd4913;
      77432:data<=16'd5724;
      77433:data<=16'd5630;
      77434:data<=16'd4899;
      77435:data<=16'd5962;
      77436:data<=16'd5006;
      77437:data<=16'd4006;
      77438:data<=16'd3563;
      77439:data<=16'd3145;
      77440:data<=16'd4005;
      77441:data<=16'd3817;
      77442:data<=16'd3560;
      77443:data<=16'd3645;
      77444:data<=16'd2696;
      77445:data<=16'd4138;
      77446:data<=16'd6711;
      77447:data<=16'd7488;
      77448:data<=16'd7765;
      77449:data<=16'd6664;
      77450:data<=16'd5383;
      77451:data<=16'd5242;
      77452:data<=16'd4743;
      77453:data<=16'd5006;
      77454:data<=16'd5312;
      77455:data<=16'd5030;
      77456:data<=16'd5770;
      77457:data<=16'd5727;
      77458:data<=16'd5104;
      77459:data<=16'd5388;
      77460:data<=16'd5292;
      77461:data<=16'd5045;
      77462:data<=16'd3838;
      77463:data<=16'd2598;
      77464:data<=16'd4064;
      77465:data<=16'd2399;
      77466:data<=-16'd5379;
      77467:data<=-16'd9988;
      77468:data<=-16'd8625;
      77469:data<=-16'd7727;
      77470:data<=-16'd7776;
      77471:data<=-16'd6887;
      77472:data<=-16'd6713;
      77473:data<=-16'd6601;
      77474:data<=-16'd6156;
      77475:data<=-16'd6716;
      77476:data<=-16'd6605;
      77477:data<=-16'd6253;
      77478:data<=-16'd6711;
      77479:data<=-16'd5388;
      77480:data<=-16'd3996;
      77481:data<=-16'd4393;
      77482:data<=-16'd4105;
      77483:data<=-16'd3727;
      77484:data<=-16'd3482;
      77485:data<=-16'd2801;
      77486:data<=-16'd3148;
      77487:data<=-16'd3683;
      77488:data<=-16'd4032;
      77489:data<=-16'd3955;
      77490:data<=-16'd3535;
      77491:data<=-16'd4937;
      77492:data<=-16'd5230;
      77493:data<=-16'd3714;
      77494:data<=-16'd3935;
      77495:data<=-16'd3344;
      77496:data<=-16'd2795;
      77497:data<=-16'd3325;
      77498:data<=-16'd1613;
      77499:data<=-16'd2275;
      77500:data<=-16'd4220;
      77501:data<=-16'd3131;
      77502:data<=-16'd4267;
      77503:data<=-16'd1013;
      77504:data<=16'd9530;
      77505:data<=16'd12082;
      77506:data<=16'd9179;
      77507:data<=16'd10461;
      77508:data<=16'd10458;
      77509:data<=16'd9338;
      77510:data<=16'd9561;
      77511:data<=16'd8505;
      77512:data<=16'd7603;
      77513:data<=16'd7074;
      77514:data<=16'd6420;
      77515:data<=16'd6748;
      77516:data<=16'd6690;
      77517:data<=16'd6199;
      77518:data<=16'd6270;
      77519:data<=16'd6511;
      77520:data<=16'd6452;
      77521:data<=16'd6111;
      77522:data<=16'd6455;
      77523:data<=16'd6648;
      77524:data<=16'd5953;
      77525:data<=16'd5905;
      77526:data<=16'd5917;
      77527:data<=16'd6075;
      77528:data<=16'd6987;
      77529:data<=16'd6566;
      77530:data<=16'd5937;
      77531:data<=16'd6561;
      77532:data<=16'd6446;
      77533:data<=16'd6018;
      77534:data<=16'd6024;
      77535:data<=16'd6297;
      77536:data<=16'd7661;
      77537:data<=16'd8469;
      77538:data<=16'd8439;
      77539:data<=16'd9515;
      77540:data<=16'd7787;
      77541:data<=16'd502;
      77542:data<=-16'd4790;
      77543:data<=-16'd4026;
      77544:data<=-16'd3432;
      77545:data<=-16'd4159;
      77546:data<=-16'd2898;
      77547:data<=-16'd2494;
      77548:data<=-16'd3454;
      77549:data<=-16'd2303;
      77550:data<=-16'd297;
      77551:data<=16'd584;
      77552:data<=16'd446;
      77553:data<=-16'd12;
      77554:data<=16'd414;
      77555:data<=16'd955;
      77556:data<=16'd943;
      77557:data<=16'd644;
      77558:data<=16'd61;
      77559:data<=16'd170;
      77560:data<=16'd221;
      77561:data<=16'd253;
      77562:data<=16'd1692;
      77563:data<=16'd2190;
      77564:data<=16'd2162;
      77565:data<=16'd3372;
      77566:data<=16'd3052;
      77567:data<=16'd2429;
      77568:data<=16'd2896;
      77569:data<=16'd2378;
      77570:data<=16'd2296;
      77571:data<=16'd2387;
      77572:data<=16'd2262;
      77573:data<=16'd3098;
      77574:data<=16'd2987;
      77575:data<=16'd4373;
      77576:data<=16'd6055;
      77577:data<=16'd3466;
      77578:data<=16'd6498;
      77579:data<=16'd15640;
      77580:data<=16'd16380;
      77581:data<=16'd13177;
      77582:data<=16'd13661;
      77583:data<=16'd12851;
      77584:data<=16'd12122;
      77585:data<=16'd12181;
      77586:data<=16'd10978;
      77587:data<=16'd11843;
      77588:data<=16'd12901;
      77589:data<=16'd12058;
      77590:data<=16'd12122;
      77591:data<=16'd11600;
      77592:data<=16'd10157;
      77593:data<=16'd10032;
      77594:data<=16'd9938;
      77595:data<=16'd9216;
      77596:data<=16'd8734;
      77597:data<=16'd8693;
      77598:data<=16'd8807;
      77599:data<=16'd8900;
      77600:data<=16'd9662;
      77601:data<=16'd9940;
      77602:data<=16'd9177;
      77603:data<=16'd9351;
      77604:data<=16'd9162;
      77605:data<=16'd7932;
      77606:data<=16'd7924;
      77607:data<=16'd7899;
      77608:data<=16'd7283;
      77609:data<=16'd7056;
      77610:data<=16'd5949;
      77611:data<=16'd5406;
      77612:data<=16'd6482;
      77613:data<=16'd7360;
      77614:data<=16'd8290;
      77615:data<=16'd6058;
      77616:data<=-16'd1792;
      77617:data<=-16'd7157;
      77618:data<=-16'd6329;
      77619:data<=-16'd5867;
      77620:data<=-16'd6661;
      77621:data<=-16'd5903;
      77622:data<=-16'd5521;
      77623:data<=-16'd5708;
      77624:data<=-16'd3955;
      77625:data<=-16'd1243;
      77626:data<=-16'd349;
      77627:data<=-16'd940;
      77628:data<=-16'd999;
      77629:data<=-16'd925;
      77630:data<=-16'd1412;
      77631:data<=-16'd1240;
      77632:data<=-16'd984;
      77633:data<=-16'd1512;
      77634:data<=-16'd1483;
      77635:data<=-16'd1516;
      77636:data<=-16'd1982;
      77637:data<=-16'd763;
      77638:data<=16'd825;
      77639:data<=16'd591;
      77640:data<=16'd26;
      77641:data<=-16'd14;
      77642:data<=-16'd38;
      77643:data<=-16'd199;
      77644:data<=-16'd432;
      77645:data<=-16'd631;
      77646:data<=-16'd1052;
      77647:data<=-16'd526;
      77648:data<=16'd293;
      77649:data<=-16'd754;
      77650:data<=16'd6;
      77651:data<=16'd1686;
      77652:data<=-16'd475;
      77653:data<=16'd2328;
      77654:data<=16'd11571;
      77655:data<=16'd13523;
      77656:data<=16'd11145;
      77657:data<=16'd11934;
      77658:data<=16'd10557;
      77659:data<=16'd9135;
      77660:data<=16'd10201;
      77661:data<=16'd9391;
      77662:data<=16'd9124;
      77663:data<=16'd9809;
      77664:data<=16'd8849;
      77665:data<=16'd8804;
      77666:data<=16'd9021;
      77667:data<=16'd8191;
      77668:data<=16'd7310;
      77669:data<=16'd5344;
      77670:data<=16'd3921;
      77671:data<=16'd4247;
      77672:data<=16'd4259;
      77673:data<=16'd3824;
      77674:data<=16'd3482;
      77675:data<=16'd4246;
      77676:data<=16'd5368;
      77677:data<=16'd4464;
      77678:data<=16'd3973;
      77679:data<=16'd4352;
      77680:data<=16'd3116;
      77681:data<=16'd2517;
      77682:data<=16'd2261;
      77683:data<=16'd1111;
      77684:data<=16'd1541;
      77685:data<=16'd1701;
      77686:data<=16'd855;
      77687:data<=16'd1504;
      77688:data<=16'd2223;
      77689:data<=16'd2984;
      77690:data<=16'd1838;
      77691:data<=-16'd5219;
      77692:data<=-16'd11423;
      77693:data<=-16'd11267;
      77694:data<=-16'd10557;
      77695:data<=-16'd11151;
      77696:data<=-16'd10783;
      77697:data<=-16'd10422;
      77698:data<=-16'd10282;
      77699:data<=-16'd9815;
      77700:data<=-16'd8534;
      77701:data<=-16'd6913;
      77702:data<=-16'd7010;
      77703:data<=-16'd7371;
      77704:data<=-16'd6376;
      77705:data<=-16'd6320;
      77706:data<=-16'd6968;
      77707:data<=-16'd6927;
      77708:data<=-16'd6852;
      77709:data<=-16'd6352;
      77710:data<=-16'd6241;
      77711:data<=-16'd7054;
      77712:data<=-16'd6264;
      77713:data<=-16'd4032;
      77714:data<=-16'd2725;
      77715:data<=-16'd2684;
      77716:data<=-16'd3002;
      77717:data<=-16'd2754;
      77718:data<=-16'd2692;
      77719:data<=-16'd2883;
      77720:data<=-16'd2590;
      77721:data<=-16'd3237;
      77722:data<=-16'd3482;
      77723:data<=-16'd2643;
      77724:data<=-16'd3556;
      77725:data<=-16'd3409;
      77726:data<=-16'd2476;
      77727:data<=-16'd4226;
      77728:data<=-16'd553;
      77729:data<=16'd8281;
      77730:data<=16'd9794;
      77731:data<=16'd7480;
      77732:data<=16'd8301;
      77733:data<=16'd8116;
      77734:data<=16'd6951;
      77735:data<=16'd6601;
      77736:data<=16'd6109;
      77737:data<=16'd5545;
      77738:data<=16'd3736;
      77739:data<=16'd2074;
      77740:data<=16'd2124;
      77741:data<=16'd1627;
      77742:data<=16'd1115;
      77743:data<=16'd1263;
      77744:data<=16'd948;
      77745:data<=16'd936;
      77746:data<=16'd597;
      77747:data<=16'd61;
      77748:data<=16'd534;
      77749:data<=-16'd18;
      77750:data<=-16'd1516;
      77751:data<=-16'd1971;
      77752:data<=-16'd2087;
      77753:data<=-16'd2209;
      77754:data<=-16'd2604;
      77755:data<=-16'd3189;
      77756:data<=-16'd2678;
      77757:data<=-16'd2494;
      77758:data<=-16'd3852;
      77759:data<=-16'd5049;
      77760:data<=-16'd5292;
      77761:data<=-16'd4748;
      77762:data<=-16'd5040;
      77763:data<=-16'd6937;
      77764:data<=-16'd7092;
      77765:data<=-16'd7570;
      77766:data<=-16'd13787;
      77767:data<=-16'd19525;
      77768:data<=-16'd18979;
      77769:data<=-16'd18073;
      77770:data<=-16'd18377;
      77771:data<=-16'd17246;
      77772:data<=-16'd16954;
      77773:data<=-16'd16841;
      77774:data<=-16'd15618;
      77775:data<=-16'd15752;
      77776:data<=-16'd16413;
      77777:data<=-16'd16298;
      77778:data<=-16'd16104;
      77779:data<=-16'd15330;
      77780:data<=-16'd14522;
      77781:data<=-16'd14129;
      77782:data<=-16'd13637;
      77783:data<=-16'd13157;
      77784:data<=-16'd12405;
      77785:data<=-16'd11817;
      77786:data<=-16'd11453;
      77787:data<=-16'd11374;
      77788:data<=-16'd12809;
      77789:data<=-16'd13634;
      77790:data<=-16'd12721;
      77791:data<=-16'd12248;
      77792:data<=-16'd11403;
      77793:data<=-16'd10655;
      77794:data<=-16'd10748;
      77795:data<=-16'd9720;
      77796:data<=-16'd9332;
      77797:data<=-16'd9426;
      77798:data<=-16'd8328;
      77799:data<=-16'd8560;
      77800:data<=-16'd8596;
      77801:data<=-16'd8740;
      77802:data<=-16'd10434;
      77803:data<=-16'd5181;
      77804:data<=16'd4984;
      77805:data<=16'd7468;
      77806:data<=16'd5567;
      77807:data<=16'd5870;
      77808:data<=16'd5852;
      77809:data<=16'd5377;
      77810:data<=16'd5366;
      77811:data<=16'd5242;
      77812:data<=16'd4423;
      77813:data<=16'd2578;
      77814:data<=16'd1898;
      77815:data<=16'd2575;
      77816:data<=16'd2475;
      77817:data<=16'd2043;
      77818:data<=16'd1889;
      77819:data<=16'd2090;
      77820:data<=16'd2364;
      77821:data<=16'd1955;
      77822:data<=16'd1721;
      77823:data<=16'd1958;
      77824:data<=16'd2056;
      77825:data<=16'd1580;
      77826:data<=16'd38;
      77827:data<=-16'd563;
      77828:data<=16'd376;
      77829:data<=16'd373;
      77830:data<=16'd115;
      77831:data<=16'd253;
      77832:data<=-16'd196;
      77833:data<=16'd318;
      77834:data<=16'd1092;
      77835:data<=16'd262;
      77836:data<=-16'd82;
      77837:data<=-16'd183;
      77838:data<=-16'd1480;
      77839:data<=-16'd1174;
      77840:data<=-16'd1559;
      77841:data<=-16'd8116;
      77842:data<=-16'd14442;
      77843:data<=-16'd13806;
      77844:data<=-16'd12396;
      77845:data<=-16'd12801;
      77846:data<=-16'd11746;
      77847:data<=-16'd11658;
      77848:data<=-16'd12401;
      77849:data<=-16'd11511;
      77850:data<=-16'd11762;
      77851:data<=-16'd12871;
      77852:data<=-16'd12286;
      77853:data<=-16'd11468;
      77854:data<=-16'd11071;
      77855:data<=-16'd10443;
      77856:data<=-16'd9861;
      77857:data<=-16'd9433;
      77858:data<=-16'd8780;
      77859:data<=-16'd7890;
      77860:data<=-16'd7893;
      77861:data<=-16'd8079;
      77862:data<=-16'd7498;
      77863:data<=-16'd8022;
      77864:data<=-16'd8792;
      77865:data<=-16'd8455;
      77866:data<=-16'd8379;
      77867:data<=-16'd7594;
      77868:data<=-16'd6590;
      77869:data<=-16'd6667;
      77870:data<=-16'd5921;
      77871:data<=-16'd5128;
      77872:data<=-16'd4645;
      77873:data<=-16'd3780;
      77874:data<=-16'd4299;
      77875:data<=-16'd4002;
      77876:data<=-16'd3711;
      77877:data<=-16'd6072;
      77878:data<=-16'd2467;
      77879:data<=16'd7210;
      77880:data<=16'd10378;
      77881:data<=16'd8746;
      77882:data<=16'd9368;
      77883:data<=16'd9700;
      77884:data<=16'd8989;
      77885:data<=16'd9057;
      77886:data<=16'd9529;
      77887:data<=16'd9162;
      77888:data<=16'd7344;
      77889:data<=16'd6297;
      77890:data<=16'd6815;
      77891:data<=16'd7230;
      77892:data<=16'd7881;
      77893:data<=16'd8304;
      77894:data<=16'd7911;
      77895:data<=16'd8155;
      77896:data<=16'd8478;
      77897:data<=16'd8241;
      77898:data<=16'd8432;
      77899:data<=16'd8379;
      77900:data<=16'd7536;
      77901:data<=16'd6661;
      77902:data<=16'd6267;
      77903:data<=16'd6496;
      77904:data<=16'd6616;
      77905:data<=16'd6475;
      77906:data<=16'd6510;
      77907:data<=16'd5890;
      77908:data<=16'd5471;
      77909:data<=16'd6185;
      77910:data<=16'd5814;
      77911:data<=16'd5195;
      77912:data<=16'd5565;
      77913:data<=16'd3977;
      77914:data<=16'd2971;
      77915:data<=16'd3644;
      77916:data<=-16'd1770;
      77917:data<=-16'd9450;
      77918:data<=-16'd9505;
      77919:data<=-16'd7517;
      77920:data<=-16'd8079;
      77921:data<=-16'd7177;
      77922:data<=-16'd6159;
      77923:data<=-16'd6141;
      77924:data<=-16'd5609;
      77925:data<=-16'd5485;
      77926:data<=-16'd5234;
      77927:data<=-16'd4842;
      77928:data<=-16'd4889;
      77929:data<=-16'd4193;
      77930:data<=-16'd3589;
      77931:data<=-16'd3436;
      77932:data<=-16'd3034;
      77933:data<=-16'd3118;
      77934:data<=-16'd2582;
      77935:data<=-16'd1516;
      77936:data<=-16'd2317;
      77937:data<=-16'd3692;
      77938:data<=-16'd3066;
      77939:data<=-16'd1319;
      77940:data<=-16'd1004;
      77941:data<=-16'd1657;
      77942:data<=-16'd910;
      77943:data<=16'd138;
      77944:data<=16'd579;
      77945:data<=16'd1011;
      77946:data<=16'd531;
      77947:data<=16'd1008;
      77948:data<=16'd2085;
      77949:data<=16'd773;
      77950:data<=16'd1579;
      77951:data<=16'd4096;
      77952:data<=16'd2896;
      77953:data<=16'd5924;
      77954:data<=16'd15414;
      77955:data<=16'd18786;
      77956:data<=16'd16202;
      77957:data<=16'd15681;
      77958:data<=16'd15735;
      77959:data<=16'd15047;
      77960:data<=16'd14722;
      77961:data<=16'd13954;
      77962:data<=16'd13467;
      77963:data<=16'd14079;
      77964:data<=16'd14973;
      77965:data<=16'd15183;
      77966:data<=16'd14448;
      77967:data<=16'd13861;
      77968:data<=16'd13659;
      77969:data<=16'd13217;
      77970:data<=16'd12821;
      77971:data<=16'd12196;
      77972:data<=16'd11723;
      77973:data<=16'd12028;
      77974:data<=16'd11717;
      77975:data<=16'd11456;
      77976:data<=16'd12416;
      77977:data<=16'd12599;
      77978:data<=16'd12328;
      77979:data<=16'd12636;
      77980:data<=16'd12358;
      77981:data<=16'd12695;
      77982:data<=16'd13274;
      77983:data<=16'd12295;
      77984:data<=16'd11811;
      77985:data<=16'd11728;
      77986:data<=16'd11044;
      77987:data<=16'd11048;
      77988:data<=16'd10686;
      77989:data<=16'd11221;
      77990:data<=16'd11873;
      77991:data<=16'd5929;
      77992:data<=-16'd1909;
      77993:data<=-16'd2767;
      77994:data<=-16'd1383;
      77995:data<=-16'd1855;
      77996:data<=-16'd1947;
      77997:data<=-16'd1738;
      77998:data<=-16'd1406;
      77999:data<=-16'd1427;
      78000:data<=-16'd1577;
      78001:data<=-16'd446;
      78002:data<=16'd318;
      78003:data<=16'd367;
      78004:data<=16'd763;
      78005:data<=16'd569;
      78006:data<=16'd508;
      78007:data<=16'd640;
      78008:data<=16'd44;
      78009:data<=16'd77;
      78010:data<=16'd552;
      78011:data<=16'd384;
      78012:data<=-16'd124;
      78013:data<=-16'd9;
      78014:data<=16'd1557;
      78015:data<=16'd2053;
      78016:data<=16'd790;
      78017:data<=16'd883;
      78018:data<=16'd939;
      78019:data<=16'd387;
      78020:data<=16'd1336;
      78021:data<=16'd1415;
      78022:data<=16'd946;
      78023:data<=16'd1397;
      78024:data<=16'd405;
      78025:data<=16'd643;
      78026:data<=16'd2030;
      78027:data<=16'd243;
      78028:data<=16'd2575;
      78029:data<=16'd11644;
      78030:data<=16'd15091;
      78031:data<=16'd12296;
      78032:data<=16'd11982;
      78033:data<=16'd12248;
      78034:data<=16'd11126;
      78035:data<=16'd11180;
      78036:data<=16'd10857;
      78037:data<=16'd9747;
      78038:data<=16'd9996;
      78039:data<=16'd10942;
      78040:data<=16'd11347;
      78041:data<=16'd10840;
      78042:data<=16'd9796;
      78043:data<=16'd8984;
      78044:data<=16'd8249;
      78045:data<=16'd8058;
      78046:data<=16'd7993;
      78047:data<=16'd6839;
      78048:data<=16'd6226;
      78049:data<=16'd6360;
      78050:data<=16'd6149;
      78051:data<=16'd6877;
      78052:data<=16'd7391;
      78053:data<=16'd6959;
      78054:data<=16'd7409;
      78055:data<=16'd7175;
      78056:data<=16'd5985;
      78057:data<=16'd5603;
      78058:data<=16'd5195;
      78059:data<=16'd5121;
      78060:data<=16'd4858;
      78061:data<=16'd3861;
      78062:data<=16'd4241;
      78063:data<=16'd4272;
      78064:data<=16'd4179;
      78065:data<=16'd5292;
      78066:data<=16'd643;
      78067:data<=-16'd7978;
      78068:data<=-16'd9952;
      78069:data<=-16'd7943;
      78070:data<=-16'd7319;
      78071:data<=-16'd6511;
      78072:data<=-16'd6194;
      78073:data<=-16'd6185;
      78074:data<=-16'd5764;
      78075:data<=-16'd6052;
      78076:data<=-16'd5627;
      78077:data<=-16'd4538;
      78078:data<=-16'd4410;
      78079:data<=-16'd4326;
      78080:data<=-16'd4126;
      78081:data<=-16'd4266;
      78082:data<=-16'd4373;
      78083:data<=-16'd4313;
      78084:data<=-16'd4037;
      78085:data<=-16'd4126;
      78086:data<=-16'd4585;
      78087:data<=-16'd4690;
      78088:data<=-16'd4011;
      78089:data<=-16'd2499;
      78090:data<=-16'd2293;
      78091:data<=-16'd3706;
      78092:data<=-16'd3715;
      78093:data<=-16'd3048;
      78094:data<=-16'd3095;
      78095:data<=-16'd2972;
      78096:data<=-16'd3500;
      78097:data<=-16'd3445;
      78098:data<=-16'd2582;
      78099:data<=-16'd3651;
      78100:data<=-16'd3560;
      78101:data<=-16'd1789;
      78102:data<=-16'd2432;
      78103:data<=16'd364;
      78104:data<=16'd8627;
      78105:data<=16'd12032;
      78106:data<=16'd10325;
      78107:data<=16'd9914;
      78108:data<=16'd9056;
      78109:data<=16'd7777;
      78110:data<=16'd8117;
      78111:data<=16'd7696;
      78112:data<=16'd6983;
      78113:data<=16'd7597;
      78114:data<=16'd7374;
      78115:data<=16'd6003;
      78116:data<=16'd4951;
      78117:data<=16'd4176;
      78118:data<=16'd3516;
      78119:data<=16'd2930;
      78120:data<=16'd2588;
      78121:data<=16'd2320;
      78122:data<=16'd1830;
      78123:data<=16'd2030;
      78124:data<=16'd2300;
      78125:data<=16'd1723;
      78126:data<=16'd1632;
      78127:data<=16'd1434;
      78128:data<=16'd506;
      78129:data<=16'd361;
      78130:data<=16'd560;
      78131:data<=16'd635;
      78132:data<=16'd177;
      78133:data<=-16'd1154;
      78134:data<=-16'd1049;
      78135:data<=-16'd737;
      78136:data<=-16'd1409;
      78137:data<=-16'd537;
      78138:data<=-16'd1759;
      78139:data<=-16'd4528;
      78140:data<=-16'd3641;
      78141:data<=-16'd7520;
      78142:data<=-16'd16921;
      78143:data<=-16'd18692;
      78144:data<=-16'd16286;
      78145:data<=-16'd16803;
      78146:data<=-16'd16149;
      78147:data<=-16'd15446;
      78148:data<=-16'd15544;
      78149:data<=-16'd14225;
      78150:data<=-16'd13876;
      78151:data<=-16'd14595;
      78152:data<=-16'd15443;
      78153:data<=-16'd16017;
      78154:data<=-16'd14766;
      78155:data<=-16'd13922;
      78156:data<=-16'd13834;
      78157:data<=-16'd13042;
      78158:data<=-16'd13138;
      78159:data<=-16'd12134;
      78160:data<=-16'd9823;
      78161:data<=-16'd9668;
      78162:data<=-16'd9818;
      78163:data<=-16'd9718;
      78164:data<=-16'd10813;
      78165:data<=-16'd11398;
      78166:data<=-16'd11717;
      78167:data<=-16'd11756;
      78168:data<=-16'd11033;
      78169:data<=-16'd10800;
      78170:data<=-16'd10160;
      78171:data<=-16'd9564;
      78172:data<=-16'd9549;
      78173:data<=-16'd8778;
      78174:data<=-16'd8889;
      78175:data<=-16'd8960;
      78176:data<=-16'd8730;
      78177:data<=-16'd10830;
      78178:data<=-16'd8126;
      78179:data<=16'd1105;
      78180:data<=16'd4811;
      78181:data<=16'd3339;
      78182:data<=16'd3589;
      78183:data<=16'd3265;
      78184:data<=16'd2922;
      78185:data<=16'd3381;
      78186:data<=16'd2452;
      78187:data<=16'd2484;
      78188:data<=16'd2787;
      78189:data<=16'd1124;
      78190:data<=16'd488;
      78191:data<=16'd608;
      78192:data<=-16'd229;
      78193:data<=-16'd315;
      78194:data<=-16'd259;
      78195:data<=-16'd690;
      78196:data<=-16'd420;
      78197:data<=-16'd220;
      78198:data<=-16'd443;
      78199:data<=-16'd347;
      78200:data<=-16'd45;
      78201:data<=-16'd182;
      78202:data<=-16'd1303;
      78203:data<=-16'd2341;
      78204:data<=-16'd2828;
      78205:data<=-16'd3400;
      78206:data<=-16'd3033;
      78207:data<=-16'd2857;
      78208:data<=-16'd3765;
      78209:data<=-16'd3115;
      78210:data<=-16'd2786;
      78211:data<=-16'd3566;
      78212:data<=-16'd2056;
      78213:data<=-16'd2272;
      78214:data<=-16'd4325;
      78215:data<=-16'd3221;
      78216:data<=-16'd6895;
      78217:data<=-16'd16126;
      78218:data<=-16'd17969;
      78219:data<=-16'd15235;
      78220:data<=-16'd15481;
      78221:data<=-16'd14853;
      78222:data<=-16'd13782;
      78223:data<=-16'd14090;
      78224:data<=-16'd13139;
      78225:data<=-16'd11967;
      78226:data<=-16'd12358;
      78227:data<=-16'd13584;
      78228:data<=-16'd13841;
      78229:data<=-16'd12625;
      78230:data<=-16'd12113;
      78231:data<=-16'd11494;
      78232:data<=-16'd10107;
      78233:data<=-16'd10293;
      78234:data<=-16'd10134;
      78235:data<=-16'd9083;
      78236:data<=-16'd9471;
      78237:data<=-16'd9012;
      78238:data<=-16'd8056;
      78239:data<=-16'd8866;
      78240:data<=-16'd9165;
      78241:data<=-16'd8934;
      78242:data<=-16'd8916;
      78243:data<=-16'd8120;
      78244:data<=-16'd7598;
      78245:data<=-16'd7101;
      78246:data<=-16'd6384;
      78247:data<=-16'd6229;
      78248:data<=-16'd5612;
      78249:data<=-16'd4675;
      78250:data<=-16'd3177;
      78251:data<=-16'd2496;
      78252:data<=-16'd5040;
      78253:data<=-16'd3169;
      78254:data<=16'd5941;
      78255:data<=16'd10451;
      78256:data<=16'd9244;
      78257:data<=16'd9276;
      78258:data<=16'd8824;
      78259:data<=16'd8276;
      78260:data<=16'd8789;
      78261:data<=16'd8056;
      78262:data<=16'd8011;
      78263:data<=16'd8363;
      78264:data<=16'd7000;
      78265:data<=16'd6234;
      78266:data<=16'd5871;
      78267:data<=16'd5156;
      78268:data<=16'd5350;
      78269:data<=16'd5197;
      78270:data<=16'd4723;
      78271:data<=16'd4875;
      78272:data<=16'd4852;
      78273:data<=16'd4808;
      78274:data<=16'd4786;
      78275:data<=16'd5092;
      78276:data<=16'd5201;
      78277:data<=16'd3494;
      78278:data<=16'd2676;
      78279:data<=16'd3800;
      78280:data<=16'd3730;
      78281:data<=16'd3662;
      78282:data<=16'd3923;
      78283:data<=16'd3127;
      78284:data<=16'd3660;
      78285:data<=16'd3892;
      78286:data<=16'd2641;
      78287:data<=16'd3535;
      78288:data<=16'd3603;
      78289:data<=16'd1821;
      78290:data<=16'd2130;
      78291:data<=-16'd1636;
      78292:data<=-16'd10648;
      78293:data<=-16'd13841;
      78294:data<=-16'd12228;
      78295:data<=-16'd12569;
      78296:data<=-16'd12140;
      78297:data<=-16'd10768;
      78298:data<=-16'd10610;
      78299:data<=-16'd9894;
      78300:data<=-16'd9047;
      78301:data<=-16'd9236;
      78302:data<=-16'd9952;
      78303:data<=-16'd10287;
      78304:data<=-16'd9133;
      78305:data<=-16'd8223;
      78306:data<=-16'd8322;
      78307:data<=-16'd7357;
      78308:data<=-16'd6234;
      78309:data<=-16'd5601;
      78310:data<=-16'd4980;
      78311:data<=-16'd5257;
      78312:data<=-16'd4824;
      78313:data<=-16'd3767;
      78314:data<=-16'd4634;
      78315:data<=-16'd6028;
      78316:data<=-16'd6454;
      78317:data<=-16'd5797;
      78318:data<=-16'd4464;
      78319:data<=-16'd4134;
      78320:data<=-16'd3688;
      78321:data<=-16'd2893;
      78322:data<=-16'd2955;
      78323:data<=-16'd2372;
      78324:data<=-16'd2259;
      78325:data<=-16'd2370;
      78326:data<=-16'd1351;
      78327:data<=-16'd2068;
      78328:data<=16'd766;
      78329:data<=16'd9993;
      78330:data<=16'd14170;
      78331:data<=16'd12900;
      78332:data<=16'd13135;
      78333:data<=16'd12565;
      78334:data<=16'd12446;
      78335:data<=16'd13059;
      78336:data<=16'd11449;
      78337:data<=16'd11709;
      78338:data<=16'd13403;
      78339:data<=16'd13665;
      78340:data<=16'd15048;
      78341:data<=16'd15470;
      78342:data<=16'd14119;
      78343:data<=16'd13940;
      78344:data<=16'd13256;
      78345:data<=16'd12472;
      78346:data<=16'd12819;
      78347:data<=16'd12290;
      78348:data<=16'd11835;
      78349:data<=16'd11536;
      78350:data<=16'd10442;
      78351:data<=16'd10953;
      78352:data<=16'd12684;
      78353:data<=16'd13443;
      78354:data<=16'd13520;
      78355:data<=16'd13029;
      78356:data<=16'd12678;
      78357:data<=16'd12633;
      78358:data<=16'd11781;
      78359:data<=16'd11271;
      78360:data<=16'd11126;
      78361:data<=16'd10501;
      78362:data<=16'd10522;
      78363:data<=16'd9688;
      78364:data<=16'd9470;
      78365:data<=16'd12366;
      78366:data<=16'd9195;
      78367:data<=-16'd974;
      78368:data<=-16'd4088;
      78369:data<=-16'd1877;
      78370:data<=-16'd2491;
      78371:data<=-16'd1983;
      78372:data<=-16'd1209;
      78373:data<=-16'd1936;
      78374:data<=-16'd1392;
      78375:data<=-16'd1727;
      78376:data<=-16'd1260;
      78377:data<=16'd1287;
      78378:data<=16'd1268;
      78379:data<=16'd754;
      78380:data<=16'd1583;
      78381:data<=16'd1513;
      78382:data<=16'd1269;
      78383:data<=16'd111;
      78384:data<=-16'd743;
      78385:data<=16'd174;
      78386:data<=16'd109;
      78387:data<=16'd3;
      78388:data<=16'd121;
      78389:data<=-16'd14;
      78390:data<=16'd1855;
      78391:data<=16'd2364;
      78392:data<=16'd960;
      78393:data<=16'd1447;
      78394:data<=16'd1691;
      78395:data<=16'd1718;
      78396:data<=16'd2053;
      78397:data<=16'd1331;
      78398:data<=16'd1877;
      78399:data<=16'd2003;
      78400:data<=16'd1448;
      78401:data<=16'd2690;
      78402:data<=16'd2467;
      78403:data<=16'd4978;
      78404:data<=16'd13329;
      78405:data<=16'd17352;
      78406:data<=16'd16076;
      78407:data<=16'd15403;
      78408:data<=16'd14777;
      78409:data<=16'd14600;
      78410:data<=16'd13937;
      78411:data<=16'd12593;
      78412:data<=16'd12778;
      78413:data<=16'd12214;
      78414:data<=16'd11937;
      78415:data<=16'd13787;
      78416:data<=16'd13383;
      78417:data<=16'd11593;
      78418:data<=16'd11562;
      78419:data<=16'd11063;
      78420:data<=16'd10158;
      78421:data<=16'd9914;
      78422:data<=16'd9309;
      78423:data<=16'd9154;
      78424:data<=16'd8995;
      78425:data<=16'd7595;
      78426:data<=16'd8079;
      78427:data<=16'd11121;
      78428:data<=16'd12275;
      78429:data<=16'd11699;
      78430:data<=16'd11796;
      78431:data<=16'd11320;
      78432:data<=16'd10431;
      78433:data<=16'd10046;
      78434:data<=16'd9488;
      78435:data<=16'd8570;
      78436:data<=16'd7724;
      78437:data<=16'd7652;
      78438:data<=16'd6784;
      78439:data<=16'd6357;
      78440:data<=16'd9045;
      78441:data<=16'd5803;
      78442:data<=-16'd4549;
      78443:data<=-16'd7333;
      78444:data<=-16'd5060;
      78445:data<=-16'd6172;
      78446:data<=-16'd5624;
      78447:data<=-16'd4942;
      78448:data<=-16'd5612;
      78449:data<=-16'd4378;
      78450:data<=-16'd4989;
      78451:data<=-16'd5745;
      78452:data<=-16'd3845;
      78453:data<=-16'd3442;
      78454:data<=-16'd3588;
      78455:data<=-16'd3163;
      78456:data<=-16'd3162;
      78457:data<=-16'd2764;
      78458:data<=-16'd2992;
      78459:data<=-16'd3078;
      78460:data<=-16'd2998;
      78461:data<=-16'd3315;
      78462:data<=-16'd2408;
      78463:data<=-16'd2851;
      78464:data<=-16'd3510;
      78465:data<=-16'd1609;
      78466:data<=-16'd1707;
      78467:data<=-16'd2393;
      78468:data<=-16'd1500;
      78469:data<=-16'd2217;
      78470:data<=-16'd2282;
      78471:data<=-16'd2617;
      78472:data<=-16'd4379;
      78473:data<=-16'd3785;
      78474:data<=-16'd3917;
      78475:data<=-16'd4563;
      78476:data<=-16'd3424;
      78477:data<=-16'd4306;
      78478:data<=-16'd1513;
      78479:data<=16'd7321;
      78480:data<=16'd11476;
      78481:data<=16'd10560;
      78482:data<=16'd9888;
      78483:data<=16'd9092;
      78484:data<=16'd8719;
      78485:data<=16'd8202;
      78486:data<=16'd7235;
      78487:data<=16'd7033;
      78488:data<=16'd6549;
      78489:data<=16'd6487;
      78490:data<=16'd7771;
      78491:data<=16'd7984;
      78492:data<=16'd6669;
      78493:data<=16'd5891;
      78494:data<=16'd5633;
      78495:data<=16'd5048;
      78496:data<=16'd4828;
      78497:data<=16'd4575;
      78498:data<=16'd3776;
      78499:data<=16'd3559;
      78500:data<=16'd3228;
      78501:data<=16'd2693;
      78502:data<=16'd3419;
      78503:data<=16'd4322;
      78504:data<=16'd4708;
      78505:data<=16'd4582;
      78506:data<=16'd3802;
      78507:data<=16'd3465;
      78508:data<=16'd3018;
      78509:data<=16'd2643;
      78510:data<=16'd2444;
      78511:data<=16'd1231;
      78512:data<=16'd1263;
      78513:data<=16'd1236;
      78514:data<=16'd632;
      78515:data<=16'd3573;
      78516:data<=16'd1642;
      78517:data<=-16'd7903;
      78518:data<=-16'd10812;
      78519:data<=-16'd8828;
      78520:data<=-16'd9746;
      78521:data<=-16'd9232;
      78522:data<=-16'd8719;
      78523:data<=-16'd9259;
      78524:data<=-16'd8270;
      78525:data<=-16'd8407;
      78526:data<=-16'd8593;
      78527:data<=-16'd8147;
      78528:data<=-16'd8693;
      78529:data<=-16'd8188;
      78530:data<=-16'd7876;
      78531:data<=-16'd8158;
      78532:data<=-16'd7454;
      78533:data<=-16'd7562;
      78534:data<=-16'd7371;
      78535:data<=-16'd6992;
      78536:data<=-16'd7928;
      78537:data<=-16'd7232;
      78538:data<=-16'd6258;
      78539:data<=-16'd7453;
      78540:data<=-16'd8727;
      78541:data<=-16'd9700;
      78542:data<=-16'd9823;
      78543:data<=-16'd9273;
      78544:data<=-16'd9498;
      78545:data<=-16'd9359;
      78546:data<=-16'd9101;
      78547:data<=-16'd8669;
      78548:data<=-16'd7712;
      78549:data<=-16'd8237;
      78550:data<=-16'd7981;
      78551:data<=-16'd6763;
      78552:data<=-16'd8681;
      78553:data<=-16'd8181;
      78554:data<=-16'd995;
      78555:data<=16'd4228;
      78556:data<=16'd3771;
      78557:data<=16'd2986;
      78558:data<=16'd3283;
      78559:data<=16'd3101;
      78560:data<=16'd2108;
      78561:data<=16'd506;
      78562:data<=16'd218;
      78563:data<=16'd1148;
      78564:data<=16'd0;
      78565:data<=-16'd2171;
      78566:data<=-16'd2736;
      78567:data<=-16'd3043;
      78568:data<=-16'd3344;
      78569:data<=-16'd3253;
      78570:data<=-16'd3519;
      78571:data<=-16'd3435;
      78572:data<=-16'd3092;
      78573:data<=-16'd2940;
      78574:data<=-16'd3036;
      78575:data<=-16'd3306;
      78576:data<=-16'd2522;
      78577:data<=-16'd2875;
      78578:data<=-16'd5265;
      78579:data<=-16'd5532;
      78580:data<=-16'd4780;
      78581:data<=-16'd4701;
      78582:data<=-16'd3852;
      78583:data<=-16'd4172;
      78584:data<=-16'd4259;
      78585:data<=-16'd3488;
      78586:data<=-16'd4619;
      78587:data<=-16'd4196;
      78588:data<=-16'd3330;
      78589:data<=-16'd4773;
      78590:data<=-16'd4608;
      78591:data<=-16'd8363;
      78592:data<=-16'd17293;
      78593:data<=-16'd19772;
      78594:data<=-16'd17993;
      78595:data<=-16'd17979;
      78596:data<=-16'd16513;
      78597:data<=-16'd15356;
      78598:data<=-16'd15244;
      78599:data<=-16'd14437;
      78600:data<=-16'd14569;
      78601:data<=-16'd13984;
      78602:data<=-16'd13295;
      78603:data<=-16'd14737;
      78604:data<=-16'd14499;
      78605:data<=-16'd12234;
      78606:data<=-16'd11006;
      78607:data<=-16'd10196;
      78608:data<=-16'd9539;
      78609:data<=-16'd9226;
      78610:data<=-16'd8690;
      78611:data<=-16'd8197;
      78612:data<=-16'd7720;
      78613:data<=-16'd7218;
      78614:data<=-16'd7292;
      78615:data<=-16'd8205;
      78616:data<=-16'd8687;
      78617:data<=-16'd8173;
      78618:data<=-16'd8504;
      78619:data<=-16'd8718;
      78620:data<=-16'd7279;
      78621:data<=-16'd6931;
      78622:data<=-16'd7286;
      78623:data<=-16'd6393;
      78624:data<=-16'd6379;
      78625:data<=-16'd5981;
      78626:data<=-16'd4502;
      78627:data<=-16'd6078;
      78628:data<=-16'd6241;
      78629:data<=16'd901;
      78630:data<=16'd7148;
      78631:data<=16'd6655;
      78632:data<=16'd5480;
      78633:data<=16'd5946;
      78634:data<=16'd5870;
      78635:data<=16'd5830;
      78636:data<=16'd5839;
      78637:data<=16'd5698;
      78638:data<=16'd5764;
      78639:data<=16'd5059;
      78640:data<=16'd3806;
      78641:data<=16'd2899;
      78642:data<=16'd2208;
      78643:data<=16'd1997;
      78644:data<=16'd2296;
      78645:data<=16'd2578;
      78646:data<=16'd2114;
      78647:data<=16'd1489;
      78648:data<=16'd2120;
      78649:data<=16'd1768;
      78650:data<=-16'd205;
      78651:data<=-16'd384;
      78652:data<=-16'd529;
      78653:data<=-16'd2014;
      78654:data<=-16'd1619;
      78655:data<=-16'd966;
      78656:data<=-16'd1277;
      78657:data<=-16'd955;
      78658:data<=-16'd1292;
      78659:data<=-16'd1102;
      78660:data<=-16'd202;
      78661:data<=-16'd902;
      78662:data<=-16'd952;
      78663:data<=-16'd914;
      78664:data<=-16'd1545;
      78665:data<=-16'd569;
      78666:data<=-16'd4454;
      78667:data<=-16'd13671;
      78668:data<=-16'd16565;
      78669:data<=-16'd14348;
      78670:data<=-16'd13825;
      78671:data<=-16'd12942;
      78672:data<=-16'd11947;
      78673:data<=-16'd11790;
      78674:data<=-16'd11276;
      78675:data<=-16'd11051;
      78676:data<=-16'd10317;
      78677:data<=-16'd9832;
      78678:data<=-16'd10658;
      78679:data<=-16'd10314;
      78680:data<=-16'd9389;
      78681:data<=-16'd9092;
      78682:data<=-16'd8299;
      78683:data<=-16'd7726;
      78684:data<=-16'd7051;
      78685:data<=-16'd6181;
      78686:data<=-16'd6281;
      78687:data<=-16'd5987;
      78688:data<=-16'd5348;
      78689:data<=-16'd5354;
      78690:data<=-16'd5322;
      78691:data<=-16'd5621;
      78692:data<=-16'd5847;
      78693:data<=-16'd5815;
      78694:data<=-16'd5379;
      78695:data<=-16'd2974;
      78696:data<=-16'd1516;
      78697:data<=-16'd2294;
      78698:data<=-16'd1651;
      78699:data<=-16'd1290;
      78700:data<=-16'd1337;
      78701:data<=16'd352;
      78702:data<=-16'd629;
      78703:data<=-16'd855;
      78704:data<=16'd6354;
      78705:data<=16'd12373;
      78706:data<=16'd11659;
      78707:data<=16'd10792;
      78708:data<=16'd11203;
      78709:data<=16'd10977;
      78710:data<=16'd10850;
      78711:data<=16'd10566;
      78712:data<=16'd10399;
      78713:data<=16'd10492;
      78714:data<=16'd9741;
      78715:data<=16'd8664;
      78716:data<=16'd7879;
      78717:data<=16'd7053;
      78718:data<=16'd6721;
      78719:data<=16'd6934;
      78720:data<=16'd6877;
      78721:data<=16'd6496;
      78722:data<=16'd6199;
      78723:data<=16'd6229;
      78724:data<=16'd6369;
      78725:data<=16'd6391;
      78726:data<=16'd6557;
      78727:data<=16'd6399;
      78728:data<=16'd6056;
      78729:data<=16'd6378;
      78730:data<=16'd6416;
      78731:data<=16'd6328;
      78732:data<=16'd6639;
      78733:data<=16'd6005;
      78734:data<=16'd5930;
      78735:data<=16'd6504;
      78736:data<=16'd5697;
      78737:data<=16'd5882;
      78738:data<=16'd5298;
      78739:data<=16'd3086;
      78740:data<=16'd4884;
      78741:data<=16'd3356;
      78742:data<=-16'd6011;
      78743:data<=-16'd9095;
      78744:data<=-16'd6291;
      78745:data<=-16'd6940;
      78746:data<=-16'd6351;
      78747:data<=-16'd4954;
      78748:data<=-16'd5850;
      78749:data<=-16'd5292;
      78750:data<=-16'd4798;
      78751:data<=-16'd4875;
      78752:data<=-16'd3391;
      78753:data<=-16'd2070;
      78754:data<=-16'd713;
      78755:data<=16'd224;
      78756:data<=16'd32;
      78757:data<=16'd259;
      78758:data<=16'd27;
      78759:data<=16'd329;
      78760:data<=16'd1424;
      78761:data<=16'd572;
      78762:data<=16'd337;
      78763:data<=16'd1377;
      78764:data<=16'd1001;
      78765:data<=16'd1688;
      78766:data<=16'd3577;
      78767:data<=16'd3929;
      78768:data<=16'd3485;
      78769:data<=16'd3269;
      78770:data<=16'd3624;
      78771:data<=16'd3839;
      78772:data<=16'd3563;
      78773:data<=16'd3721;
      78774:data<=16'd3378;
      78775:data<=16'd3380;
      78776:data<=16'd4329;
      78777:data<=16'd3845;
      78778:data<=16'd5768;
      78779:data<=16'd13341;
      78780:data<=16'd19237;
      78781:data<=16'd19071;
      78782:data<=16'd17414;
      78783:data<=16'd17773;
      78784:data<=16'd18832;
      78785:data<=16'd18201;
      78786:data<=16'd16812;
      78787:data<=16'd16824;
      78788:data<=16'd17007;
      78789:data<=16'd16060;
      78790:data<=16'd15837;
      78791:data<=16'd16697;
      78792:data<=16'd16351;
      78793:data<=16'd15402;
      78794:data<=16'd15409;
      78795:data<=16'd14768;
      78796:data<=16'd13471;
      78797:data<=16'd13019;
      78798:data<=16'd12618;
      78799:data<=16'd12037;
      78800:data<=16'd11588;
      78801:data<=16'd10937;
      78802:data<=16'd10983;
      78803:data<=16'd12043;
      78804:data<=16'd12392;
      78805:data<=16'd11326;
      78806:data<=16'd10830;
      78807:data<=16'd10936;
      78808:data<=16'd9800;
      78809:data<=16'd9359;
      78810:data<=16'd9404;
      78811:data<=16'd7934;
      78812:data<=16'd8135;
      78813:data<=16'd8185;
      78814:data<=16'd6485;
      78815:data<=16'd8464;
      78816:data<=16'd7024;
      78817:data<=-16'd2387;
      78818:data<=-16'd5923;
      78819:data<=-16'd3507;
      78820:data<=-16'd4425;
      78821:data<=-16'd4475;
      78822:data<=-16'd3242;
      78823:data<=-16'd4087;
      78824:data<=-16'd4276;
      78825:data<=-16'd4077;
      78826:data<=-16'd4173;
      78827:data<=-16'd3704;
      78828:data<=-16'd3680;
      78829:data<=-16'd3539;
      78830:data<=-16'd2948;
      78831:data<=-16'd2453;
      78832:data<=-16'd2385;
      78833:data<=-16'd3016;
      78834:data<=-16'd2541;
      78835:data<=-16'd1518;
      78836:data<=-16'd2167;
      78837:data<=-16'd2507;
      78838:data<=-16'd1859;
      78839:data<=-16'd1838;
      78840:data<=-16'd1456;
      78841:data<=-16'd100;
      78842:data<=16'd590;
      78843:data<=-16'd287;
      78844:data<=-16'd652;
      78845:data<=16'd525;
      78846:data<=16'd488;
      78847:data<=-16'd388;
      78848:data<=-16'd70;
      78849:data<=-16'd326;
      78850:data<=-16'd434;
      78851:data<=16'd581;
      78852:data<=-16'd325;
      78853:data<=16'd329;
      78854:data<=16'd7891;
      78855:data<=16'd15148;
      78856:data<=16'd15186;
      78857:data<=16'd13198;
      78858:data<=16'd12566;
      78859:data<=16'd11782;
      78860:data<=16'd11749;
      78861:data<=16'd11456;
      78862:data<=16'd10323;
      78863:data<=16'd10326;
      78864:data<=16'd9843;
      78865:data<=16'd9230;
      78866:data<=16'd10390;
      78867:data<=16'd10234;
      78868:data<=16'd9039;
      78869:data<=16'd9204;
      78870:data<=16'd8696;
      78871:data<=16'd7618;
      78872:data<=16'd7642;
      78873:data<=16'd8156;
      78874:data<=16'd8216;
      78875:data<=16'd7512;
      78876:data<=16'd6825;
      78877:data<=16'd6084;
      78878:data<=16'd6164;
      78879:data<=16'd7926;
      78880:data<=16'd7856;
      78881:data<=16'd6502;
      78882:data<=16'd6611;
      78883:data<=16'd5826;
      78884:data<=16'd5456;
      78885:data<=16'd5676;
      78886:data<=16'd4184;
      78887:data<=16'd4601;
      78888:data<=16'd4646;
      78889:data<=16'd2714;
      78890:data<=16'd4367;
      78891:data<=16'd2170;
      78892:data<=-16'd7072;
      78893:data<=-16'd10308;
      78894:data<=-16'd8298;
      78895:data<=-16'd8757;
      78896:data<=-16'd8925;
      78897:data<=-16'd8325;
      78898:data<=-16'd8345;
      78899:data<=-16'd8140;
      78900:data<=-16'd8282;
      78901:data<=-16'd8452;
      78902:data<=-16'd8119;
      78903:data<=-16'd7081;
      78904:data<=-16'd5777;
      78905:data<=-16'd5668;
      78906:data<=-16'd5723;
      78907:data<=-16'd5184;
      78908:data<=-16'd5140;
      78909:data<=-16'd4937;
      78910:data<=-16'd4567;
      78911:data<=-16'd4918;
      78912:data<=-16'd5084;
      78913:data<=-16'd4667;
      78914:data<=-16'd4622;
      78915:data<=-16'd4566;
      78916:data<=-16'd3585;
      78917:data<=-16'd3321;
      78918:data<=-16'd4783;
      78919:data<=-16'd5676;
      78920:data<=-16'd5241;
      78921:data<=-16'd4952;
      78922:data<=-16'd5022;
      78923:data<=-16'd4717;
      78924:data<=-16'd4554;
      78925:data<=-16'd5147;
      78926:data<=-16'd4655;
      78927:data<=-16'd4071;
      78928:data<=-16'd4402;
      78929:data<=16'd828;
      78930:data<=16'd8881;
      78931:data<=16'd9244;
      78932:data<=16'd7089;
      78933:data<=16'd7926;
      78934:data<=16'd7300;
      78935:data<=16'd6684;
      78936:data<=16'd6652;
      78937:data<=16'd5670;
      78938:data<=16'd5909;
      78939:data<=16'd5473;
      78940:data<=16'd3929;
      78941:data<=16'd2793;
      78942:data<=16'd1022;
      78943:data<=16'd869;
      78944:data<=16'd1434;
      78945:data<=16'd478;
      78946:data<=16'd593;
      78947:data<=16'd373;
      78948:data<=-16'd488;
      78949:data<=16'd39;
      78950:data<=-16'd349;
      78951:data<=-16'd649;
      78952:data<=-16'd291;
      78953:data<=-16'd1560;
      78954:data<=-16'd2796;
      78955:data<=-16'd3554;
      78956:data<=-16'd3500;
      78957:data<=-16'd2608;
      78958:data<=-16'd3259;
      78959:data<=-16'd3274;
      78960:data<=-16'd2875;
      78961:data<=-16'd3325;
      78962:data<=-16'd1245;
      78963:data<=-16'd716;
      78964:data<=-16'd2276;
      78965:data<=-16'd773;
      78966:data<=-16'd4921;
      78967:data<=-16'd15493;
      78968:data<=-16'd18616;
      78969:data<=-16'd16098;
      78970:data<=-16'd15578;
      78971:data<=-16'd15104;
      78972:data<=-16'd14587;
      78973:data<=-16'd14552;
      78974:data<=-16'd13712;
      78975:data<=-16'd13227;
      78976:data<=-16'd13126;
      78977:data<=-16'd12393;
      78978:data<=-16'd12548;
      78979:data<=-16'd13808;
      78980:data<=-16'd13667;
      78981:data<=-16'd12619;
      78982:data<=-16'd12463;
      78983:data<=-16'd12019;
      78984:data<=-16'd11288;
      78985:data<=-16'd10778;
      78986:data<=-16'd9973;
      78987:data<=-16'd10058;
      78988:data<=-16'd10052;
      78989:data<=-16'd8734;
      78990:data<=-16'd8866;
      78991:data<=-16'd10414;
      78992:data<=-16'd10583;
      78993:data<=-16'd9737;
      78994:data<=-16'd9535;
      78995:data<=-16'd9535;
      78996:data<=-16'd8943;
      78997:data<=-16'd8987;
      78998:data<=-16'd8863;
      78999:data<=-16'd7733;
      79000:data<=-16'd7937;
      79001:data<=-16'd7335;
      79002:data<=-16'd6296;
      79003:data<=-16'd8222;
      79004:data<=-16'd4434;
      79005:data<=16'd4993;
      79006:data<=16'd5712;
      79007:data<=16'd1692;
      79008:data<=16'd2015;
      79009:data<=16'd2355;
      79010:data<=16'd2197;
      79011:data<=16'd2432;
      79012:data<=16'd1841;
      79013:data<=16'd2215;
      79014:data<=16'd2229;
      79015:data<=16'd1397;
      79016:data<=16'd749;
      79017:data<=-16'd572;
      79018:data<=-16'd698;
      79019:data<=-16'd300;
      79020:data<=-16'd996;
      79021:data<=-16'd564;
      79022:data<=-16'd511;
      79023:data<=-16'd1403;
      79024:data<=-16'd769;
      79025:data<=-16'd194;
      79026:data<=-16'd209;
      79027:data<=-16'd288;
      79028:data<=-16'd1356;
      79029:data<=-16'd2517;
      79030:data<=-16'd3435;
      79031:data<=-16'd3639;
      79032:data<=-16'd3074;
      79033:data<=-16'd3071;
      79034:data<=-16'd2440;
      79035:data<=-16'd2123;
      79036:data<=-16'd2820;
      79037:data<=-16'd1676;
      79038:data<=-16'd1883;
      79039:data<=-16'd3378;
      79040:data<=-16'd1384;
      79041:data<=-16'd4414;
      79042:data<=-16'd14897;
      79043:data<=-16'd18792;
      79044:data<=-16'd16219;
      79045:data<=-16'd15785;
      79046:data<=-16'd14939;
      79047:data<=-16'd13515;
      79048:data<=-16'd14022;
      79049:data<=-16'd13803;
      79050:data<=-16'd12678;
      79051:data<=-16'd11251;
      79052:data<=-16'd9247;
      79053:data<=-16'd9148;
      79054:data<=-16'd10395;
      79055:data<=-16'd10363;
      79056:data<=-16'd9702;
      79057:data<=-16'd9037;
      79058:data<=-16'd8436;
      79059:data<=-16'd7900;
      79060:data<=-16'd7081;
      79061:data<=-16'd6760;
      79062:data<=-16'd6677;
      79063:data<=-16'd6354;
      79064:data<=-16'd6081;
      79065:data<=-16'd5178;
      79066:data<=-16'd5265;
      79067:data<=-16'd6593;
      79068:data<=-16'd6211;
      79069:data<=-16'd5803;
      79070:data<=-16'd5941;
      79071:data<=-16'd4589;
      79072:data<=-16'd4504;
      79073:data<=-16'd4793;
      79074:data<=-16'd3685;
      79075:data<=-16'd4165;
      79076:data<=-16'd3344;
      79077:data<=-16'd1859;
      79078:data<=-16'd3802;
      79079:data<=-16'd367;
      79080:data<=16'd8587;
      79081:data<=16'd10392;
      79082:data<=16'd8114;
      79083:data<=16'd8335;
      79084:data<=16'd8073;
      79085:data<=16'd8176;
      79086:data<=16'd8765;
      79087:data<=16'd8178;
      79088:data<=16'd8436;
      79089:data<=16'd8545;
      79090:data<=16'd7890;
      79091:data<=16'd7473;
      79092:data<=16'd5518;
      79093:data<=16'd4241;
      79094:data<=16'd5344;
      79095:data<=16'd4684;
      79096:data<=16'd2617;
      79097:data<=16'd1988;
      79098:data<=16'd2006;
      79099:data<=16'd2467;
      79100:data<=16'd2855;
      79101:data<=16'd2441;
      79102:data<=16'd2255;
      79103:data<=16'd1992;
      79104:data<=16'd1051;
      79105:data<=16'd352;
      79106:data<=16'd470;
      79107:data<=16'd881;
      79108:data<=16'd1007;
      79109:data<=16'd1371;
      79110:data<=16'd1410;
      79111:data<=16'd919;
      79112:data<=16'd1591;
      79113:data<=16'd1289;
      79114:data<=16'd453;
      79115:data<=16'd2560;
      79116:data<=-16'd714;
      79117:data<=-16'd11391;
      79118:data<=-16'd14932;
      79119:data<=-16'd12076;
      79120:data<=-16'd12310;
      79121:data<=-16'd11887;
      79122:data<=-16'd10789;
      79123:data<=-16'd11336;
      79124:data<=-16'd10002;
      79125:data<=-16'd8974;
      79126:data<=-16'd9130;
      79127:data<=-16'd7915;
      79128:data<=-16'd7464;
      79129:data<=-16'd7251;
      79130:data<=-16'd6490;
      79131:data<=-16'd6649;
      79132:data<=-16'd5718;
      79133:data<=-16'd4610;
      79134:data<=-16'd4880;
      79135:data<=-16'd4228;
      79136:data<=-16'd3647;
      79137:data<=-16'd3665;
      79138:data<=-16'd3052;
      79139:data<=-16'd2939;
      79140:data<=-16'd1997;
      79141:data<=16'd466;
      79142:data<=16'd2208;
      79143:data<=16'd2948;
      79144:data<=16'd2587;
      79145:data<=16'd2343;
      79146:data<=16'd3130;
      79147:data<=16'd2887;
      79148:data<=16'd3289;
      79149:data<=16'd4196;
      79150:data<=16'd2666;
      79151:data<=16'd3280;
      79152:data<=16'd4954;
      79153:data<=16'd3159;
      79154:data<=16'd7817;
      79155:data<=16'd18498;
      79156:data<=16'd20422;
      79157:data<=16'd17638;
      79158:data<=16'd18204;
      79159:data<=16'd17475;
      79160:data<=16'd16695;
      79161:data<=16'd17256;
      79162:data<=16'd15978;
      79163:data<=16'd15362;
      79164:data<=16'd15080;
      79165:data<=16'd13628;
      79166:data<=16'd14404;
      79167:data<=16'd15750;
      79168:data<=16'd15264;
      79169:data<=16'd14944;
      79170:data<=16'd14589;
      79171:data<=16'd13940;
      79172:data<=16'd13540;
      79173:data<=16'd13054;
      79174:data<=16'd12727;
      79175:data<=16'd12236;
      79176:data<=16'd11861;
      79177:data<=16'd11580;
      79178:data<=16'd10965;
      79179:data<=16'd11697;
      79180:data<=16'd12502;
      79181:data<=16'd11664;
      79182:data<=16'd11647;
      79183:data<=16'd11775;
      79184:data<=16'd10463;
      79185:data<=16'd9022;
      79186:data<=16'd7856;
      79187:data<=16'd7756;
      79188:data<=16'd7329;
      79189:data<=16'd6088;
      79190:data<=16'd7321;
      79191:data<=16'd5758;
      79192:data<=-16'd2041;
      79193:data<=-16'd5971;
      79194:data<=-16'd4613;
      79195:data<=-16'd4575;
      79196:data<=-16'd4052;
      79197:data<=-16'd3247;
      79198:data<=-16'd4168;
      79199:data<=-16'd3733;
      79200:data<=-16'd2898;
      79201:data<=-16'd3498;
      79202:data<=-16'd3309;
      79203:data<=-16'd2635;
      79204:data<=-16'd2062;
      79205:data<=-16'd963;
      79206:data<=-16'd567;
      79207:data<=-16'd596;
      79208:data<=-16'd314;
      79209:data<=-16'd429;
      79210:data<=-16'd309;
      79211:data<=-16'd212;
      79212:data<=-16'd660;
      79213:data<=-16'd476;
      79214:data<=-16'd469;
      79215:data<=-16'd754;
      79216:data<=16'd355;
      79217:data<=16'd1801;
      79218:data<=16'd2425;
      79219:data<=16'd2083;
      79220:data<=16'd1521;
      79221:data<=16'd2147;
      79222:data<=16'd1927;
      79223:data<=16'd1387;
      79224:data<=16'd2405;
      79225:data<=16'd1586;
      79226:data<=16'd1544;
      79227:data<=16'd3102;
      79228:data<=16'd1096;
      79229:data<=16'd5835;
      79230:data<=16'd18729;
      79231:data<=16'd20994;
      79232:data<=16'd16894;
      79233:data<=16'd17986;
      79234:data<=16'd17088;
      79235:data<=16'd15312;
      79236:data<=16'd15934;
      79237:data<=16'd14650;
      79238:data<=16'd14031;
      79239:data<=16'd13752;
      79240:data<=16'd12187;
      79241:data<=16'd12930;
      79242:data<=16'd13840;
      79243:data<=16'd13552;
      79244:data<=16'd13490;
      79245:data<=16'd12396;
      79246:data<=16'd11805;
      79247:data<=16'd11634;
      79248:data<=16'd10627;
      79249:data<=16'd10527;
      79250:data<=16'd10125;
      79251:data<=16'd9210;
      79252:data<=16'd9072;
      79253:data<=16'd8542;
      79254:data<=16'd8385;
      79255:data<=16'd8536;
      79256:data<=16'd8395;
      79257:data<=16'd8910;
      79258:data<=16'd8431;
      79259:data<=16'd7454;
      79260:data<=16'd7144;
      79261:data<=16'd6103;
      79262:data<=16'd6067;
      79263:data<=16'd6011;
      79264:data<=16'd4623;
      79265:data<=16'd5562;
      79266:data<=16'd3985;
      79267:data<=-16'd3588;
      79268:data<=-16'd7413;
      79269:data<=-16'd6297;
      79270:data<=-16'd6710;
      79271:data<=-16'd6498;
      79272:data<=-16'd5410;
      79273:data<=-16'd6683;
      79274:data<=-16'd8029;
      79275:data<=-16'd8155;
      79276:data<=-16'd8147;
      79277:data<=-16'd7573;
      79278:data<=-16'd7266;
      79279:data<=-16'd7022;
      79280:data<=-16'd5601;
      79281:data<=-16'd4890;
      79282:data<=-16'd5172;
      79283:data<=-16'd4934;
      79284:data<=-16'd5086;
      79285:data<=-16'd5369;
      79286:data<=-16'd5260;
      79287:data<=-16'd5342;
      79288:data<=-16'd4930;
      79289:data<=-16'd5019;
      79290:data<=-16'd5580;
      79291:data<=-16'd4250;
      79292:data<=-16'd2543;
      79293:data<=-16'd2208;
      79294:data<=-16'd2617;
      79295:data<=-16'd2904;
      79296:data<=-16'd2008;
      79297:data<=-16'd1932;
      79298:data<=-16'd2628;
      79299:data<=-16'd2087;
      79300:data<=-16'd2769;
      79301:data<=-16'd2481;
      79302:data<=-16'd1196;
      79303:data<=-16'd3748;
      79304:data<=-16'd38;
      79305:data<=16'd11793;
      79306:data<=16'd14627;
      79307:data<=16'd11132;
      79308:data<=16'd11106;
      79309:data<=16'd9988;
      79310:data<=16'd9188;
      79311:data<=16'd9612;
      79312:data<=16'd8106;
      79313:data<=16'd8126;
      79314:data<=16'd7970;
      79315:data<=16'd6302;
      79316:data<=16'd7232;
      79317:data<=16'd8081;
      79318:data<=16'd8188;
      79319:data<=16'd9711;
      79320:data<=16'd9652;
      79321:data<=16'd8539;
      79322:data<=16'd8002;
      79323:data<=16'd7027;
      79324:data<=16'd6707;
      79325:data<=16'd6698;
      79326:data<=16'd6038;
      79327:data<=16'd5454;
      79328:data<=16'd5027;
      79329:data<=16'd4687;
      79330:data<=16'd3885;
      79331:data<=16'd3369;
      79332:data<=16'd3536;
      79333:data<=16'd2511;
      79334:data<=16'd2058;
      79335:data<=16'd2743;
      79336:data<=16'd1803;
      79337:data<=16'd1256;
      79338:data<=16'd990;
      79339:data<=-16'd65;
      79340:data<=16'd1394;
      79341:data<=-16'd716;
      79342:data<=-16'd10599;
      79343:data<=-16'd16163;
      79344:data<=-16'd14592;
      79345:data<=-16'd14557;
      79346:data<=-16'd14674;
      79347:data<=-16'd13198;
      79348:data<=-16'd13455;
      79349:data<=-16'd13591;
      79350:data<=-16'd12660;
      79351:data<=-16'd12736;
      79352:data<=-16'd12364;
      79353:data<=-16'd11233;
      79354:data<=-16'd11758;
      79355:data<=-16'd13236;
      79356:data<=-16'd13379;
      79357:data<=-16'd12727;
      79358:data<=-16'd12734;
      79359:data<=-16'd12542;
      79360:data<=-16'd11787;
      79361:data<=-16'd11973;
      79362:data<=-16'd12252;
      79363:data<=-16'd11928;
      79364:data<=-16'd12722;
      79365:data<=-16'd13089;
      79366:data<=-16'd11908;
      79367:data<=-16'd12040;
      79368:data<=-16'd12919;
      79369:data<=-16'd12689;
      79370:data<=-16'd12317;
      79371:data<=-16'd11975;
      79372:data<=-16'd11950;
      79373:data<=-16'd11702;
      79374:data<=-16'd10754;
      79375:data<=-16'd10836;
      79376:data<=-16'd9919;
      79377:data<=-16'd8630;
      79378:data<=-16'd10458;
      79379:data<=-16'd7462;
      79380:data<=16'd1406;
      79381:data<=16'd3319;
      79382:data<=16'd1037;
      79383:data<=16'd1898;
      79384:data<=16'd1007;
      79385:data<=-16'd117;
      79386:data<=16'd849;
      79387:data<=16'd378;
      79388:data<=16'd466;
      79389:data<=16'd743;
      79390:data<=-16'd159;
      79391:data<=16'd600;
      79392:data<=16'd206;
      79393:data<=-16'd1607;
      79394:data<=-16'd922;
      79395:data<=-16'd679;
      79396:data<=-16'd1422;
      79397:data<=-16'd928;
      79398:data<=-16'd1165;
      79399:data<=-16'd1483;
      79400:data<=-16'd1072;
      79401:data<=-16'd1280;
      79402:data<=-16'd1395;
      79403:data<=-16'd1817;
      79404:data<=-16'd3057;
      79405:data<=-16'd4220;
      79406:data<=-16'd4598;
      79407:data<=-16'd3365;
      79408:data<=-16'd2205;
      79409:data<=-16'd2036;
      79410:data<=-16'd1428;
      79411:data<=-16'd1436;
      79412:data<=-16'd1641;
      79413:data<=-16'd1507;
      79414:data<=-16'd2149;
      79415:data<=-16'd1098;
      79416:data<=-16'd2181;
      79417:data<=-16'd10778;
      79418:data<=-16'd17215;
      79419:data<=-16'd16104;
      79420:data<=-16'd15074;
      79421:data<=-16'd14781;
      79422:data<=-16'd13461;
      79423:data<=-16'd13339;
      79424:data<=-16'd12939;
      79425:data<=-16'd11935;
      79426:data<=-16'd11847;
      79427:data<=-16'd11492;
      79428:data<=-16'd11151;
      79429:data<=-16'd11872;
      79430:data<=-16'd12800;
      79431:data<=-16'd12857;
      79432:data<=-16'd12094;
      79433:data<=-16'd11999;
      79434:data<=-16'd11964;
      79435:data<=-16'd10575;
      79436:data<=-16'd9777;
      79437:data<=-16'd9741;
      79438:data<=-16'd9189;
      79439:data<=-16'd9323;
      79440:data<=-16'd8783;
      79441:data<=-16'd7153;
      79442:data<=-16'd7764;
      79443:data<=-16'd9053;
      79444:data<=-16'd8523;
      79445:data<=-16'd7827;
      79446:data<=-16'd7253;
      79447:data<=-16'd7015;
      79448:data<=-16'd6975;
      79449:data<=-16'd6376;
      79450:data<=-16'd6493;
      79451:data<=-16'd5692;
      79452:data<=-16'd5219;
      79453:data<=-16'd8216;
      79454:data<=-16'd5559;
      79455:data<=16'd3692;
      79456:data<=16'd5736;
      79457:data<=16'd3607;
      79458:data<=16'd4837;
      79459:data<=16'd4309;
      79460:data<=16'd3805;
      79461:data<=16'd5112;
      79462:data<=16'd4422;
      79463:data<=16'd4455;
      79464:data<=16'd4883;
      79465:data<=16'd3977;
      79466:data<=16'd4399;
      79467:data<=16'd3791;
      79468:data<=16'd2150;
      79469:data<=16'd2431;
      79470:data<=16'd2423;
      79471:data<=16'd2447;
      79472:data<=16'd2993;
      79473:data<=16'd2397;
      79474:data<=16'd2519;
      79475:data<=16'd2911;
      79476:data<=16'd2279;
      79477:data<=16'd2262;
      79478:data<=16'd2378;
      79479:data<=16'd1591;
      79480:data<=-16'd12;
      79481:data<=-16'd831;
      79482:data<=16'd118;
      79483:data<=-16'd36;
      79484:data<=-16'd408;
      79485:data<=16'd696;
      79486:data<=16'd362;
      79487:data<=16'd391;
      79488:data<=16'd1152;
      79489:data<=16'd23;
      79490:data<=16'd816;
      79491:data<=-16'd65;
      79492:data<=-16'd8364;
      79493:data<=-16'd14301;
      79494:data<=-16'd13676;
      79495:data<=-16'd13400;
      79496:data<=-16'd12546;
      79497:data<=-16'd9823;
      79498:data<=-16'd8486;
      79499:data<=-16'd8178;
      79500:data<=-16'd7961;
      79501:data<=-16'd7685;
      79502:data<=-16'd6954;
      79503:data<=-16'd6554;
      79504:data<=-16'd6827;
      79505:data<=-16'd7752;
      79506:data<=-16'd8314;
      79507:data<=-16'd7503;
      79508:data<=-16'd7235;
      79509:data<=-16'd7341;
      79510:data<=-16'd5927;
      79511:data<=-16'd5150;
      79512:data<=-16'd5348;
      79513:data<=-16'd4807;
      79514:data<=-16'd4807;
      79515:data<=-16'd4384;
      79516:data<=-16'd3033;
      79517:data<=-16'd3432;
      79518:data<=-16'd4000;
      79519:data<=-16'd3694;
      79520:data<=-16'd3971;
      79521:data<=-16'd3400;
      79522:data<=-16'd3011;
      79523:data<=-16'd3154;
      79524:data<=-16'd2085;
      79525:data<=-16'd2340;
      79526:data<=-16'd2149;
      79527:data<=-16'd669;
      79528:data<=-16'd2287;
      79529:data<=16'd579;
      79530:data<=16'd10190;
      79531:data<=16'd13336;
      79532:data<=16'd11570;
      79533:data<=16'd12117;
      79534:data<=16'd11450;
      79535:data<=16'd10968;
      79536:data<=16'd11724;
      79537:data<=16'd11019;
      79538:data<=16'd10705;
      79539:data<=16'd10621;
      79540:data<=16'd10199;
      79541:data<=16'd9649;
      79542:data<=16'd8305;
      79543:data<=16'd9081;
      79544:data<=16'd10440;
      79545:data<=16'd9600;
      79546:data<=16'd9867;
      79547:data<=16'd9683;
      79548:data<=16'd8170;
      79549:data<=16'd8564;
      79550:data<=16'd8381;
      79551:data<=16'd7868;
      79552:data<=16'd8642;
      79553:data<=16'd7577;
      79554:data<=16'd6666;
      79555:data<=16'd8228;
      79556:data<=16'd10097;
      79557:data<=16'd11063;
      79558:data<=16'd10332;
      79559:data<=16'd10003;
      79560:data<=16'd10695;
      79561:data<=16'd9724;
      79562:data<=16'd9285;
      79563:data<=16'd9248;
      79564:data<=16'd8119;
      79565:data<=16'd9107;
      79566:data<=16'd7721;
      79567:data<=16'd1093;
      79568:data<=-16'd1923;
      79569:data<=-16'd737;
      79570:data<=-16'd782;
      79571:data<=-16'd605;
      79572:data<=-16'd230;
      79573:data<=-16'd666;
      79574:data<=-16'd446;
      79575:data<=-16'd368;
      79576:data<=-16'd634;
      79577:data<=-16'd212;
      79578:data<=-16'd33;
      79579:data<=-16'd249;
      79580:data<=16'd364;
      79581:data<=16'd1522;
      79582:data<=16'd1836;
      79583:data<=16'd1481;
      79584:data<=16'd1715;
      79585:data<=16'd2077;
      79586:data<=16'd1944;
      79587:data<=16'd2161;
      79588:data<=16'd2356;
      79589:data<=16'd1962;
      79590:data<=16'd2020;
      79591:data<=16'd2331;
      79592:data<=16'd2737;
      79593:data<=16'd4058;
      79594:data<=16'd4567;
      79595:data<=16'd3911;
      79596:data<=16'd4118;
      79597:data<=16'd4029;
      79598:data<=16'd3750;
      79599:data<=16'd4293;
      79600:data<=16'd3592;
      79601:data<=16'd3573;
      79602:data<=16'd4340;
      79603:data<=16'd2578;
      79604:data<=16'd5130;
      79605:data<=16'd13517;
      79606:data<=16'd16525;
      79607:data<=16'd15027;
      79608:data<=16'd15201;
      79609:data<=16'd14481;
      79610:data<=16'd13517;
      79611:data<=16'd13573;
      79612:data<=16'd12828;
      79613:data<=16'd12251;
      79614:data<=16'd11679;
      79615:data<=16'd10945;
      79616:data<=16'd11016;
      79617:data<=16'd11248;
      79618:data<=16'd12119;
      79619:data<=16'd12414;
      79620:data<=16'd11166;
      79621:data<=16'd11116;
      79622:data<=16'd11027;
      79623:data<=16'd9492;
      79624:data<=16'd9138;
      79625:data<=16'd9077;
      79626:data<=16'd8476;
      79627:data<=16'd8545;
      79628:data<=16'd7900;
      79629:data<=16'd6810;
      79630:data<=16'd7392;
      79631:data<=16'd9007;
      79632:data<=16'd9307;
      79633:data<=16'd8046;
      79634:data<=16'd7635;
      79635:data<=16'd7582;
      79636:data<=16'd6520;
      79637:data<=16'd6516;
      79638:data<=16'd6328;
      79639:data<=16'd5063;
      79640:data<=16'd5829;
      79641:data<=16'd4962;
      79642:data<=-16'd513;
      79643:data<=-16'd4167;
      79644:data<=-16'd4167;
      79645:data<=-16'd3865;
      79646:data<=-16'd3378;
      79647:data<=-16'd3456;
      79648:data<=-16'd4200;
      79649:data<=-16'd3891;
      79650:data<=-16'd3433;
      79651:data<=-16'd3500;
      79652:data<=-16'd3571;
      79653:data<=-16'd4168;
      79654:data<=-16'd4281;
      79655:data<=-16'd2886;
      79656:data<=-16'd1565;
      79657:data<=-16'd1409;
      79658:data<=-16'd1794;
      79659:data<=-16'd1764;
      79660:data<=-16'd1283;
      79661:data<=-16'd1343;
      79662:data<=-16'd1666;
      79663:data<=-16'd1604;
      79664:data<=-16'd1692;
      79665:data<=-16'd1760;
      79666:data<=-16'd1712;
      79667:data<=-16'd1336;
      79668:data<=16'd117;
      79669:data<=16'd895;
      79670:data<=16'd438;
      79671:data<=16'd664;
      79672:data<=16'd599;
      79673:data<=16'd328;
      79674:data<=16'd872;
      79675:data<=16'd372;
      79676:data<=16'd361;
      79677:data<=16'd860;
      79678:data<=-16'd895;
      79679:data<=16'd1579;
      79680:data<=16'd9922;
      79681:data<=16'd13332;
      79682:data<=16'd11794;
      79683:data<=16'd11852;
      79684:data<=16'd11449;
      79685:data<=16'd10336;
      79686:data<=16'd10304;
      79687:data<=16'd9611;
      79688:data<=16'd8813;
      79689:data<=16'd8768;
      79690:data<=16'd8285;
      79691:data<=16'd7708;
      79692:data<=16'd7955;
      79693:data<=16'd8890;
      79694:data<=16'd9212;
      79695:data<=16'd8627;
      79696:data<=16'd8334;
      79697:data<=16'd7629;
      79698:data<=16'd6511;
      79699:data<=16'd6475;
      79700:data<=16'd6332;
      79701:data<=16'd5780;
      79702:data<=16'd5792;
      79703:data<=16'd5059;
      79704:data<=16'd4387;
      79705:data<=16'd5427;
      79706:data<=16'd6203;
      79707:data<=16'd5718;
      79708:data<=16'd5303;
      79709:data<=16'd5410;
      79710:data<=16'd5143;
      79711:data<=16'd3785;
      79712:data<=16'd2955;
      79713:data<=16'd3215;
      79714:data<=16'd3040;
      79715:data<=16'd3325;
      79716:data<=16'd2461;
      79717:data<=-16'd2678;
      79718:data<=-16'd6959;
      79719:data<=-16'd6578;
      79720:data<=-16'd6123;
      79721:data<=-16'd6666;
      79722:data<=-16'd6341;
      79723:data<=-16'd6302;
      79724:data<=-16'd6625;
      79725:data<=-16'd6717;
      79726:data<=-16'd6575;
      79727:data<=-16'd6143;
      79728:data<=-16'd6219;
      79729:data<=-16'd6351;
      79730:data<=-16'd6246;
      79731:data<=-16'd6692;
      79732:data<=-16'd6457;
      79733:data<=-16'd5844;
      79734:data<=-16'd6217;
      79735:data<=-16'd5973;
      79736:data<=-16'd5585;
      79737:data<=-16'd6334;
      79738:data<=-16'd6334;
      79739:data<=-16'd5883;
      79740:data<=-16'd6200;
      79741:data<=-16'd5994;
      79742:data<=-16'd5518;
      79743:data<=-16'd6308;
      79744:data<=-16'd7782;
      79745:data<=-16'd7797;
      79746:data<=-16'd6784;
      79747:data<=-16'd7248;
      79748:data<=-16'd7517;
      79749:data<=-16'd6687;
      79750:data<=-16'd7379;
      79751:data<=-16'd7045;
      79752:data<=-16'd5944;
      79753:data<=-16'd7741;
      79754:data<=-16'd5060;
      79755:data<=16'd2657;
      79756:data<=16'd3404;
      79757:data<=16'd920;
      79758:data<=16'd2393;
      79759:data<=16'd1541;
      79760:data<=-16'd317;
      79761:data<=16'd928;
      79762:data<=16'd664;
      79763:data<=-16'd194;
      79764:data<=16'd443;
      79765:data<=-16'd33;
      79766:data<=-16'd83;
      79767:data<=16'd485;
      79768:data<=-16'd1019;
      79769:data<=-16'd2698;
      79770:data<=-16'd2575;
      79771:data<=-16'd2200;
      79772:data<=-16'd2775;
      79773:data<=-16'd3195;
      79774:data<=-16'd2781;
      79775:data<=-16'd2631;
      79776:data<=-16'd2190;
      79777:data<=-16'd1645;
      79778:data<=-16'd2447;
      79779:data<=-16'd2608;
      79780:data<=-16'd2522;
      79781:data<=-16'd4432;
      79782:data<=-16'd5571;
      79783:data<=-16'd5318;
      79784:data<=-16'd5192;
      79785:data<=-16'd4526;
      79786:data<=-16'd4819;
      79787:data<=-16'd5391;
      79788:data<=-16'd4526;
      79789:data<=-16'd4517;
      79790:data<=-16'd4337;
      79791:data<=-16'd4414;
      79792:data<=-16'd9291;
      79793:data<=-16'd15060;
      79794:data<=-16'd16301;
      79795:data<=-16'd15497;
      79796:data<=-16'd14945;
      79797:data<=-16'd14827;
      79798:data<=-16'd14728;
      79799:data<=-16'd13972;
      79800:data<=-16'd13406;
      79801:data<=-16'd12827;
      79802:data<=-16'd12122;
      79803:data<=-16'd12031;
      79804:data<=-16'd11376;
      79805:data<=-16'd11019;
      79806:data<=-16'd12340;
      79807:data<=-16'd12756;
      79808:data<=-16'd11834;
      79809:data<=-16'd11458;
      79810:data<=-16'd11082;
      79811:data<=-16'd10689;
      79812:data<=-16'd10602;
      79813:data<=-16'd10002;
      79814:data<=-16'd9465;
      79815:data<=-16'd9580;
      79816:data<=-16'd9532;
      79817:data<=-16'd9015;
      79818:data<=-16'd8793;
      79819:data<=-16'd9329;
      79820:data<=-16'd9339;
      79821:data<=-16'd8684;
      79822:data<=-16'd8819;
      79823:data<=-16'd8196;
      79824:data<=-16'd6975;
      79825:data<=-16'd7548;
      79826:data<=-16'd6980;
      79827:data<=-16'd5977;
      79828:data<=-16'd7662;
      79829:data<=-16'd4723;
      79830:data<=16'd2466;
      79831:data<=16'd3295;
      79832:data<=16'd1524;
      79833:data<=16'd2359;
      79834:data<=16'd1744;
      79835:data<=16'd1662;
      79836:data<=16'd2631;
      79837:data<=16'd2055;
      79838:data<=16'd2907;
      79839:data<=16'd3560;
      79840:data<=16'd1921;
      79841:data<=16'd1823;
      79842:data<=16'd2557;
      79843:data<=16'd1845;
      79844:data<=16'd381;
      79845:data<=-16'd617;
      79846:data<=16'd494;
      79847:data<=16'd1416;
      79848:data<=16'd505;
      79849:data<=16'd567;
      79850:data<=16'd1045;
      79851:data<=16'd907;
      79852:data<=16'd1074;
      79853:data<=16'd919;
      79854:data<=16'd957;
      79855:data<=16'd581;
      79856:data<=-16'd977;
      79857:data<=-16'd1475;
      79858:data<=-16'd1428;
      79859:data<=-16'd1509;
      79860:data<=-16'd831;
      79861:data<=-16'd1151;
      79862:data<=-16'd1365;
      79863:data<=-16'd350;
      79864:data<=-16'd772;
      79865:data<=-16'd561;
      79866:data<=16'd308;
      79867:data<=-16'd4247;
      79868:data<=-16'd11047;
      79869:data<=-16'd12747;
      79870:data<=-16'd11759;
      79871:data<=-16'd11233;
      79872:data<=-16'd10191;
      79873:data<=-16'd9588;
      79874:data<=-16'd9749;
      79875:data<=-16'd9417;
      79876:data<=-16'd8666;
      79877:data<=-16'd7888;
      79878:data<=-16'd7661;
      79879:data<=-16'd7533;
      79880:data<=-16'd7037;
      79881:data<=-16'd7814;
      79882:data<=-16'd8551;
      79883:data<=-16'd7711;
      79884:data<=-16'd7711;
      79885:data<=-16'd7520;
      79886:data<=-16'd6323;
      79887:data<=-16'd6549;
      79888:data<=-16'd6120;
      79889:data<=-16'd4778;
      79890:data<=-16'd5222;
      79891:data<=-16'd5404;
      79892:data<=-16'd4675;
      79893:data<=-16'd4575;
      79894:data<=-16'd5065;
      79895:data<=-16'd5600;
      79896:data<=-16'd4560;
      79897:data<=-16'd3792;
      79898:data<=-16'd4581;
      79899:data<=-16'd3835;
      79900:data<=-16'd3101;
      79901:data<=-16'd2864;
      79902:data<=-16'd2149;
      79903:data<=-16'd3771;
      79904:data<=-16'd1521;
      79905:data<=16'd6907;
      79906:data<=16'd9544;
      79907:data<=16'd6808;
      79908:data<=16'd6329;
      79909:data<=16'd6250;
      79910:data<=16'd6589;
      79911:data<=16'd7271;
      79912:data<=16'd6573;
      79913:data<=16'd6581;
      79914:data<=16'd6449;
      79915:data<=16'd5318;
      79916:data<=16'd5356;
      79917:data<=16'd5786;
      79918:data<=16'd4971;
      79919:data<=16'd3482;
      79920:data<=16'd3331;
      79921:data<=16'd4131;
      79922:data<=16'd3460;
      79923:data<=16'd2927;
      79924:data<=16'd3626;
      79925:data<=16'd3747;
      79926:data<=16'd3485;
      79927:data<=16'd3140;
      79928:data<=16'd3410;
      79929:data<=16'd4255;
      79930:data<=16'd3856;
      79931:data<=16'd3673;
      79932:data<=16'd4035;
      79933:data<=16'd3344;
      79934:data<=16'd3369;
      79935:data<=16'd3970;
      79936:data<=16'd3833;
      79937:data<=16'd3962;
      79938:data<=16'd3774;
      79939:data<=16'd3242;
      79940:data<=16'd4044;
      79941:data<=16'd4441;
      79942:data<=-16'd67;
      79943:data<=-16'd6463;
      79944:data<=-16'd6185;
      79945:data<=-16'd3363;
      79946:data<=-16'd4911;
      79947:data<=-16'd5037;
      79948:data<=-16'd3504;
      79949:data<=-16'd4328;
      79950:data<=-16'd3670;
      79951:data<=-16'd2561;
      79952:data<=-16'd2980;
      79953:data<=-16'd2268;
      79954:data<=-16'd1999;
      79955:data<=-16'd2167;
      79956:data<=-16'd899;
      79957:data<=16'd409;
      79958:data<=16'd870;
      79959:data<=16'd440;
      79960:data<=16'd682;
      79961:data<=16'd1597;
      79962:data<=16'd1568;
      79963:data<=16'd2335;
      79964:data<=16'd2591;
      79965:data<=16'd1404;
      79966:data<=16'd1703;
      79967:data<=16'd1685;
      79968:data<=16'd1909;
      79969:data<=16'd3921;
      79970:data<=16'd3965;
      79971:data<=16'd3715;
      79972:data<=16'd4545;
      79973:data<=16'd4053;
      79974:data<=16'd3771;
      79975:data<=16'd3673;
      79976:data<=16'd4235;
      79977:data<=16'd4605;
      79978:data<=16'd2394;
      79979:data<=16'd4965;
      79980:data<=16'd12330;
      79981:data<=16'd14742;
      79982:data<=16'd14924;
      79983:data<=16'd15412;
      79984:data<=16'd13960;
      79985:data<=16'd13599;
      79986:data<=16'd13775;
      79987:data<=16'd13587;
      79988:data<=16'd13315;
      79989:data<=16'd11362;
      79990:data<=16'd10834;
      79991:data<=16'd11471;
      79992:data<=16'd10592;
      79993:data<=16'd10777;
      79994:data<=16'd11094;
      79995:data<=16'd10748;
      79996:data<=16'd11021;
      79997:data<=16'd10319;
      79998:data<=16'd10026;
      79999:data<=16'd9849;
      80000:data<=16'd8296;
      80001:data<=16'd8583;
      80002:data<=16'd9235;
      80003:data<=16'd8150;
      80004:data<=16'd7955;
      80005:data<=16'd7938;
      80006:data<=16'd8005;
      80007:data<=16'd9112;
      80008:data<=16'd8947;
      80009:data<=16'd7937;
      80010:data<=16'd7879;
      80011:data<=16'd7790;
      80012:data<=16'd7385;
      80013:data<=16'd6743;
      80014:data<=16'd5234;
      80015:data<=16'd5224;
      80016:data<=16'd6884;
      80017:data<=16'd3136;
      80018:data<=-16'd4215;
      80019:data<=-16'd4928;
      80020:data<=-16'd2566;
      80021:data<=-16'd3010;
      80022:data<=-16'd2875;
      80023:data<=-16'd2984;
      80024:data<=-16'd3127;
      80025:data<=-16'd2008;
      80026:data<=-16'd2958;
      80027:data<=-16'd3243;
      80028:data<=-16'd1850;
      80029:data<=-16'd2391;
      80030:data<=-16'd2064;
      80031:data<=-16'd628;
      80032:data<=-16'd14;
      80033:data<=16'd848;
      80034:data<=16'd755;
      80035:data<=16'd876;
      80036:data<=16'd1339;
      80037:data<=-16'd64;
      80038:data<=-16'd496;
      80039:data<=16'd244;
      80040:data<=16'd223;
      80041:data<=16'd143;
      80042:data<=-16'd331;
      80043:data<=16'd91;
      80044:data<=16'd807;
      80045:data<=16'd748;
      80046:data<=16'd1977;
      80047:data<=16'd1903;
      80048:data<=16'd899;
      80049:data<=16'd1609;
      80050:data<=16'd610;
      80051:data<=16'd699;
      80052:data<=16'd2311;
      80053:data<=16'd252;
      80054:data<=16'd1861;
      80055:data<=16'd8877;
      80056:data<=16'd11859;
      80057:data<=16'd12078;
      80058:data<=16'd12552;
      80059:data<=16'd12188;
      80060:data<=16'd11632;
      80061:data<=16'd10050;
      80062:data<=16'd9312;
      80063:data<=16'd10366;
      80064:data<=16'd9696;
      80065:data<=16'd7864;
      80066:data<=16'd6960;
      80067:data<=16'd7236;
      80068:data<=16'd8190;
      80069:data<=16'd7915;
      80070:data<=16'd7191;
      80071:data<=16'd7547;
      80072:data<=16'd7891;
      80073:data<=16'd7582;
      80074:data<=16'd6831;
      80075:data<=16'd6140;
      80076:data<=16'd5424;
      80077:data<=16'd5124;
      80078:data<=16'd6072;
      80079:data<=16'd5702;
      80080:data<=16'd3946;
      80081:data<=16'd4637;
      80082:data<=16'd6208;
      80083:data<=16'd5821;
      80084:data<=16'd5328;
      80085:data<=16'd5607;
      80086:data<=16'd5122;
      80087:data<=16'd4657;
      80088:data<=16'd5298;
      80089:data<=16'd4114;
      80090:data<=16'd2482;
      80091:data<=16'd3823;
      80092:data<=16'd728;
      80093:data<=-16'd7195;
      80094:data<=-16'd8205;
      80095:data<=-16'd5222;
      80096:data<=-16'd5868;
      80097:data<=-16'd6156;
      80098:data<=-16'd5504;
      80099:data<=-16'd6178;
      80100:data<=-16'd6467;
      80101:data<=-16'd6037;
      80102:data<=-16'd5883;
      80103:data<=-16'd6159;
      80104:data<=-16'd5841;
      80105:data<=-16'd5369;
      80106:data<=-16'd4790;
      80107:data<=-16'd2322;
      80108:data<=-16'd1621;
      80109:data<=-16'd3668;
      80110:data<=-16'd3385;
      80111:data<=-16'd2761;
      80112:data<=-16'd2995;
      80113:data<=-16'd2303;
      80114:data<=-16'd3112;
      80115:data<=-16'd3151;
      80116:data<=-16'd2182;
      80117:data<=-16'd3515;
      80118:data<=-16'd3374;
      80119:data<=-16'd2088;
      80120:data<=-16'd1589;
      80121:data<=-16'd92;
      80122:data<=-16'd836;
      80123:data<=-16'd1789;
      80124:data<=-16'd325;
      80125:data<=-16'd1048;
      80126:data<=-16'd1049;
      80127:data<=-16'd317;
      80128:data<=-16'd2379;
      80129:data<=16'd590;
      80130:data<=16'd7521;
      80131:data<=16'd9145;
      80132:data<=16'd8061;
      80133:data<=16'd7517;
      80134:data<=16'd7397;
      80135:data<=16'd7650;
      80136:data<=16'd6208;
      80137:data<=16'd5312;
      80138:data<=16'd6166;
      80139:data<=16'd5824;
      80140:data<=16'd5281;
      80141:data<=16'd4940;
      80142:data<=16'd3882;
      80143:data<=16'd3489;
      80144:data<=16'd2736;
      80145:data<=16'd904;
      80146:data<=-16'd39;
      80147:data<=16'd0;
      80148:data<=16'd450;
      80149:data<=16'd1274;
      80150:data<=16'd1227;
      80151:data<=16'd77;
      80152:data<=-16'd519;
      80153:data<=-16'd466;
      80154:data<=-16'd318;
      80155:data<=16'd211;
      80156:data<=-16'd641;
      80157:data<=-16'd2863;
      80158:data<=-16'd3353;
      80159:data<=-16'd2949;
      80160:data<=-16'd3192;
      80161:data<=-16'd3295;
      80162:data<=-16'd3439;
      80163:data<=-16'd3037;
      80164:data<=-16'd3151;
      80165:data<=-16'd4167;
      80166:data<=-16'd3597;
      80167:data<=-16'd5732;
      80168:data<=-16'd12141;
      80169:data<=-16'd14938;
      80170:data<=-16'd14559;
      80171:data<=-16'd15114;
      80172:data<=-16'd15015;
      80173:data<=-16'd14938;
      80174:data<=-16'd14421;
      80175:data<=-16'd13209;
      80176:data<=-16'd13335;
      80177:data<=-16'd12446;
      80178:data<=-16'd11142;
      80179:data<=-16'd11230;
      80180:data<=-16'd10257;
      80181:data<=-16'd10577;
      80182:data<=-16'd12296;
      80183:data<=-16'd11512;
      80184:data<=-16'd11094;
      80185:data<=-16'd11914;
      80186:data<=-16'd11579;
      80187:data<=-16'd10827;
      80188:data<=-16'd9743;
      80189:data<=-16'd9800;
      80190:data<=-16'd10402;
      80191:data<=-16'd9051;
      80192:data<=-16'd8909;
      80193:data<=-16'd9802;
      80194:data<=-16'd9304;
      80195:data<=-16'd9644;
      80196:data<=-16'd9606;
      80197:data<=-16'd8877;
      80198:data<=-16'd9044;
      80199:data<=-16'd8252;
      80200:data<=-16'd8229;
      80201:data<=-16'd8484;
      80202:data<=-16'd7206;
      80203:data<=-16'd8416;
      80204:data<=-16'd7086;
      80205:data<=16'd547;
      80206:data<=16'd4061;
      80207:data<=16'd2811;
      80208:data<=16'd2470;
      80209:data<=16'd1383;
      80210:data<=16'd1720;
      80211:data<=16'd3055;
      80212:data<=16'd1754;
      80213:data<=16'd1372;
      80214:data<=16'd1909;
      80215:data<=16'd1362;
      80216:data<=16'd2176;
      80217:data<=16'd2485;
      80218:data<=16'd1457;
      80219:data<=16'd1239;
      80220:data<=-16'd180;
      80221:data<=-16'd1506;
      80222:data<=-16'd265;
      80223:data<=-16'd47;
      80224:data<=-16'd1174;
      80225:data<=-16'd758;
      80226:data<=16'd117;
      80227:data<=16'd311;
      80228:data<=-16'd215;
      80229:data<=-16'd1021;
      80230:data<=-16'd723;
      80231:data<=-16'd723;
      80232:data<=-16'd2173;
      80233:data<=-16'd3083;
      80234:data<=-16'd3065;
      80235:data<=-16'd2464;
      80236:data<=-16'd1848;
      80237:data<=-16'd2441;
      80238:data<=-16'd2493;
      80239:data<=-16'd1612;
      80240:data<=-16'd995;
      80241:data<=-16'd14;
      80242:data<=-16'd2742;
      80243:data<=-16'd9914;
      80244:data<=-16'd13153;
      80245:data<=-16'd12016;
      80246:data<=-16'd11426;
      80247:data<=-16'd11204;
      80248:data<=-16'd11773;
      80249:data<=-16'd11808;
      80250:data<=-16'd10402;
      80251:data<=-16'd10217;
      80252:data<=-16'd9574;
      80253:data<=-16'd8536;
      80254:data<=-16'd9182;
      80255:data<=-16'd8264;
      80256:data<=-16'd7239;
      80257:data<=-16'd8931;
      80258:data<=-16'd9633;
      80259:data<=-16'd9066;
      80260:data<=-16'd8981;
      80261:data<=-16'd8507;
      80262:data<=-16'd7644;
      80263:data<=-16'd6628;
      80264:data<=-16'd6223;
      80265:data<=-16'd6012;
      80266:data<=-16'd5403;
      80267:data<=-16'd5682;
      80268:data<=-16'd5389;
      80269:data<=-16'd4871;
      80270:data<=-16'd6018;
      80271:data<=-16'd5956;
      80272:data<=-16'd5184;
      80273:data<=-16'd5298;
      80274:data<=-16'd4548;
      80275:data<=-16'd4513;
      80276:data<=-16'd4132;
      80277:data<=-16'd2732;
      80278:data<=-16'd3583;
      80279:data<=-16'd1471;
      80280:data<=16'd5166;
      80281:data<=16'd7633;
      80282:data<=16'd6472;
      80283:data<=16'd6246;
      80284:data<=16'd5988;
      80285:data<=16'd5773;
      80286:data<=16'd5486;
      80287:data<=16'd5101;
      80288:data<=16'd5597;
      80289:data<=16'd6018;
      80290:data<=16'd5791;
      80291:data<=16'd5473;
      80292:data<=16'd5830;
      80293:data<=16'd6566;
      80294:data<=16'd5934;
      80295:data<=16'd4461;
      80296:data<=16'd3755;
      80297:data<=16'd3603;
      80298:data<=16'd3369;
      80299:data<=16'd3371;
      80300:data<=16'd3865;
      80301:data<=16'd3307;
      80302:data<=16'd2754;
      80303:data<=16'd4155;
      80304:data<=16'd4061;
      80305:data<=16'd3083;
      80306:data<=16'd4372;
      80307:data<=16'd3703;
      80308:data<=16'd1163;
      80309:data<=16'd970;
      80310:data<=16'd1240;
      80311:data<=16'd1137;
      80312:data<=16'd1868;
      80313:data<=16'd2146;
      80314:data<=16'd936;
      80315:data<=16'd792;
      80316:data<=16'd2822;
      80317:data<=-16'd382;
      80318:data<=-16'd8147;
      80319:data<=-16'd9882;
      80320:data<=-16'd9297;
      80321:data<=-16'd10637;
      80322:data<=-16'd9494;
      80323:data<=-16'd9480;
      80324:data<=-16'd9843;
      80325:data<=-16'd7429;
      80326:data<=-16'd7075;
      80327:data<=-16'd7015;
      80328:data<=-16'd6190;
      80329:data<=-16'd6419;
      80330:data<=-16'd5001;
      80331:data<=-16'd5062;
      80332:data<=-16'd5873;
      80333:data<=-16'd4206;
      80334:data<=-16'd4831;
      80335:data<=-16'd5143;
      80336:data<=-16'd3785;
      80337:data<=-16'd4493;
      80338:data<=-16'd3163;
      80339:data<=-16'd2158;
      80340:data<=-16'd3610;
      80341:data<=-16'd2507;
      80342:data<=-16'd2366;
      80343:data<=-16'd2687;
      80344:data<=-16'd373;
      80345:data<=16'd223;
      80346:data<=16'd320;
      80347:data<=16'd138;
      80348:data<=-16'd543;
      80349:data<=16'd1342;
      80350:data<=16'd1004;
      80351:data<=16'd177;
      80352:data<=16'd2485;
      80353:data<=16'd1124;
      80354:data<=16'd1759;
      80355:data<=16'd9480;
      80356:data<=16'd13247;
      80357:data<=16'd12960;
      80358:data<=16'd15177;
      80359:data<=16'd16880;
      80360:data<=16'd16028;
      80361:data<=16'd14880;
      80362:data<=16'd14628;
      80363:data<=16'd13888;
      80364:data<=16'd12836;
      80365:data<=16'd13068;
      80366:data<=16'd13001;
      80367:data<=16'd12363;
      80368:data<=16'd11647;
      80369:data<=16'd10945;
      80370:data<=16'd12334;
      80371:data<=16'd13273;
      80372:data<=16'd12091;
      80373:data<=16'd12022;
      80374:data<=16'd11546;
      80375:data<=16'd10384;
      80376:data<=16'd10555;
      80377:data<=16'd10103;
      80378:data<=16'd9897;
      80379:data<=16'd10645;
      80380:data<=16'd10187;
      80381:data<=16'd9653;
      80382:data<=16'd10211;
      80383:data<=16'd10947;
      80384:data<=16'd10378;
      80385:data<=16'd9139;
      80386:data<=16'd9538;
      80387:data<=16'd9448;
      80388:data<=16'd7579;
      80389:data<=16'd6467;
      80390:data<=16'd7401;
      80391:data<=16'd9691;
      80392:data<=16'd7197;
      80393:data<=-16'd558;
      80394:data<=-16'd3272;
      80395:data<=-16'd1618;
      80396:data<=-16'd1327;
      80397:data<=-16'd229;
      80398:data<=-16'd100;
      80399:data<=-16'd1024;
      80400:data<=16'd82;
      80401:data<=16'd406;
      80402:data<=16'd218;
      80403:data<=16'd1136;
      80404:data<=16'd1424;
      80405:data<=16'd1130;
      80406:data<=16'd42;
      80407:data<=16'd85;
      80408:data<=16'd2685;
      80409:data<=16'd3888;
      80410:data<=16'd2901;
      80411:data<=16'd1237;
      80412:data<=16'd26;
      80413:data<=16'd1372;
      80414:data<=16'd2729;
      80415:data<=16'd2381;
      80416:data<=16'd2147;
      80417:data<=16'd961;
      80418:data<=16'd100;
      80419:data<=16'd1519;
      80420:data<=16'd2611;
      80421:data<=16'd2914;
      80422:data<=16'd3748;
      80423:data<=16'd4187;
      80424:data<=16'd3586;
      80425:data<=16'd3133;
      80426:data<=16'd3586;
      80427:data<=16'd3011;
      80428:data<=16'd1694;
      80429:data<=16'd3829;
      80430:data<=16'd9488;
      80431:data<=16'd13699;
      80432:data<=16'd13741;
      80433:data<=16'd13191;
      80434:data<=16'd15317;
      80435:data<=16'd15985;
      80436:data<=16'd13593;
      80437:data<=16'd12944;
      80438:data<=16'd13367;
      80439:data<=16'd11489;
      80440:data<=16'd9702;
      80441:data<=16'd10314;
      80442:data<=16'd10915;
      80443:data<=16'd9633;
      80444:data<=16'd8906;
      80445:data<=16'd9679;
      80446:data<=16'd9559;
      80447:data<=16'd9414;
      80448:data<=16'd10392;
      80449:data<=16'd9708;
      80450:data<=16'd7523;
      80451:data<=16'd7380;
      80452:data<=16'd8481;
      80453:data<=16'd7541;
      80454:data<=16'd5758;
      80455:data<=16'd5007;
      80456:data<=16'd4346;
      80457:data<=16'd4783;
      80458:data<=16'd6229;
      80459:data<=16'd6296;
      80460:data<=16'd5852;
      80461:data<=16'd5379;
      80462:data<=16'd5054;
      80463:data<=16'd5230;
      80464:data<=16'd3436;
      80465:data<=16'd3397;
      80466:data<=16'd6548;
      80467:data<=16'd2209;
      80468:data<=-16'd7269;
      80469:data<=-16'd8822;
      80470:data<=-16'd5647;
      80471:data<=-16'd5245;
      80472:data<=-16'd6088;
      80473:data<=-16'd5993;
      80474:data<=-16'd5039;
      80475:data<=-16'd4293;
      80476:data<=-16'd3436;
      80477:data<=-16'd2927;
      80478:data<=-16'd3982;
      80479:data<=-16'd3794;
      80480:data<=-16'd3389;
      80481:data<=-16'd5545;
      80482:data<=-16'd5571;
      80483:data<=-16'd3357;
      80484:data<=-16'd2974;
      80485:data<=-16'd2338;
      80486:data<=-16'd1882;
      80487:data<=-16'd3107;
      80488:data<=-16'd3189;
      80489:data<=-16'd3125;
      80490:data<=-16'd4303;
      80491:data<=-16'd3891;
      80492:data<=-16'd2690;
      80493:data<=-16'd3664;
      80494:data<=-16'd4252;
      80495:data<=-16'd1720;
      80496:data<=-16'd341;
      80497:data<=-16'd2071;
      80498:data<=-16'd1512;
      80499:data<=16'd741;
      80500:data<=-16'd646;
      80501:data<=-16'd2505;
      80502:data<=-16'd1650;
      80503:data<=-16'd1871;
      80504:data<=-16'd1149;
      80505:data<=16'd4881;
      80506:data<=16'd9570;
      80507:data<=16'd8907;
      80508:data<=16'd9794;
      80509:data<=16'd11594;
      80510:data<=16'd9462;
      80511:data<=16'd7943;
      80512:data<=16'd7882;
      80513:data<=16'd5965;
      80514:data<=16'd5714;
      80515:data<=16'd6805;
      80516:data<=16'd5501;
      80517:data<=16'd4907;
      80518:data<=16'd5685;
      80519:data<=16'd4608;
      80520:data<=16'd4241;
      80521:data<=16'd6449;
      80522:data<=16'd6443;
      80523:data<=16'd3920;
      80524:data<=16'd4259;
      80525:data<=16'd5198;
      80526:data<=16'd3312;
      80527:data<=16'd3409;
      80528:data<=16'd5234;
      80529:data<=16'd4726;
      80530:data<=16'd3891;
      80531:data<=16'd3228;
      80532:data<=16'd2911;
      80533:data<=16'd3204;
      80534:data<=16'd1353;
      80535:data<=16'd399;
      80536:data<=16'd837;
      80537:data<=-16'd1057;
      80538:data<=-16'd253;
      80539:data<=16'd1162;
      80540:data<=-16'd2707;
      80541:data<=-16'd5471;
      80542:data<=-16'd9552;
      80543:data<=-16'd17861;
      80544:data<=-16'd19855;
      80545:data<=-16'd18069;
      80546:data<=-16'd18562;
      80547:data<=-16'd17920;
      80548:data<=-16'd19133;
      80549:data<=-16'd19415;
      80550:data<=-16'd15411;
      80551:data<=-16'd16930;
      80552:data<=-16'd21892;
      80553:data<=-16'd22495;
      80554:data<=-16'd22868;
      80555:data<=-16'd22556;
      80556:data<=-16'd21003;
      80557:data<=-16'd22331;
      80558:data<=-16'd22600;
      80559:data<=-16'd20375;
      80560:data<=-16'd19409;
      80561:data<=-16'd16995;
      80562:data<=-16'd13723;
      80563:data<=-16'd15167;
      80564:data<=-16'd17106;
      80565:data<=-16'd14436;
      80566:data<=-16'd13444;
      80567:data<=-16'd15723;
      80568:data<=-16'd14880;
      80569:data<=-16'd12319;
      80570:data<=-16'd10787;
      80571:data<=-16'd9899;
      80572:data<=-16'd11323;
      80573:data<=-16'd11016;
      80574:data<=-16'd8677;
      80575:data<=-16'd14478;
      80576:data<=-16'd26821;
      80577:data<=-16'd32878;
      80578:data<=-16'd26715;
      80579:data<=-16'd13585;
      80580:data<=-16'd7022;
      80581:data<=-16'd12751;
      80582:data<=-16'd21353;
      80583:data<=-16'd21325;
      80584:data<=-16'd11388;
      80585:data<=-16'd5565;
      80586:data<=-16'd11301;
      80587:data<=-16'd15738;
      80588:data<=-16'd14645;
      80589:data<=-16'd12819;
      80590:data<=-16'd7457;
      80591:data<=-16'd5278;
      80592:data<=-16'd9295;
      80593:data<=-16'd1500;
      80594:data<=16'd15575;
      80595:data<=16'd15773;
      80596:data<=16'd2632;
      80597:data<=-16'd1005;
      80598:data<=16'd3580;
      80599:data<=16'd7608;
      80600:data<=16'd10542;
      80601:data<=16'd6478;
      80602:data<=-16'd1384;
      80603:data<=16'd825;
      80604:data<=16'd10237;
      80605:data<=16'd13368;
      80606:data<=16'd6934;
      80607:data<=16'd1336;
      80608:data<=16'd4417;
      80609:data<=16'd6393;
      80610:data<=16'd5221;
      80611:data<=16'd7385;
      80612:data<=16'd3154;
      80613:data<=-16'd981;
      80614:data<=16'd7850;
      80615:data<=16'd6213;
      80616:data<=-16'd8047;
      80617:data<=-16'd5448;
      80618:data<=16'd2487;
      80619:data<=-16'd3240;
      80620:data<=-16'd6097;
      80621:data<=-16'd2927;
      80622:data<=-16'd3774;
      80623:data<=-16'd1089;
      80624:data<=16'd4379;
      80625:data<=16'd2999;
      80626:data<=16'd3277;
      80627:data<=16'd8011;
      80628:data<=16'd3004;
      80629:data<=-16'd8740;
      80630:data<=-16'd12654;
      80631:data<=-16'd10742;
      80632:data<=-16'd10662;
      80633:data<=-16'd8044;
      80634:data<=-16'd654;
      80635:data<=-16'd5767;
      80636:data<=-16'd24272;
      80637:data<=-16'd26530;
      80638:data<=-16'd17764;
      80639:data<=-16'd22747;
      80640:data<=-16'd25927;
      80641:data<=-16'd21270;
      80642:data<=-16'd21106;
      80643:data<=-16'd16474;
      80644:data<=-16'd12216;
      80645:data<=-16'd16997;
      80646:data<=-16'd17805;
      80647:data<=-16'd14193;
      80648:data<=-16'd11858;
      80649:data<=-16'd12595;
      80650:data<=-16'd16048;
      80651:data<=-16'd13016;
      80652:data<=-16'd11767;
      80653:data<=-16'd15412;
      80654:data<=-16'd7573;
      80655:data<=-16'd4006;
      80656:data<=-16'd14277;
      80657:data<=-16'd15282;
      80658:data<=-16'd11600;
      80659:data<=-16'd11539;
      80660:data<=-16'd6357;
      80661:data<=-16'd7197;
      80662:data<=-16'd17779;
      80663:data<=-16'd21193;
      80664:data<=-16'd15518;
      80665:data<=-16'd11126;
      80666:data<=-16'd8727;
      80667:data<=-16'd4704;
      80668:data<=-16'd5476;
      80669:data<=-16'd9004;
      80670:data<=-16'd4138;
      80671:data<=-16'd1380;
      80672:data<=-16'd4896;
      80673:data<=16'd197;
      80674:data<=16'd7256;
      80675:data<=16'd6032;
      80676:data<=16'd3418;
      80677:data<=16'd6598;
      80678:data<=16'd18551;
      80679:data<=16'd29016;
      80680:data<=16'd30590;
      80681:data<=16'd29157;
      80682:data<=16'd22328;
      80683:data<=16'd17362;
      80684:data<=16'd24216;
      80685:data<=16'd28765;
      80686:data<=16'd26900;
      80687:data<=16'd25147;
      80688:data<=16'd21808;
      80689:data<=16'd23099;
      80690:data<=16'd27943;
      80691:data<=16'd26729;
      80692:data<=16'd22559;
      80693:data<=16'd22668;
      80694:data<=16'd29540;
      80695:data<=16'd30949;
      80696:data<=16'd20086;
      80697:data<=16'd17576;
      80698:data<=16'd23044;
      80699:data<=16'd19012;
      80700:data<=16'd17353;
      80701:data<=16'd20281;
      80702:data<=16'd15672;
      80703:data<=16'd15396;
      80704:data<=16'd21406;
      80705:data<=16'd20648;
      80706:data<=16'd20598;
      80707:data<=16'd24683;
      80708:data<=16'd22174;
      80709:data<=16'd18682;
      80710:data<=16'd20281;
      80711:data<=16'd18804;
      80712:data<=16'd17687;
      80713:data<=16'd21006;
      80714:data<=16'd19176;
      80715:data<=16'd14613;
      80716:data<=16'd14747;
      80717:data<=16'd16633;
      80718:data<=16'd17561;
      80719:data<=16'd13135;
      80720:data<=16'd5025;
      80721:data<=-16'd1069;
      80722:data<=-16'd6699;
      80723:data<=-16'd4664;
      80724:data<=16'd1811;
      80725:data<=-16'd1915;
      80726:data<=-16'd1362;
      80727:data<=16'd7101;
      80728:data<=16'd4152;
      80729:data<=-16'd1163;
      80730:data<=-16'd2855;
      80731:data<=-16'd7941;
      80732:data<=-16'd6310;
      80733:data<=-16'd2179;
      80734:data<=-16'd5453;
      80735:data<=-16'd6320;
      80736:data<=-16'd4807;
      80737:data<=-16'd8379;
      80738:data<=-16'd11250;
      80739:data<=-16'd6115;
      80740:data<=-16'd1359;
      80741:data<=-16'd5256;
      80742:data<=-16'd4513;
      80743:data<=16'd523;
      80744:data<=-16'd2447;
      80745:data<=16'd702;
      80746:data<=16'd6182;
      80747:data<=-16'd3257;
      80748:data<=-16'd9192;
      80749:data<=-16'd7009;
      80750:data<=-16'd8334;
      80751:data<=-16'd3479;
      80752:data<=16'd2020;
      80753:data<=-16'd1668;
      80754:data<=-16'd1648;
      80755:data<=16'd3265;
      80756:data<=16'd1483;
      80757:data<=-16'd2672;
      80758:data<=16'd3313;
      80759:data<=16'd9799;
      80760:data<=16'd5573;
      80761:data<=16'd9318;
      80762:data<=16'd19996;
      80763:data<=16'd19120;
      80764:data<=16'd19701;
      80765:data<=16'd21211;
      80766:data<=16'd15430;
      80767:data<=16'd18812;
      80768:data<=16'd20498;
      80769:data<=16'd10675;
      80770:data<=16'd10144;
      80771:data<=16'd14891;
      80772:data<=16'd14384;
      80773:data<=16'd11869;
      80774:data<=16'd9036;
      80775:data<=16'd12557;
      80776:data<=16'd11376;
      80777:data<=16'd2878;
      80778:data<=16'd11041;
      80779:data<=16'd18965;
      80780:data<=16'd7218;
      80781:data<=16'd5231;
      80782:data<=16'd15518;
      80783:data<=16'd14371;
      80784:data<=16'd7423;
      80785:data<=16'd6109;
      80786:data<=16'd10287;
      80787:data<=16'd13147;
      80788:data<=16'd6639;
      80789:data<=-16'd1024;
      80790:data<=-16'd431;
      80791:data<=-16'd118;
      80792:data<=-16'd837;
      80793:data<=16'd5497;
      80794:data<=16'd6208;
      80795:data<=-16'd3112;
      80796:data<=-16'd2130;
      80797:data<=16'd3865;
      80798:data<=-16'd85;
      80799:data<=-16'd4131;
      80800:data<=-16'd7003;
      80801:data<=-16'd7186;
      80802:data<=-16'd634;
      80803:data<=-16'd5821;
      80804:data<=-16'd18813;
      80805:data<=-16'd20997;
      80806:data<=-16'd21663;
      80807:data<=-16'd20938;
      80808:data<=-16'd17001;
      80809:data<=-16'd21076;
      80810:data<=-16'd23951;
      80811:data<=-16'd20830;
      80812:data<=-16'd19558;
      80813:data<=-16'd17179;
      80814:data<=-16'd16768;
      80815:data<=-16'd19535;
      80816:data<=-16'd20136;
      80817:data<=-16'd20067;
      80818:data<=-16'd17020;
      80819:data<=-16'd15590;
      80820:data<=-16'd20776;
      80821:data<=-16'd19708;
      80822:data<=-16'd14505;
      80823:data<=-16'd17790;
      80824:data<=-16'd19312;
      80825:data<=-16'd12982;
      80826:data<=-16'd12627;
      80827:data<=-16'd18939;
      80828:data<=-16'd19776;
      80829:data<=-16'd20039;
      80830:data<=-16'd24353;
      80831:data<=-16'd23975;
      80832:data<=-16'd23695;
      80833:data<=-16'd23905;
      80834:data<=-16'd18703;
      80835:data<=-16'd21566;
      80836:data<=-16'd24598;
      80837:data<=-16'd16192;
      80838:data<=-16'd17364;
      80839:data<=-16'd20868;
      80840:data<=-16'd16258;
      80841:data<=-16'd21282;
      80842:data<=-16'd21086;
      80843:data<=-16'd11717;
      80844:data<=-16'd14058;
      80845:data<=-16'd10408;
      80846:data<=16'd1277;
      80847:data<=16'd1069;
      80848:data<=16'd2491;
      80849:data<=16'd7150;
      80850:data<=16'd2546;
      80851:data<=16'd26;
      80852:data<=16'd3024;
      80853:data<=-16'd132;
      80854:data<=-16'd4276;
      80855:data<=16'd1318;
      80856:data<=16'd2267;
      80857:data<=-16'd7040;
      80858:data<=-16'd3991;
      80859:data<=16'd2902;
      80860:data<=-16'd2573;
      80861:data<=-16'd2828;
      80862:data<=-16'd1051;
      80863:data<=-16'd3753;
      80864:data<=16'd246;
      80865:data<=16'd1124;
      80866:data<=-16'd402;
      80867:data<=-16'd549;
      80868:data<=-16'd7841;
      80869:data<=-16'd4385;
      80870:data<=16'd5441;
      80871:data<=16'd745;
      80872:data<=16'd152;
      80873:data<=16'd4308;
      80874:data<=16'd2678;
      80875:data<=16'd5495;
      80876:data<=16'd3873;
      80877:data<=-16'd693;
      80878:data<=16'd5357;
      80879:data<=16'd13091;
      80880:data<=16'd18392;
      80881:data<=16'd17620;
      80882:data<=16'd12953;
      80883:data<=16'd17051;
      80884:data<=16'd18125;
      80885:data<=16'd15036;
      80886:data<=16'd18951;
      80887:data<=16'd12461;
      80888:data<=-16'd3428;
      80889:data<=-16'd7028;
      80890:data<=-16'd2121;
      80891:data<=-16'd1225;
      80892:data<=-16'd5251;
      80893:data<=-16'd4420;
      80894:data<=16'd1145;
      80895:data<=16'd1119;
      80896:data<=16'd1929;
      80897:data<=16'd4276;
      80898:data<=16'd159;
      80899:data<=-16'd4778;
      80900:data<=-16'd8331;
      80901:data<=-16'd5844;
      80902:data<=16'd1952;
      80903:data<=16'd961;
      80904:data<=-16'd89;
      80905:data<=16'd3785;
      80906:data<=16'd1251;
      80907:data<=16'd1058;
      80908:data<=16'd3469;
      80909:data<=16'd3007;
      80910:data<=16'd9104;
      80911:data<=16'd13599;
      80912:data<=16'd8904;
      80913:data<=16'd4046;
      80914:data<=16'd2455;
      80915:data<=16'd4846;
      80916:data<=16'd6523;
      80917:data<=16'd7739;
      80918:data<=16'd11670;
      80919:data<=16'd7192;
      80920:data<=16'd1177;
      80921:data<=16'd5512;
      80922:data<=16'd8523;
      80923:data<=16'd10446;
      80924:data<=16'd12182;
      80925:data<=16'd7009;
      80926:data<=16'd6319;
      80927:data<=16'd10249;
      80928:data<=16'd9218;
      80929:data<=16'd8611;
      80930:data<=16'd9834;
      80931:data<=16'd12029;
      80932:data<=16'd15459;
      80933:data<=16'd17931;
      80934:data<=16'd20729;
      80935:data<=16'd19843;
      80936:data<=16'd16208;
      80937:data<=16'd16207;
      80938:data<=16'd15321;
      80939:data<=16'd14043;
      80940:data<=16'd13835;
      80941:data<=16'd10810;
      80942:data<=16'd12091;
      80943:data<=16'd18201;
      80944:data<=16'd20835;
      80945:data<=16'd20450;
      80946:data<=16'd16051;
      80947:data<=16'd10919;
      80948:data<=16'd13471;
      80949:data<=16'd16079;
      80950:data<=16'd10765;
      80951:data<=16'd9288;
      80952:data<=16'd14492;
      80953:data<=16'd11086;
      80954:data<=16'd6137;
      80955:data<=16'd11906;
      80956:data<=16'd12516;
      80957:data<=16'd11341;
      80958:data<=16'd18307;
      80959:data<=16'd13279;
      80960:data<=16'd6050;
      80961:data<=16'd12279;
      80962:data<=16'd9392;
      80963:data<=16'd3591;
      80964:data<=16'd8668;
      80965:data<=16'd8439;
      80966:data<=16'd6974;
      80967:data<=16'd9702;
      80968:data<=16'd7488;
      80969:data<=16'd4511;
      80970:data<=16'd3357;
      80971:data<=16'd2373;
      80972:data<=-16'd2834;
      80973:data<=-16'd13392;
      80974:data<=-16'd15417;
      80975:data<=-16'd10751;
      80976:data<=-16'd10608;
      80977:data<=-16'd14832;
      80978:data<=-16'd21673;
      80979:data<=-16'd17132;
      80980:data<=-16'd5506;
      80981:data<=-16'd7197;
      80982:data<=-16'd6052;
      80983:data<=-16'd3;
      80984:data<=-16'd6717;
      80985:data<=-16'd9821;
      80986:data<=-16'd8113;
      80987:data<=-16'd12777;
      80988:data<=-16'd12248;
      80989:data<=-16'd8596;
      80990:data<=-16'd6505;
      80991:data<=-16'd5841;
      80992:data<=-16'd9852;
      80993:data<=-16'd8661;
      80994:data<=-16'd6185;
      80995:data<=-16'd8904;
      80996:data<=-16'd8267;
      80997:data<=-16'd11113;
      80998:data<=-16'd11864;
      80999:data<=-16'd4234;
      81000:data<=-16'd8034;
      81001:data<=-16'd14421;
      81002:data<=-16'd13113;
      81003:data<=-16'd16349;
      81004:data<=-16'd13530;
      81005:data<=-16'd9151;
      81006:data<=-16'd15150;
      81007:data<=-16'd13177;
      81008:data<=-16'd8188;
      81009:data<=-16'd10699;
      81010:data<=-16'd8294;
      81011:data<=-16'd6834;
      81012:data<=-16'd8335;
      81013:data<=-16'd4067;
      81014:data<=-16'd2484;
      81015:data<=-16'd3410;
      81016:data<=16'd763;
      81017:data<=16'd5456;
      81018:data<=16'd7909;
      81019:data<=16'd7785;
      81020:data<=16'd3410;
      81021:data<=-16'd1066;
      81022:data<=-16'd610;
      81023:data<=-16'd206;
      81024:data<=-16'd3809;
      81025:data<=-16'd3697;
      81026:data<=-16'd613;
      81027:data<=16'd802;
      81028:data<=16'd3277;
      81029:data<=-16'd1691;
      81030:data<=-16'd12043;
      81031:data<=-16'd11649;
      81032:data<=-16'd8053;
      81033:data<=-16'd8739;
      81034:data<=-16'd9699;
      81035:data<=-16'd12643;
      81036:data<=-16'd10948;
      81037:data<=-16'd8486;
      81038:data<=-16'd13900;
      81039:data<=-16'd12175;
      81040:data<=-16'd5037;
      81041:data<=-16'd7553;
      81042:data<=-16'd11588;
      81043:data<=-16'd10405;
      81044:data<=-16'd5541;
      81045:data<=-16'd2458;
      81046:data<=-16'd8947;
      81047:data<=-16'd15033;
      81048:data<=-16'd12148;
      81049:data<=-16'd7906;
      81050:data<=-16'd7421;
      81051:data<=-16'd10372;
      81052:data<=-16'd10931;
      81053:data<=-16'd8041;
      81054:data<=-16'd8029;
      81055:data<=-16'd10411;
      81056:data<=-16'd17385;
      81057:data<=-16'd26329;
      81058:data<=-16'd25980;
      81059:data<=-16'd22685;
      81060:data<=-16'd23278;
      81061:data<=-16'd21678;
      81062:data<=-16'd19763;
      81063:data<=-16'd20343;
      81064:data<=-16'd19499;
      81065:data<=-16'd15224;
      81066:data<=-16'd14207;
      81067:data<=-16'd19012;
      81068:data<=-16'd16134;
      81069:data<=-16'd10875;
      81070:data<=-16'd15864;
      81071:data<=-16'd14034;
      81072:data<=-16'd6815;
      81073:data<=-16'd8834;
      81074:data<=-16'd8489;
      81075:data<=-16'd6905;
      81076:data<=-16'd5626;
      81077:data<=16'd802;
      81078:data<=-16'd3163;
      81079:data<=-16'd5600;
      81080:data<=16'd7232;
      81081:data<=16'd7714;
      81082:data<=16'd1381;
      81083:data<=16'd7242;
      81084:data<=16'd9362;
      81085:data<=16'd9462;
      81086:data<=16'd12185;
      81087:data<=16'd6724;
      81088:data<=16'd2990;
      81089:data<=16'd8251;
      81090:data<=16'd13603;
      81091:data<=16'd13785;
      81092:data<=16'd8769;
      81093:data<=16'd6561;
      81094:data<=16'd9400;
      81095:data<=16'd10425;
      81096:data<=16'd9380;
      81097:data<=16'd9894;
      81098:data<=16'd18882;
      81099:data<=16'd31076;
      81100:data<=16'd29625;
      81101:data<=16'd23619;
      81102:data<=16'd25511;
      81103:data<=16'd26562;
      81104:data<=16'd26786;
      81105:data<=16'd26920;
      81106:data<=16'd25135;
      81107:data<=16'd27558;
      81108:data<=16'd26166;
      81109:data<=16'd20609;
      81110:data<=16'd24635;
      81111:data<=16'd26356;
      81112:data<=16'd20941;
      81113:data<=16'd23096;
      81114:data<=16'd24565;
      81115:data<=16'd22092;
      81116:data<=16'd24964;
      81117:data<=16'd22870;
      81118:data<=16'd16874;
      81119:data<=16'd18901;
      81120:data<=16'd20633;
      81121:data<=16'd18468;
      81122:data<=16'd16543;
      81123:data<=16'd15117;
      81124:data<=16'd19158;
      81125:data<=16'd20545;
      81126:data<=16'd13041;
      81127:data<=16'd14404;
      81128:data<=16'd21828;
      81129:data<=16'd16207;
      81130:data<=16'd6578;
      81131:data<=16'd3987;
      81132:data<=16'd3873;
      81133:data<=16'd4855;
      81134:data<=16'd5836;
      81135:data<=16'd5800;
      81136:data<=16'd4746;
      81137:data<=16'd2608;
      81138:data<=16'd3562;
      81139:data<=16'd4202;
      81140:data<=-16'd1865;
      81141:data<=-16'd8837;
      81142:data<=-16'd11711;
      81143:data<=-16'd10837;
      81144:data<=-16'd7827;
      81145:data<=-16'd6067;
      81146:data<=-16'd5066;
      81147:data<=-16'd7163;
      81148:data<=-16'd11550;
      81149:data<=-16'd9212;
      81150:data<=-16'd5859;
      81151:data<=-16'd7116;
      81152:data<=-16'd5292;
      81153:data<=-16'd3917;
      81154:data<=-16'd4034;
      81155:data<=-16'd1929;
      81156:data<=-16'd3738;
      81157:data<=-16'd3228;
      81158:data<=16'd1629;
      81159:data<=-16'd746;
      81160:data<=-16'd3400;
      81161:data<=-16'd2367;
      81162:data<=-16'd3122;
      81163:data<=-16'd1600;
      81164:data<=-16'd1923;
      81165:data<=-16'd3767;
      81166:data<=-16'd3139;
      81167:data<=-16'd7194;
      81168:data<=-16'd6643;
      81169:data<=-16'd347;
      81170:data<=-16'd2720;
      81171:data<=-16'd2578;
      81172:data<=-16'd83;
      81173:data<=-16'd5071;
      81174:data<=-16'd3900;
      81175:data<=-16'd2372;
      81176:data<=-16'd5943;
      81177:data<=-16'd3899;
      81178:data<=-16'd7694;
      81179:data<=-16'd9253;
      81180:data<=16'd3454;
      81181:data<=16'd5648;
      81182:data<=16'd5110;
      81183:data<=16'd17841;
      81184:data<=16'd19519;
      81185:data<=16'd13121;
      81186:data<=16'd14716;
      81187:data<=16'd15250;
      81188:data<=16'd16362;
      81189:data<=16'd16020;
      81190:data<=16'd8314;
      81191:data<=16'd6714;
      81192:data<=16'd8862;
      81193:data<=16'd4491;
      81194:data<=16'd4111;
      81195:data<=16'd6922;
      81196:data<=16'd3263;
      81197:data<=16'd735;
      81198:data<=16'd2171;
      81199:data<=16'd1434;
      81200:data<=16'd94;
      81201:data<=-16'd3271;
      81202:data<=-16'd7891;
      81203:data<=-16'd4513;
      81204:data<=16'd1253;
      81205:data<=16'd373;
      81206:data<=-16'd902;
      81207:data<=-16'd1495;
      81208:data<=-16'd3048;
      81209:data<=-16'd2743;
      81210:data<=-16'd3183;
      81211:data<=-16'd2540;
      81212:data<=-16'd584;
      81213:data<=-16'd3169;
      81214:data<=-16'd6455;
      81215:data<=-16'd7850;
      81216:data<=-16'd7671;
      81217:data<=-16'd6551;
      81218:data<=-16'd9453;
      81219:data<=-16'd5802;
      81220:data<=16'd1481;
      81221:data<=-16'd10157;
      81222:data<=-16'd18950;
      81223:data<=-16'd9227;
      81224:data<=-16'd13435;
      81225:data<=-16'd27014;
      81226:data<=-16'd27065;
      81227:data<=-16'd23281;
      81228:data<=-16'd19429;
      81229:data<=-16'd21103;
      81230:data<=-16'd31492;
      81231:data<=-16'd34329;
      81232:data<=-16'd33909;
      81233:data<=-16'd35621;
      81234:data<=-16'd29666;
      81235:data<=-16'd26809;
      81236:data<=-16'd30876;
      81237:data<=-16'd29378;
      81238:data<=-16'd25372;
      81239:data<=-16'd24209;
      81240:data<=-16'd25561;
      81241:data<=-16'd26884;
      81242:data<=-16'd25689;
      81243:data<=-16'd24940;
      81244:data<=-16'd20495;
      81245:data<=-16'd14698;
      81246:data<=-16'd18060;
      81247:data<=-16'd20566;
      81248:data<=-16'd17791;
      81249:data<=-16'd19755;
      81250:data<=-16'd22266;
      81251:data<=-16'd22700;
      81252:data<=-16'd20776;
      81253:data<=-16'd13838;
      81254:data<=-16'd11371;
      81255:data<=-16'd13671;
      81256:data<=-16'd13038;
      81257:data<=-16'd12607;
      81258:data<=-16'd12675;
      81259:data<=-16'd12337;
      81260:data<=-16'd11726;
      81261:data<=-16'd10887;
      81262:data<=-16'd11953;
      81263:data<=-16'd8643;
      81264:data<=-16'd6237;
      81265:data<=-16'd13121;
      81266:data<=-16'd10188;
      81267:data<=16'd3159;
      81268:data<=16'd8936;
      81269:data<=16'd11468;
      81270:data<=16'd7799;
      81271:data<=16'd2702;
      81272:data<=16'd13670;
      81273:data<=16'd19532;
      81274:data<=16'd9385;
      81275:data<=16'd7655;
      81276:data<=16'd12813;
      81277:data<=16'd14411;
      81278:data<=16'd14659;
      81279:data<=16'd12113;
      81280:data<=16'd13647;
      81281:data<=16'd20724;
      81282:data<=16'd22030;
      81283:data<=16'd19062;
      81284:data<=16'd19229;
      81285:data<=16'd20030;
      81286:data<=16'd16650;
      81287:data<=16'd14035;
      81288:data<=16'd16791;
      81289:data<=16'd16791;
      81290:data<=16'd14910;
      81291:data<=16'd16992;
      81292:data<=16'd16248;
      81293:data<=16'd15951;
      81294:data<=16'd18830;
      81295:data<=16'd16716;
      81296:data<=16'd16349;
      81297:data<=16'd17992;
      81298:data<=16'd15007;
      81299:data<=16'd18218;
      81300:data<=16'd21616;
      81301:data<=16'd14339;
      81302:data<=16'd13057;
      81303:data<=16'd19555;
      81304:data<=16'd19085;
      81305:data<=16'd15038;
      81306:data<=16'd15183;
      81307:data<=16'd16842;
      81308:data<=16'd10096;
      81309:data<=-16'd1814;
      81310:data<=-16'd1142;
      81311:data<=16'd4473;
      81312:data<=-16'd569;
      81313:data<=-16'd3841;
      81314:data<=16'd926;
      81315:data<=16'd3979;
      81316:data<=16'd1727;
      81317:data<=-16'd4341;
      81318:data<=-16'd5049;
      81319:data<=16'd540;
      81320:data<=16'd737;
      81321:data<=16'd884;
      81322:data<=16'd6091;
      81323:data<=16'd6949;
      81324:data<=16'd6040;
      81325:data<=16'd6346;
      81326:data<=16'd4363;
      81327:data<=16'd4488;
      81328:data<=16'd5841;
      81329:data<=16'd6561;
      81330:data<=16'd6907;
      81331:data<=-16'd1386;
      81332:data<=-16'd8869;
      81333:data<=-16'd1959;
      81334:data<=-16'd494;
      81335:data<=-16'd10234;
      81336:data<=-16'd8934;
      81337:data<=-16'd3033;
      81338:data<=-16'd4300;
      81339:data<=-16'd1574;
      81340:data<=16'd1864;
      81341:data<=16'd1733;
      81342:data<=16'd3230;
      81343:data<=-16'd3149;
      81344:data<=-16'd9109;
      81345:data<=-16'd1039;
      81346:data<=16'd1657;
      81347:data<=-16'd297;
      81348:data<=16'd4548;
      81349:data<=16'd2099;
      81350:data<=16'd4681;
      81351:data<=16'd19406;
      81352:data<=16'd20812;
      81353:data<=16'd18369;
      81354:data<=16'd22248;
      81355:data<=16'd18422;
      81356:data<=16'd16777;
      81357:data<=16'd20033;
      81358:data<=16'd20174;
      81359:data<=16'd21217;
      81360:data<=16'd18854;
      81361:data<=16'd17925;
      81362:data<=16'd19146;
      81363:data<=16'd10035;
      81364:data<=16'd4444;
      81365:data<=16'd8170;
      81366:data<=16'd9803;
      81367:data<=16'd12974;
      81368:data<=16'd12760;
      81369:data<=16'd9177;
      81370:data<=16'd8621;
      81371:data<=16'd4839;
      81372:data<=16'd7567;
      81373:data<=16'd13712;
      81374:data<=16'd6379;
      81375:data<=16'd2088;
      81376:data<=16'd5820;
      81377:data<=16'd5189;
      81378:data<=16'd3589;
      81379:data<=-16'd1234;
      81380:data<=-16'd3668;
      81381:data<=16'd2990;
      81382:data<=16'd6601;
      81383:data<=16'd5838;
      81384:data<=16'd4528;
      81385:data<=16'd5109;
      81386:data<=16'd8587;
      81387:data<=16'd5890;
      81388:data<=16'd4384;
      81389:data<=16'd7635;
      81390:data<=16'd4404;
      81391:data<=16'd3636;
      81392:data<=16'd1334;
      81393:data<=-16'd12552;
      81394:data<=-16'd19103;
      81395:data<=-16'd17092;
      81396:data<=-16'd18387;
      81397:data<=-16'd18622;
      81398:data<=-16'd18070;
      81399:data<=-16'd19244;
      81400:data<=-16'd20428;
      81401:data<=-16'd17758;
      81402:data<=-16'd14856;
      81403:data<=-16'd18295;
      81404:data<=-16'd15770;
      81405:data<=-16'd10710;
      81406:data<=-16'd15158;
      81407:data<=-16'd14255;
      81408:data<=-16'd14090;
      81409:data<=-16'd19996;
      81410:data<=-16'd14528;
      81411:data<=-16'd13684;
      81412:data<=-16'd19191;
      81413:data<=-16'd11799;
      81414:data<=-16'd9779;
      81415:data<=-16'd15593;
      81416:data<=-16'd14504;
      81417:data<=-16'd13339;
      81418:data<=-16'd13180;
      81419:data<=-16'd14530;
      81420:data<=-16'd16390;
      81421:data<=-16'd15167;
      81422:data<=-16'd14731;
      81423:data<=-16'd9923;
      81424:data<=-16'd7591;
      81425:data<=-16'd13553;
      81426:data<=-16'd13844;
      81427:data<=-16'd14963;
      81428:data<=-16'd16754;
      81429:data<=-16'd14310;
      81430:data<=-16'd20918;
      81431:data<=-16'd19538;
      81432:data<=-16'd12780;
      81433:data<=-16'd24166;
      81434:data<=-16'd21200;
      81435:data<=-16'd1701;
      81436:data<=16'd597;
      81437:data<=-16'd1410;
      81438:data<=-16'd2256;
      81439:data<=-16'd3333;
      81440:data<=16'd3139;
      81441:data<=16'd2631;
      81442:data<=-16'd1959;
      81443:data<=-16'd2796;
      81444:data<=-16'd3876;
      81445:data<=16'd1295;
      81446:data<=16'd411;
      81447:data<=-16'd4184;
      81448:data<=16'd3700;
      81449:data<=16'd843;
      81450:data<=-16'd7808;
      81451:data<=-16'd519;
      81452:data<=16'd144;
      81453:data<=-16'd4757;
      81454:data<=-16'd2578;
      81455:data<=-16'd7210;
      81456:data<=-16'd10270;
      81457:data<=-16'd4596;
      81458:data<=-16'd2437;
      81459:data<=-16'd2652;
      81460:data<=-16'd4434;
      81461:data<=-16'd7122;
      81462:data<=-16'd2637;
      81463:data<=16'd3618;
      81464:data<=-16'd55;
      81465:data<=-16'd7645;
      81466:data<=-16'd5298;
      81467:data<=16'd165;
      81468:data<=-16'd1522;
      81469:data<=-16'd1334;
      81470:data<=16'd393;
      81471:data<=-16'd476;
      81472:data<=16'd4528;
      81473:data<=16'd8408;
      81474:data<=16'd4267;
      81475:data<=16'd722;
      81476:data<=-16'd4684;
      81477:data<=-16'd11256;
      81478:data<=-16'd10909;
      81479:data<=-16'd10170;
      81480:data<=-16'd10182;
      81481:data<=-16'd4106;
      81482:data<=-16'd343;
      81483:data<=-16'd3425;
      81484:data<=-16'd2693;
      81485:data<=16'd288;
      81486:data<=-16'd778;
      81487:data<=16'd3538;
      81488:data<=16'd10140;
      81489:data<=16'd6260;
      81490:data<=16'd2520;
      81491:data<=16'd4564;
      81492:data<=16'd4405;
      81493:data<=16'd5952;
      81494:data<=16'd6219;
      81495:data<=16'd4238;
      81496:data<=16'd8725;
      81497:data<=16'd8028;
      81498:data<=16'd2231;
      81499:data<=16'd6355;
      81500:data<=16'd8631;
      81501:data<=16'd6855;
      81502:data<=16'd9166;
      81503:data<=16'd7404;
      81504:data<=16'd10204;
      81505:data<=16'd16386;
      81506:data<=16'd9283;
      81507:data<=16'd6316;
      81508:data<=16'd10812;
      81509:data<=16'd5491;
      81510:data<=16'd4062;
      81511:data<=16'd7738;
      81512:data<=16'd6470;
      81513:data<=16'd10481;
      81514:data<=16'd13617;
      81515:data<=16'd12073;
      81516:data<=16'd14763;
      81517:data<=16'd12863;
      81518:data<=16'd10707;
      81519:data<=16'd17990;
      81520:data<=16'd23645;
      81521:data<=16'd26790;
      81522:data<=16'd28125;
      81523:data<=16'd25532;
      81524:data<=16'd27904;
      81525:data<=16'd28938;
      81526:data<=16'd23634;
      81527:data<=16'd23831;
      81528:data<=16'd25607;
      81529:data<=16'd21478;
      81530:data<=16'd16730;
      81531:data<=16'd15904;
      81532:data<=16'd17202;
      81533:data<=16'd11771;
      81534:data<=16'd5359;
      81535:data<=16'd10709;
      81536:data<=16'd15549;
      81537:data<=16'd14057;
      81538:data<=16'd16571;
      81539:data<=16'd18346;
      81540:data<=16'd17684;
      81541:data<=16'd19329;
      81542:data<=16'd18450;
      81543:data<=16'd16126;
      81544:data<=16'd15797;
      81545:data<=16'd15180;
      81546:data<=16'd15077;
      81547:data<=16'd15576;
      81548:data<=16'd15141;
      81549:data<=16'd13788;
      81550:data<=16'd12672;
      81551:data<=16'd12904;
      81552:data<=16'd12684;
      81553:data<=16'd12722;
      81554:data<=16'd13738;
      81555:data<=16'd13241;
      81556:data<=16'd13344;
      81557:data<=16'd12742;
      81558:data<=16'd10026;
      81559:data<=16'd11311;
      81560:data<=16'd9682;
      81561:data<=-16'd1571;
      81562:data<=-16'd8175;
      81563:data<=-16'd5441;
      81564:data<=-16'd4631;
      81565:data<=-16'd7961;
      81566:data<=-16'd9260;
      81567:data<=-16'd6802;
      81568:data<=-16'd7006;
      81569:data<=-16'd10178;
      81570:data<=-16'd9277;
      81571:data<=-16'd8179;
      81572:data<=-16'd9843;
      81573:data<=-16'd9420;
      81574:data<=-16'd9138;
      81575:data<=-16'd9321;
      81576:data<=-16'd8185;
      81577:data<=-16'd8795;
      81578:data<=-16'd9426;
      81579:data<=-16'd9982;
      81580:data<=-16'd10269;
      81581:data<=-16'd4915;
      81582:data<=-16'd191;
      81583:data<=-16'd1935;
      81584:data<=-16'd2820;
      81585:data<=-16'd2050;
      81586:data<=-16'd2977;
      81587:data<=-16'd4288;
      81588:data<=-16'd5066;
      81589:data<=-16'd4108;
      81590:data<=-16'd3879;
      81591:data<=-16'd6314;
      81592:data<=-16'd7683;
      81593:data<=-16'd8489;
      81594:data<=-16'd9991;
      81595:data<=-16'd10093;
      81596:data<=-16'd9477;
      81597:data<=-16'd9367;
      81598:data<=-16'd10410;
      81599:data<=-16'd10681;
      81600:data<=-16'd9104;
      81601:data<=-16'd9817;
      81602:data<=-16'd7993;
      81603:data<=16'd1257;
      81604:data<=16'd7103;
      81605:data<=16'd6255;
      81606:data<=16'd5470;
      81607:data<=16'd4350;
      81608:data<=16'd3603;
      81609:data<=16'd3770;
      81610:data<=16'd2109;
      81611:data<=16'd1054;
      81612:data<=16'd1384;
      81613:data<=16'd737;
      81614:data<=16'd508;
      81615:data<=16'd828;
      81616:data<=-16'd644;
      81617:data<=-16'd2764;
      81618:data<=-16'd3016;
      81619:data<=-16'd3316;
      81620:data<=-16'd4143;
      81621:data<=-16'd3243;
      81622:data<=-16'd4502;
      81623:data<=-16'd7215;
      81624:data<=-16'd5862;
      81625:data<=-16'd5571;
      81626:data<=-16'd6469;
      81627:data<=-16'd4861;
      81628:data<=-16'd7163;
      81629:data<=-16'd9132;
      81630:data<=-16'd7476;
      81631:data<=-16'd12058;
      81632:data<=-16'd16528;
      81633:data<=-16'd15302;
      81634:data<=-16'd17014;
      81635:data<=-16'd17587;
      81636:data<=-16'd14847;
      81637:data<=-16'd15033;
      81638:data<=-16'd15167;
      81639:data<=-16'd14578;
      81640:data<=-16'd14763;
      81641:data<=-16'd14750;
      81642:data<=-16'd15452;
      81643:data<=-16'd13399;
      81644:data<=-16'd12988;
      81645:data<=-16'd22633;
      81646:data<=-16'd31651;
      81647:data<=-16'd31490;
      81648:data<=-16'd29194;
      81649:data<=-16'd27881;
      81650:data<=-16'd27082;
      81651:data<=-16'd26500;
      81652:data<=-16'd25219;
      81653:data<=-16'd25314;
      81654:data<=-16'd26254;
      81655:data<=-16'd25396;
      81656:data<=-16'd23754;
      81657:data<=-16'd22861;
      81658:data<=-16'd22403;
      81659:data<=-16'd21444;
      81660:data<=-16'd20632;
      81661:data<=-16'd20626;
      81662:data<=-16'd19860;
      81663:data<=-16'd18359;
      81664:data<=-16'd17258;
      81665:data<=-16'd16604;
      81666:data<=-16'd16137;
      81667:data<=-16'd14998;
      81668:data<=-16'd14069;
      81669:data<=-16'd13480;
      81670:data<=-16'd12110;
      81671:data<=-16'd11768;
      81672:data<=-16'd10402;
      81673:data<=-16'd7122;
      81674:data<=-16'd7944;
      81675:data<=-16'd9515;
      81676:data<=-16'd7644;
      81677:data<=-16'd7363;
      81678:data<=-16'd6191;
      81679:data<=-16'd4225;
      81680:data<=-16'd5494;
      81681:data<=-16'd1577;
      81682:data<=16'd5524;
      81683:data<=16'd5677;
      81684:data<=16'd5183;
      81685:data<=16'd6382;
      81686:data<=16'd7964;
      81687:data<=16'd16624;
      81688:data<=16'd25073;
      81689:data<=16'd24512;
      81690:data<=16'd23212;
      81691:data<=16'd24586;
      81692:data<=16'd24450;
      81693:data<=16'd23065;
      81694:data<=16'd22268;
      81695:data<=16'd22196;
      81696:data<=16'd21362;
      81697:data<=16'd21341;
      81698:data<=16'd23074;
      81699:data<=16'd22406;
      81700:data<=16'd20347;
      81701:data<=16'd19323;
      81702:data<=16'd18045;
      81703:data<=16'd18460;
      81704:data<=16'd19253;
      81705:data<=16'd18524;
      81706:data<=16'd18776;
      81707:data<=16'd16841;
      81708:data<=16'd13687;
      81709:data<=16'd15141;
      81710:data<=16'd16280;
      81711:data<=16'd14872;
      81712:data<=16'd15029;
      81713:data<=16'd14809;
      81714:data<=16'd14161;
      81715:data<=16'd14894;
      81716:data<=16'd15377;
      81717:data<=16'd15277;
      81718:data<=16'd14804;
      81719:data<=16'd14495;
      81720:data<=16'd13925;
      81721:data<=16'd13126;
      81722:data<=16'd14854;
      81723:data<=16'd16178;
      81724:data<=16'd14872;
      81725:data<=16'd14069;
      81726:data<=16'd11838;
      81727:data<=16'd10836;
      81728:data<=16'd12624;
      81729:data<=16'd6611;
      81730:data<=-16'd3321;
      81731:data<=-16'd7181;
      81732:data<=-16'd11338;
      81733:data<=-16'd14310;
      81734:data<=-16'd11759;
      81735:data<=-16'd11157;
      81736:data<=-16'd11122;
      81737:data<=-16'd9461;
      81738:data<=-16'd10756;
      81739:data<=-16'd10568;
      81740:data<=-16'd7388;
      81741:data<=-16'd6628;
      81742:data<=-16'd6763;
      81743:data<=-16'd6187;
      81744:data<=-16'd6410;
      81745:data<=-16'd6560;
      81746:data<=-16'd5670;
      81747:data<=-16'd3873;
      81748:data<=-16'd2369;
      81749:data<=-16'd1683;
      81750:data<=-16'd1104;
      81751:data<=-16'd1360;
      81752:data<=-16'd2402;
      81753:data<=-16'd2406;
      81754:data<=-16'd887;
      81755:data<=16'd212;
      81756:data<=-16'd629;
      81757:data<=-16'd984;
      81758:data<=16'd218;
      81759:data<=16'd372;
      81760:data<=16'd156;
      81761:data<=16'd981;
      81762:data<=16'd1444;
      81763:data<=16'd782;
      81764:data<=-16'd108;
      81765:data<=16'd517;
      81766:data<=16'd828;
      81767:data<=-16'd171;
      81768:data<=16'd1240;
      81769:data<=16'd977;
      81770:data<=-16'd1648;
      81771:data<=16'd4620;
      81772:data<=16'd14216;
      81773:data<=16'd15021;
      81774:data<=16'd13634;
      81775:data<=16'd13496;
      81776:data<=16'd12013;
      81777:data<=16'd11916;
      81778:data<=16'd11024;
      81779:data<=16'd8311;
      81780:data<=16'd7835;
      81781:data<=16'd10568;
      81782:data<=16'd15053;
      81783:data<=16'd16566;
      81784:data<=16'd14486;
      81785:data<=16'd13160;
      81786:data<=16'd11364;
      81787:data<=16'd9843;
      81788:data<=16'd10158;
      81789:data<=16'd9435;
      81790:data<=16'd8834;
      81791:data<=16'd7322;
      81792:data<=16'd4250;
      81793:data<=16'd3968;
      81794:data<=16'd3562;
      81795:data<=16'd2910;
      81796:data<=16'd4423;
      81797:data<=16'd2463;
      81798:data<=16'd446;
      81799:data<=16'd1589;
      81800:data<=-16'd456;
      81801:data<=-16'd1662;
      81802:data<=16'd188;
      81803:data<=-16'd566;
      81804:data<=-16'd2344;
      81805:data<=-16'd3112;
      81806:data<=-16'd2235;
      81807:data<=-16'd1633;
      81808:data<=-16'd3245;
      81809:data<=-16'd2394;
      81810:data<=-16'd3310;
      81811:data<=-16'd6645;
      81812:data<=-16'd4097;
      81813:data<=-16'd8146;
      81814:data<=-16'd20992;
      81815:data<=-16'd23690;
      81816:data<=-16'd22504;
      81817:data<=-16'd24547;
      81818:data<=-16'd22152;
      81819:data<=-16'd21237;
      81820:data<=-16'd21690;
      81821:data<=-16'd19071;
      81822:data<=-16'd20363;
      81823:data<=-16'd22239;
      81824:data<=-16'd20492;
      81825:data<=-16'd20163;
      81826:data<=-16'd20127;
      81827:data<=-16'd19425;
      81828:data<=-16'd19382;
      81829:data<=-16'd18516;
      81830:data<=-16'd17655;
      81831:data<=-16'd19064;
      81832:data<=-16'd22453;
      81833:data<=-16'd23795;
      81834:data<=-16'd23241;
      81835:data<=-16'd24288;
      81836:data<=-16'd23209;
      81837:data<=-16'd20870;
      81838:data<=-16'd21347;
      81839:data<=-16'd20205;
      81840:data<=-16'd19258;
      81841:data<=-16'd20898;
      81842:data<=-16'd19917;
      81843:data<=-16'd18492;
      81844:data<=-16'd18280;
      81845:data<=-16'd17217;
      81846:data<=-16'd16715;
      81847:data<=-16'd16251;
      81848:data<=-16'd17262;
      81849:data<=-16'd17764;
      81850:data<=-16'd14727;
      81851:data<=-16'd14747;
      81852:data<=-16'd14783;
      81853:data<=-16'd12621;
      81854:data<=-16'd15955;
      81855:data<=-16'd11702;
      81856:data<=16'd3512;
      81857:data<=16'd7780;
      81858:data<=16'd5045;
      81859:data<=16'd6451;
      81860:data<=16'd5015;
      81861:data<=16'd3935;
      81862:data<=16'd5585;
      81863:data<=16'd4623;
      81864:data<=16'd3914;
      81865:data<=16'd3952;
      81866:data<=16'd4077;
      81867:data<=16'd6055;
      81868:data<=16'd6266;
      81869:data<=16'd4880;
      81870:data<=16'd4831;
      81871:data<=16'd4569;
      81872:data<=16'd5312;
      81873:data<=16'd7288;
      81874:data<=16'd6393;
      81875:data<=16'd4637;
      81876:data<=16'd5912;
      81877:data<=16'd6464;
      81878:data<=16'd5565;
      81879:data<=16'd6954;
      81880:data<=16'd7567;
      81881:data<=16'd8795;
      81882:data<=16'd15361;
      81883:data<=16'd18682;
      81884:data<=16'd16449;
      81885:data<=16'd17211;
      81886:data<=16'd18254;
      81887:data<=16'd17525;
      81888:data<=16'd17517;
      81889:data<=16'd15869;
      81890:data<=16'd15558;
      81891:data<=16'd17192;
      81892:data<=16'd16989;
      81893:data<=16'd17526;
      81894:data<=16'd17311;
      81895:data<=16'd16625;
      81896:data<=16'd18140;
      81897:data<=16'd12310;
      81898:data<=16'd652;
      81899:data<=-16'd2843;
      81900:data<=-16'd1145;
      81901:data<=-16'd1131;
      81902:data<=-16'd1227;
      81903:data<=-16'd564;
      81904:data<=16'd1547;
      81905:data<=16'd2899;
      81906:data<=16'd2252;
      81907:data<=16'd2171;
      81908:data<=16'd1130;
      81909:data<=16'd176;
      81910:data<=16'd2181;
      81911:data<=16'd3328;
      81912:data<=16'd3297;
      81913:data<=16'd4631;
      81914:data<=16'd4502;
      81915:data<=16'd3099;
      81916:data<=16'd4526;
      81917:data<=16'd7376;
      81918:data<=16'd7498;
      81919:data<=16'd6686;
      81920:data<=16'd7709;
      81921:data<=16'd7865;
      81922:data<=16'd7562;
      81923:data<=16'd8975;
      81924:data<=16'd8719;
      81925:data<=16'd7436;
      81926:data<=16'd8388;
      81927:data<=16'd9025;
      81928:data<=16'd8517;
      81929:data<=16'd8805;
      81930:data<=16'd9762;
      81931:data<=16'd8348;
      81932:data<=16'd2212;
      81933:data<=-16'd1936;
      81934:data<=-16'd403;
      81935:data<=16'd588;
      81936:data<=16'd1992;
      81937:data<=16'd3002;
      81938:data<=-16'd212;
      81939:data<=16'd4159;
      81940:data<=16'd16524;
      81941:data<=16'd20266;
      81942:data<=16'd18810;
      81943:data<=16'd19892;
      81944:data<=16'd18621;
      81945:data<=16'd16856;
      81946:data<=16'd16662;
      81947:data<=16'd16493;
      81948:data<=16'd17866;
      81949:data<=16'd18131;
      81950:data<=16'd16941;
      81951:data<=16'd16792;
      81952:data<=16'd15458;
      81953:data<=16'd14651;
      81954:data<=16'd15940;
      81955:data<=16'd15729;
      81956:data<=16'd14471;
      81957:data<=16'd13743;
      81958:data<=16'd13109;
      81959:data<=16'd12498;
      81960:data<=16'd12390;
      81961:data<=16'd13608;
      81962:data<=16'd13303;
      81963:data<=16'd11195;
      81964:data<=16'd11115;
      81965:data<=16'd10824;
      81966:data<=16'd10293;
      81967:data<=16'd11640;
      81968:data<=16'd10575;
      81969:data<=16'd8182;
      81970:data<=16'd7692;
      81971:data<=16'd7319;
      81972:data<=16'd7047;
      81973:data<=16'd5513;
      81974:data<=16'd3709;
      81975:data<=16'd3466;
      81976:data<=16'd1983;
      81977:data<=16'd2293;
      81978:data<=16'd3159;
      81979:data<=16'd364;
      81980:data<=16'd385;
      81981:data<=-16'd2300;
      81982:data<=-16'd11420;
      81983:data<=-16'd11436;
      81984:data<=-16'd7125;
      81985:data<=-16'd9884;
      81986:data<=-16'd11402;
      81987:data<=-16'd11785;
      81988:data<=-16'd13091;
      81989:data<=-16'd11201;
      81990:data<=-16'd10290;
      81991:data<=-16'd10971;
      81992:data<=-16'd11823;
      81993:data<=-16'd13532;
      81994:data<=-16'd12818;
      81995:data<=-16'd11822;
      81996:data<=-16'd11899;
      81997:data<=-16'd11197;
      81998:data<=-16'd12455;
      81999:data<=-16'd13279;
      82000:data<=-16'd12370;
      82001:data<=-16'd13104;
      82002:data<=-16'd12627;
      82003:data<=-16'd11186;
      82004:data<=-16'd11900;
      82005:data<=-16'd12806;
      82006:data<=-16'd12857;
      82007:data<=-16'd12560;
      82008:data<=-16'd12878;
      82009:data<=-16'd12881;
      82010:data<=-16'd12167;
      82011:data<=-16'd13512;
      82012:data<=-16'd14041;
      82013:data<=-16'd13470;
      82014:data<=-16'd14395;
      82015:data<=-16'd12320;
      82016:data<=-16'd11671;
      82017:data<=-16'd14979;
      82018:data<=-16'd13946;
      82019:data<=-16'd13438;
      82020:data<=-16'd14242;
      82021:data<=-16'd11611;
      82022:data<=-16'd13245;
      82023:data<=-16'd11030;
      82024:data<=16'd1206;
      82025:data<=16'd5964;
      82026:data<=16'd3724;
      82027:data<=16'd4256;
      82028:data<=16'd3883;
      82029:data<=16'd3160;
      82030:data<=16'd3243;
      82031:data<=16'd2598;
      82032:data<=-16'd1209;
      82033:data<=-16'd7950;
      82034:data<=-16'd8301;
      82035:data<=-16'd5953;
      82036:data<=-16'd9028;
      82037:data<=-16'd9400;
      82038:data<=-16'd8238;
      82039:data<=-16'd9485;
      82040:data<=-16'd8301;
      82041:data<=-16'd8922;
      82042:data<=-16'd10483;
      82043:data<=-16'd8874;
      82044:data<=-16'd8681;
      82045:data<=-16'd8322;
      82046:data<=-16'd8334;
      82047:data<=-16'd10235;
      82048:data<=-16'd9219;
      82049:data<=-16'd8743;
      82050:data<=-16'd9063;
      82051:data<=-16'd6789;
      82052:data<=-16'd6599;
      82053:data<=-16'd7131;
      82054:data<=-16'd7371;
      82055:data<=-16'd8751;
      82056:data<=-16'd7706;
      82057:data<=-16'd7585;
      82058:data<=-16'd7991;
      82059:data<=-16'd5891;
      82060:data<=-16'd6828;
      82061:data<=-16'd7500;
      82062:data<=-16'd6901;
      82063:data<=-16'd8355;
      82064:data<=-16'd5705;
      82065:data<=-16'd8460;
      82066:data<=-16'd21303;
      82067:data<=-16'd24654;
      82068:data<=-16'd21194;
      82069:data<=-16'd21919;
      82070:data<=-16'd19842;
      82071:data<=-16'd18516;
      82072:data<=-16'd20192;
      82073:data<=-16'd17243;
      82074:data<=-16'd14249;
      82075:data<=-16'd14487;
      82076:data<=-16'd13423;
      82077:data<=-16'd12187;
      82078:data<=-16'd11937;
      82079:data<=-16'd10099;
      82080:data<=-16'd7994;
      82081:data<=-16'd8153;
      82082:data<=-16'd5049;
      82083:data<=16'd2382;
      82084:data<=16'd4305;
      82085:data<=16'd3169;
      82086:data<=16'd5509;
      82087:data<=16'd5391;
      82088:data<=16'd4223;
      82089:data<=16'd5694;
      82090:data<=16'd5395;
      82091:data<=16'd5535;
      82092:data<=16'd7188;
      82093:data<=16'd6711;
      82094:data<=16'd6120;
      82095:data<=16'd6672;
      82096:data<=16'd7103;
      82097:data<=16'd6693;
      82098:data<=16'd6948;
      82099:data<=16'd8937;
      82100:data<=16'd8366;
      82101:data<=16'd7535;
      82102:data<=16'd9016;
      82103:data<=16'd7112;
      82104:data<=16'd7753;
      82105:data<=16'd11283;
      82106:data<=16'd7777;
      82107:data<=16'd10818;
      82108:data<=16'd23839;
      82109:data<=16'd26256;
      82110:data<=16'd23514;
      82111:data<=16'd26269;
      82112:data<=16'd25564;
      82113:data<=16'd23414;
      82114:data<=16'd24221;
      82115:data<=16'd22824;
      82116:data<=16'd21349;
      82117:data<=16'd22877;
      82118:data<=16'd23534;
      82119:data<=16'd21869;
      82120:data<=16'd21064;
      82121:data<=16'd21399;
      82122:data<=16'd20528;
      82123:data<=16'd19908;
      82124:data<=16'd19694;
      82125:data<=16'd18732;
      82126:data<=16'd19332;
      82127:data<=16'd19538;
      82128:data<=16'd17908;
      82129:data<=16'd18266;
      82130:data<=16'd19317;
      82131:data<=16'd18437;
      82132:data<=16'd15007;
      82133:data<=16'd9347;
      82134:data<=16'd6589;
      82135:data<=16'd7362;
      82136:data<=16'd8196;
      82137:data<=16'd9277;
      82138:data<=16'd8707;
      82139:data<=16'd7018;
      82140:data<=16'd6537;
      82141:data<=16'd5680;
      82142:data<=16'd6610;
      82143:data<=16'd8241;
      82144:data<=16'd7145;
      82145:data<=16'd7480;
      82146:data<=16'd7081;
      82147:data<=16'd4824;
      82148:data<=16'd7236;
      82149:data<=16'd5712;
      82150:data<=-16'd4864;
      82151:data<=-16'd10334;
      82152:data<=-16'd9693;
      82153:data<=-16'd10622;
      82154:data<=-16'd9238;
      82155:data<=-16'd6351;
      82156:data<=-16'd6842;
      82157:data<=-16'd7207;
      82158:data<=-16'd6117;
      82159:data<=-16'd6370;
      82160:data<=-16'd6200;
      82161:data<=-16'd4740;
      82162:data<=-16'd4146;
      82163:data<=-16'd3839;
      82164:data<=-16'd4109;
      82165:data<=-16'd5201;
      82166:data<=-16'd4361;
      82167:data<=-16'd3677;
      82168:data<=-16'd5125;
      82169:data<=-16'd5096;
      82170:data<=-16'd4757;
      82171:data<=-16'd5697;
      82172:data<=-16'd5485;
      82173:data<=-16'd5357;
      82174:data<=-16'd5824;
      82175:data<=-16'd6499;
      82176:data<=-16'd7859;
      82177:data<=-16'd7086;
      82178:data<=-16'd5952;
      82179:data<=-16'd7318;
      82180:data<=-16'd8273;
      82181:data<=-16'd9013;
      82182:data<=-16'd7068;
      82183:data<=-16'd647;
      82184:data<=16'd1595;
      82185:data<=16'd0;
      82186:data<=-16'd176;
      82187:data<=-16'd2079;
      82188:data<=-16'd1768;
      82189:data<=16'd120;
      82190:data<=-16'd3256;
      82191:data<=-16'd631;
      82192:data<=16'd10472;
      82193:data<=16'd14142;
      82194:data<=16'd12375;
      82195:data<=16'd12630;
      82196:data<=16'd11532;
      82197:data<=16'd10730;
      82198:data<=16'd10392;
      82199:data<=16'd8028;
      82200:data<=16'd6777;
      82201:data<=16'd6519;
      82202:data<=16'd6485;
      82203:data<=16'd7330;
      82204:data<=16'd5482;
      82205:data<=16'd2302;
      82206:data<=16'd2006;
      82207:data<=16'd2094;
      82208:data<=16'd1213;
      82209:data<=16'd1374;
      82210:data<=16'd1794;
      82211:data<=16'd617;
      82212:data<=-16'd1169;
      82213:data<=-16'd1377;
      82214:data<=-16'd1350;
      82215:data<=-16'd2187;
      82216:data<=-16'd2074;
      82217:data<=-16'd2561;
      82218:data<=-16'd4191;
      82219:data<=-16'd4334;
      82220:data<=-16'd4525;
      82221:data<=-16'd4825;
      82222:data<=-16'd3533;
      82223:data<=-16'd4188;
      82224:data<=-16'd6664;
      82225:data<=-16'd6883;
      82226:data<=-16'd6499;
      82227:data<=-16'd7106;
      82228:data<=-16'd6664;
      82229:data<=-16'd6217;
      82230:data<=-16'd7627;
      82231:data<=-16'd7738;
      82232:data<=-16'd7344;
      82233:data<=-16'd15158;
      82234:data<=-16'd28297;
      82235:data<=-16'd33663;
      82236:data<=-16'd32540;
      82237:data<=-16'd32163;
      82238:data<=-16'd31019;
      82239:data<=-16'd29179;
      82240:data<=-16'd28333;
      82241:data<=-16'd27602;
      82242:data<=-16'd27560;
      82243:data<=-16'd27871;
      82244:data<=-16'd27613;
      82245:data<=-16'd26680;
      82246:data<=-16'd24674;
      82247:data<=-16'd23340;
      82248:data<=-16'd23649;
      82249:data<=-16'd23708;
      82250:data<=-16'd22830;
      82251:data<=-16'd21758;
      82252:data<=-16'd21074;
      82253:data<=-16'd20313;
      82254:data<=-16'd19687;
      82255:data<=-16'd20257;
      82256:data<=-16'd20165;
      82257:data<=-16'd18651;
      82258:data<=-16'd17390;
      82259:data<=-16'd16001;
      82260:data<=-16'd15497;
      82261:data<=-16'd16220;
      82262:data<=-16'd15700;
      82263:data<=-16'd14525;
      82264:data<=-16'd13391;
      82265:data<=-16'd12528;
      82266:data<=-16'd12587;
      82267:data<=-16'd11156;
      82268:data<=-16'd9624;
      82269:data<=-16'd10120;
      82270:data<=-16'd9417;
      82271:data<=-16'd8774;
      82272:data<=-16'd8739;
      82273:data<=-16'd6519;
      82274:data<=-16'd5398;
      82275:data<=-16'd2538;
      82276:data<=16'd7413;
      82277:data<=16'd14986;
      82278:data<=16'd14694;
      82279:data<=16'd14390;
      82280:data<=16'd15890;
      82281:data<=16'd15688;
      82282:data<=16'd16477;
      82283:data<=16'd20956;
      82284:data<=16'd24069;
      82285:data<=16'd23250;
      82286:data<=16'd23487;
      82287:data<=16'd24228;
      82288:data<=16'd22745;
      82289:data<=16'd22639;
      82290:data<=16'd23132;
      82291:data<=16'd21704;
      82292:data<=16'd21384;
      82293:data<=16'd22115;
      82294:data<=16'd22116;
      82295:data<=16'd22190;
      82296:data<=16'd21949;
      82297:data<=16'd21076;
      82298:data<=16'd20328;
      82299:data<=16'd20595;
      82300:data<=16'd21202;
      82301:data<=16'd20310;
      82302:data<=16'd19343;
      82303:data<=16'd19041;
      82304:data<=16'd18506;
      82305:data<=16'd19308;
      82306:data<=16'd19587;
      82307:data<=16'd18119;
      82308:data<=16'd17973;
      82309:data<=16'd16847;
      82310:data<=16'd15109;
      82311:data<=16'd16953;
      82312:data<=16'd17729;
      82313:data<=16'd16433;
      82314:data<=16'd16780;
      82315:data<=16'd15638;
      82316:data<=16'd14844;
      82317:data<=16'd14654;
      82318:data<=16'd7078;
      82319:data<=-16'd1485;
      82320:data<=-16'd1870;
      82321:data<=-16'd1328;
      82322:data<=-16'd2488;
      82323:data<=-16'd1222;
      82324:data<=16'd115;
      82325:data<=16'd493;
      82326:data<=16'd949;
      82327:data<=16'd1157;
      82328:data<=16'd1601;
      82329:data<=16'd1124;
      82330:data<=16'd926;
      82331:data<=16'd3268;
      82332:data<=16'd3257;
      82333:data<=-16'd1199;
      82334:data<=-16'd4502;
      82335:data<=-16'd5057;
      82336:data<=-16'd4181;
      82337:data<=-16'd2259;
      82338:data<=-16'd1833;
      82339:data<=-16'd2543;
      82340:data<=-16'd2038;
      82341:data<=-16'd2164;
      82342:data<=-16'd2234;
      82343:data<=16'd89;
      82344:data<=16'd1028;
      82345:data<=-16'd297;
      82346:data<=-16'd158;
      82347:data<=16'd109;
      82348:data<=16'd11;
      82349:data<=16'd1495;
      82350:data<=16'd2285;
      82351:data<=16'd2059;
      82352:data<=16'd2234;
      82353:data<=16'd1638;
      82354:data<=16'd1712;
      82355:data<=16'd2890;
      82356:data<=16'd3400;
      82357:data<=16'd4055;
      82358:data<=16'd3421;
      82359:data<=16'd3562;
      82360:data<=16'd11248;
      82361:data<=16'd20336;
      82362:data<=16'd21688;
      82363:data<=16'd20400;
      82364:data<=16'd20359;
      82365:data<=16'd18856;
      82366:data<=16'd17170;
      82367:data<=16'd16618;
      82368:data<=16'd15911;
      82369:data<=16'd15082;
      82370:data<=16'd14910;
      82371:data<=16'd15104;
      82372:data<=16'd13809;
      82373:data<=16'd11514;
      82374:data<=16'd11191;
      82375:data<=16'd11395;
      82376:data<=16'd9838;
      82377:data<=16'd8857;
      82378:data<=16'd8957;
      82379:data<=16'd8311;
      82380:data<=16'd7347;
      82381:data<=16'd5929;
      82382:data<=16'd4854;
      82383:data<=16'd7127;
      82384:data<=16'd10472;
      82385:data<=16'd10437;
      82386:data<=16'd8822;
      82387:data<=16'd7800;
      82388:data<=16'd6634;
      82389:data<=16'd5905;
      82390:data<=16'd5294;
      82391:data<=16'd4416;
      82392:data<=16'd3970;
      82393:data<=16'd2275;
      82394:data<=16'd626;
      82395:data<=16'd1519;
      82396:data<=16'd1081;
      82397:data<=-16'd191;
      82398:data<=16'd845;
      82399:data<=-16'd743;
      82400:data<=-16'd2933;
      82401:data<=-16'd2208;
      82402:data<=-16'd8984;
      82403:data<=-16'd20095;
      82404:data<=-16'd20833;
      82405:data<=-16'd18715;
      82406:data<=-16'd21282;
      82407:data<=-16'd20315;
      82408:data<=-16'd18246;
      82409:data<=-16'd19520;
      82410:data<=-16'd18547;
      82411:data<=-16'd17047;
      82412:data<=-16'd18550;
      82413:data<=-16'd19146;
      82414:data<=-16'd18242;
      82415:data<=-16'd17834;
      82416:data<=-16'd17291;
      82417:data<=-16'd17068;
      82418:data<=-16'd18240;
      82419:data<=-16'd19199;
      82420:data<=-16'd18616;
      82421:data<=-16'd18196;
      82422:data<=-16'd17685;
      82423:data<=-16'd16307;
      82424:data<=-16'd17515;
      82425:data<=-16'd19626;
      82426:data<=-16'd17934;
      82427:data<=-16'd16463;
      82428:data<=-16'd16557;
      82429:data<=-16'd14913;
      82430:data<=-16'd15690;
      82431:data<=-16'd18016;
      82432:data<=-16'd15870;
      82433:data<=-16'd15603;
      82434:data<=-16'd20017;
      82435:data<=-16'd20072;
      82436:data<=-16'd18243;
      82437:data<=-16'd20398;
      82438:data<=-16'd20074;
      82439:data<=-16'd18133;
      82440:data<=-16'd19314;
      82441:data<=-16'd17370;
      82442:data<=-16'd15499;
      82443:data<=-16'd18252;
      82444:data<=-16'd12466;
      82445:data<=-16'd273;
      82446:data<=16'd2337;
      82447:data<=16'd1011;
      82448:data<=16'd2023;
      82449:data<=16'd92;
      82450:data<=-16'd1315;
      82451:data<=-16'd187;
      82452:data<=16'd39;
      82453:data<=16'd487;
      82454:data<=16'd582;
      82455:data<=-16'd287;
      82456:data<=-16'd787;
      82457:data<=-16'd1296;
      82458:data<=-16'd1052;
      82459:data<=-16'd511;
      82460:data<=-16'd164;
      82461:data<=16'd247;
      82462:data<=-16'd1550;
      82463:data<=-16'd2892;
      82464:data<=-16'd1116;
      82465:data<=-16'd356;
      82466:data<=-16'd393;
      82467:data<=-16'd52;
      82468:data<=-16'd779;
      82469:data<=-16'd408;
      82470:data<=16'd296;
      82471:data<=16'd217;
      82472:data<=16'd1136;
      82473:data<=16'd1202;
      82474:data<=16'd1495;
      82475:data<=16'd3294;
      82476:data<=16'd3011;
      82477:data<=16'd2388;
      82478:data<=16'd2930;
      82479:data<=16'd2551;
      82480:data<=16'd3570;
      82481:data<=16'd5297;
      82482:data<=16'd4839;
      82483:data<=16'd5718;
      82484:data<=16'd10481;
      82485:data<=16'd13389;
      82486:data<=16'd6848;
      82487:data<=-16'd3651;
      82488:data<=-16'd6081;
      82489:data<=-16'd3806;
      82490:data<=-16'd3950;
      82491:data<=-16'd3711;
      82492:data<=-16'd2922;
      82493:data<=-16'd2544;
      82494:data<=-16'd1146;
      82495:data<=-16'd403;
      82496:data<=-16'd182;
      82497:data<=16'd61;
      82498:data<=-16'd422;
      82499:data<=16'd743;
      82500:data<=16'd2441;
      82501:data<=16'd1851;
      82502:data<=16'd1556;
      82503:data<=16'd1882;
      82504:data<=16'd1196;
      82505:data<=16'd1762;
      82506:data<=16'd3072;
      82507:data<=16'd2698;
      82508:data<=16'd2964;
      82509:data<=16'd4035;
      82510:data<=16'd3096;
      82511:data<=16'd3216;
      82512:data<=16'd5683;
      82513:data<=16'd5882;
      82514:data<=16'd5109;
      82515:data<=16'd5645;
      82516:data<=16'd5187;
      82517:data<=16'd5595;
      82518:data<=16'd7791;
      82519:data<=16'd8810;
      82520:data<=16'd8824;
      82521:data<=16'd8293;
      82522:data<=16'd7984;
      82523:data<=16'd7905;
      82524:data<=16'd6928;
      82525:data<=16'd8413;
      82526:data<=16'd9245;
      82527:data<=16'd6141;
      82528:data<=16'd11634;
      82529:data<=16'd23886;
      82530:data<=16'd25995;
      82531:data<=16'd24103;
      82532:data<=16'd25749;
      82533:data<=16'd22521;
      82534:data<=16'd17150;
      82535:data<=16'd15597;
      82536:data<=16'd15238;
      82537:data<=16'd15908;
      82538:data<=16'd16063;
      82539:data<=16'd14598;
      82540:data<=16'd14175;
      82541:data<=16'd13605;
      82542:data<=16'd13063;
      82543:data<=16'd14178;
      82544:data<=16'd14184;
      82545:data<=16'd13308;
      82546:data<=16'd13426;
      82547:data<=16'd12707;
      82548:data<=16'd11553;
      82549:data<=16'd12026;
      82550:data<=16'd12777;
      82551:data<=16'd12201;
      82552:data<=16'd11652;
      82553:data<=16'd11515;
      82554:data<=16'd10223;
      82555:data<=16'd9715;
      82556:data<=16'd11558;
      82557:data<=16'd12082;
      82558:data<=16'd10402;
      82559:data<=16'd9216;
      82560:data<=16'd8616;
      82561:data<=16'd8114;
      82562:data<=16'd8140;
      82563:data<=16'd8310;
      82564:data<=16'd7471;
      82565:data<=16'd6710;
      82566:data<=16'd7558;
      82567:data<=16'd6516;
      82568:data<=16'd4945;
      82569:data<=16'd7045;
      82570:data<=16'd2540;
      82571:data<=-16'd10596;
      82572:data<=-16'd15296;
      82573:data<=-16'd12404;
      82574:data<=-16'd13353;
      82575:data<=-16'd14187;
      82576:data<=-16'd13543;
      82577:data<=-16'd14465;
      82578:data<=-16'd14292;
      82579:data<=-16'd13465;
      82580:data<=-16'd13248;
      82581:data<=-16'd13673;
      82582:data<=-16'd14926;
      82583:data<=-16'd13271;
      82584:data<=-16'd8987;
      82585:data<=-16'd6996;
      82586:data<=-16'd7401;
      82587:data<=-16'd8407;
      82588:data<=-16'd8994;
      82589:data<=-16'd8827;
      82590:data<=-16'd8887;
      82591:data<=-16'd8711;
      82592:data<=-16'd8346;
      82593:data<=-16'd9030;
      82594:data<=-16'd9785;
      82595:data<=-16'd9401;
      82596:data<=-16'd9185;
      82597:data<=-16'd9931;
      82598:data<=-16'd9612;
      82599:data<=-16'd9048;
      82600:data<=-16'd10352;
      82601:data<=-16'd10238;
      82602:data<=-16'd9330;
      82603:data<=-16'd10395;
      82604:data<=-16'd9295;
      82605:data<=-16'd8011;
      82606:data<=-16'd10061;
      82607:data<=-16'd10907;
      82608:data<=-16'd10948;
      82609:data<=-16'd9967;
      82610:data<=-16'd7852;
      82611:data<=-16'd9912;
      82612:data<=-16'd7054;
      82613:data<=16'd4704;
      82614:data<=16'd8721;
      82615:data<=16'd5888;
      82616:data<=16'd6534;
      82617:data<=16'd6253;
      82618:data<=16'd4910;
      82619:data<=16'd4487;
      82620:data<=16'd3248;
      82621:data<=16'd2814;
      82622:data<=16'd2003;
      82623:data<=16'd1416;
      82624:data<=16'd1742;
      82625:data<=-16'd681;
      82626:data<=-16'd1756;
      82627:data<=16'd102;
      82628:data<=-16'd385;
      82629:data<=-16'd444;
      82630:data<=-16'd14;
      82631:data<=-16'd2144;
      82632:data<=-16'd2106;
      82633:data<=-16'd1665;
      82634:data<=-16'd5976;
      82635:data<=-16'd9054;
      82636:data<=-16'd7767;
      82637:data<=-16'd8261;
      82638:data<=-16'd10436;
      82639:data<=-16'd9577;
      82640:data<=-16'd8736;
      82641:data<=-16'd9846;
      82642:data<=-16'd9206;
      82643:data<=-16'd8904;
      82644:data<=-16'd10066;
      82645:data<=-16'd9562;
      82646:data<=-16'd9621;
      82647:data<=-16'd9967;
      82648:data<=-16'd8830;
      82649:data<=-16'd9075;
      82650:data<=-16'd9618;
      82651:data<=-16'd10161;
      82652:data<=-16'd10009;
      82653:data<=-16'd6607;
      82654:data<=-16'd10255;
      82655:data<=-16'd23050;
      82656:data<=-16'd28335;
      82657:data<=-16'd25761;
      82658:data<=-16'd24879;
      82659:data<=-16'd24090;
      82660:data<=-16'd23355;
      82661:data<=-16'd23309;
      82662:data<=-16'd22706;
      82663:data<=-16'd22521;
      82664:data<=-16'd21353;
      82665:data<=-16'd20227;
      82666:data<=-16'd20133;
      82667:data<=-16'd18283;
      82668:data<=-16'd17179;
      82669:data<=-16'd17508;
      82670:data<=-16'd15954;
      82671:data<=-16'd14813;
      82672:data<=-16'd14552;
      82673:data<=-16'd13129;
      82674:data<=-16'd11626;
      82675:data<=-16'd9975;
      82676:data<=-16'd8648;
      82677:data<=-16'd8226;
      82678:data<=-16'd7547;
      82679:data<=-16'd6848;
      82680:data<=-16'd5413;
      82681:data<=-16'd3783;
      82682:data<=-16'd3974;
      82683:data<=-16'd2846;
      82684:data<=16'd1513;
      82685:data<=16'd4952;
      82686:data<=16'd5392;
      82687:data<=16'd5720;
      82688:data<=16'd7400;
      82689:data<=16'd7808;
      82690:data<=16'd7709;
      82691:data<=16'd8607;
      82692:data<=16'd7738;
      82693:data<=16'd8422;
      82694:data<=16'd10772;
      82695:data<=16'd8525;
      82696:data<=16'd11890;
      82697:data<=16'd24742;
      82698:data<=16'd29055;
      82699:data<=16'd25878;
      82700:data<=16'd27070;
      82701:data<=16'd27390;
      82702:data<=16'd25927;
      82703:data<=16'd25895;
      82704:data<=16'd24163;
      82705:data<=16'd22920;
      82706:data<=16'd23852;
      82707:data<=16'd24140;
      82708:data<=16'd23470;
      82709:data<=16'd22395;
      82710:data<=16'd21761;
      82711:data<=16'd21091;
      82712:data<=16'd20580;
      82713:data<=16'd21735;
      82714:data<=16'd21596;
      82715:data<=16'd20330;
      82716:data<=16'd20535;
      82717:data<=16'd19320;
      82718:data<=16'd18557;
      82719:data<=16'd20533;
      82720:data<=16'd20582;
      82721:data<=16'd19255;
      82722:data<=16'd18607;
      82723:data<=16'd17364;
      82724:data<=16'd17274;
      82725:data<=16'd18031;
      82726:data<=16'd17491;
      82727:data<=16'd16531;
      82728:data<=16'd15902;
      82729:data<=16'd15171;
      82730:data<=16'd13998;
      82731:data<=16'd14082;
      82732:data<=16'd15097;
      82733:data<=16'd13675;
      82734:data<=16'd11000;
      82735:data<=16'd7498;
      82736:data<=16'd4781;
      82737:data<=16'd7652;
      82738:data<=16'd5497;
      82739:data<=-16'd7125;
      82740:data<=-16'd12123;
      82741:data<=-16'd8868;
      82742:data<=-16'd10006;
      82743:data<=-16'd9615;
      82744:data<=-16'd6763;
      82745:data<=-16'd7612;
      82746:data<=-16'd7589;
      82747:data<=-16'd6529;
      82748:data<=-16'd7268;
      82749:data<=-16'd6818;
      82750:data<=-16'd5554;
      82751:data<=-16'd4996;
      82752:data<=-16'd4467;
      82753:data<=-16'd4043;
      82754:data<=-16'd3814;
      82755:data<=-16'd3961;
      82756:data<=-16'd3374;
      82757:data<=-16'd2006;
      82758:data<=-16'd2077;
      82759:data<=-16'd2564;
      82760:data<=-16'd2253;
      82761:data<=-16'd2215;
      82762:data<=-16'd1533;
      82763:data<=-16'd158;
      82764:data<=16'd126;
      82765:data<=-16'd403;
      82766:data<=-16'd394;
      82767:data<=16'd168;
      82768:data<=16'd102;
      82769:data<=-16'd408;
      82770:data<=-16'd405;
      82771:data<=-16'd294;
      82772:data<=-16'd70;
      82773:data<=-16'd42;
      82774:data<=-16'd552;
      82775:data<=-16'd855;
      82776:data<=-16'd1498;
      82777:data<=-16'd1394;
      82778:data<=-16'd869;
      82779:data<=-16'd2881;
      82780:data<=16'd55;
      82781:data<=16'd11194;
      82782:data<=16'd15227;
      82783:data<=16'd11035;
      82784:data<=16'd12795;
      82785:data<=16'd17264;
      82786:data<=16'd17250;
      82787:data<=16'd16026;
      82788:data<=16'd14322;
      82789:data<=16'd12646;
      82790:data<=16'd12483;
      82791:data<=16'd12199;
      82792:data<=16'd11586;
      82793:data<=16'd10252;
      82794:data<=16'd8267;
      82795:data<=16'd7770;
      82796:data<=16'd7696;
      82797:data<=16'd7004;
      82798:data<=16'd6645;
      82799:data<=16'd5671;
      82800:data<=16'd4182;
      82801:data<=16'd3576;
      82802:data<=16'd3571;
      82803:data<=16'd3099;
      82804:data<=16'd2299;
      82805:data<=16'd2305;
      82806:data<=16'd1700;
      82807:data<=-16'd149;
      82808:data<=-16'd496;
      82809:data<=-16'd415;
      82810:data<=-16'd1157;
      82811:data<=-16'd723;
      82812:data<=-16'd1089;
      82813:data<=-16'd3007;
      82814:data<=-16'd3565;
      82815:data<=-16'd3509;
      82816:data<=-16'd4099;
      82817:data<=-16'd4602;
      82818:data<=-16'd4811;
      82819:data<=-16'd5832;
      82820:data<=-16'd6986;
      82821:data<=-16'd5432;
      82822:data<=-16'd7984;
      82823:data<=-16'd19235;
      82824:data<=-16'd25109;
      82825:data<=-16'd23123;
      82826:data<=-16'd24175;
      82827:data<=-16'd23910;
      82828:data<=-16'd21896;
      82829:data<=-16'd22971;
      82830:data<=-16'd20970;
      82831:data<=-16'd19763;
      82832:data<=-16'd22471;
      82833:data<=-16'd20674;
      82834:data<=-16'd20732;
      82835:data<=-16'd25760;
      82836:data<=-16'd25162;
      82837:data<=-16'd23397;
      82838:data<=-16'd25464;
      82839:data<=-16'd24862;
      82840:data<=-16'd23393;
      82841:data<=-16'd23400;
      82842:data<=-16'd21497;
      82843:data<=-16'd20274;
      82844:data<=-16'd21547;
      82845:data<=-16'd21367;
      82846:data<=-16'd20142;
      82847:data<=-16'd20301;
      82848:data<=-16'd19237;
      82849:data<=-16'd17247;
      82850:data<=-16'd17810;
      82851:data<=-16'd18202;
      82852:data<=-16'd16792;
      82853:data<=-16'd16316;
      82854:data<=-16'd15415;
      82855:data<=-16'd13779;
      82856:data<=-16'd14143;
      82857:data<=-16'd15074;
      82858:data<=-16'd14222;
      82859:data<=-16'd13016;
      82860:data<=-16'd12907;
      82861:data<=-16'd11550;
      82862:data<=-16'd10308;
      82863:data<=-16'd13082;
      82864:data<=-16'd10580;
      82865:data<=16'd1553;
      82866:data<=16'd7811;
      82867:data<=16'd6176;
      82868:data<=16'd6722;
      82869:data<=16'd6664;
      82870:data<=16'd6084;
      82871:data<=16'd7480;
      82872:data<=16'd6699;
      82873:data<=16'd6194;
      82874:data<=16'd7507;
      82875:data<=16'd7700;
      82876:data<=16'd8520;
      82877:data<=16'd9063;
      82878:data<=16'd8657;
      82879:data<=16'd8957;
      82880:data<=16'd8360;
      82881:data<=16'd9068;
      82882:data<=16'd10848;
      82883:data<=16'd9843;
      82884:data<=16'd11421;
      82885:data<=16'd16123;
      82886:data<=16'd16525;
      82887:data<=16'd15702;
      82888:data<=16'd17432;
      82889:data<=16'd17749;
      82890:data<=16'd16641;
      82891:data<=16'd16167;
      82892:data<=16'd15197;
      82893:data<=16'd14304;
      82894:data<=16'd15458;
      82895:data<=16'd16665;
      82896:data<=16'd15565;
      82897:data<=16'd14572;
      82898:data<=16'd14398;
      82899:data<=16'd13335;
      82900:data<=16'd13308;
      82901:data<=16'd14522;
      82902:data<=16'd14352;
      82903:data<=16'd13000;
      82904:data<=16'd12308;
      82905:data<=16'd13324;
      82906:data<=16'd11361;
      82907:data<=16'd2138;
      82908:data<=-16'd5048;
      82909:data<=-16'd3817;
      82910:data<=-16'd2337;
      82911:data<=-16'd3237;
      82912:data<=-16'd2717;
      82913:data<=-16'd1880;
      82914:data<=-16'd1394;
      82915:data<=-16'd1010;
      82916:data<=-16'd1157;
      82917:data<=-16'd1178;
      82918:data<=-16'd966;
      82919:data<=16'd384;
      82920:data<=16'd1988;
      82921:data<=16'd1468;
      82922:data<=16'd1089;
      82923:data<=16'd1506;
      82924:data<=16'd949;
      82925:data<=16'd1841;
      82926:data<=16'd3620;
      82927:data<=16'd3283;
      82928:data<=16'd2701;
      82929:data<=16'd2928;
      82930:data<=16'd2805;
      82931:data<=16'd2934;
      82932:data<=16'd4040;
      82933:data<=16'd4605;
      82934:data<=16'd2388;
      82935:data<=-16'd652;
      82936:data<=-16'd1794;
      82937:data<=-16'd1949;
      82938:data<=-16'd540;
      82939:data<=16'd1441;
      82940:data<=16'd1048;
      82941:data<=16'd731;
      82942:data<=16'd1246;
      82943:data<=16'd346;
      82944:data<=16'd379;
      82945:data<=16'd2300;
      82946:data<=16'd2942;
      82947:data<=16'd1274;
      82948:data<=16'd2863;
      82949:data<=16'd12460;
      82950:data<=16'd20706;
      82951:data<=16'd19936;
      82952:data<=16'd18114;
      82953:data<=16'd18560;
      82954:data<=16'd18199;
      82955:data<=16'd18073;
      82956:data<=16'd17611;
      82957:data<=16'd17391;
      82958:data<=16'd17878;
      82959:data<=16'd16760;
      82960:data<=16'd16008;
      82961:data<=16'd15691;
      82962:data<=16'd14512;
      82963:data<=16'd15164;
      82964:data<=16'd15773;
      82965:data<=16'd14744;
      82966:data<=16'd14043;
      82967:data<=16'd12783;
      82968:data<=16'd12069;
      82969:data<=16'd12022;
      82970:data<=16'd10828;
      82971:data<=16'd10481;
      82972:data<=16'd10070;
      82973:data<=16'd8895;
      82974:data<=16'd9042;
      82975:data<=16'd8012;
      82976:data<=16'd5668;
      82977:data<=16'd4605;
      82978:data<=16'd4212;
      82979:data<=16'd4187;
      82980:data<=16'd3237;
      82981:data<=16'd1532;
      82982:data<=16'd578;
      82983:data<=-16'd638;
      82984:data<=16'd473;
      82985:data<=16'd4199;
      82986:data<=16'd5676;
      82987:data<=16'd4954;
      82988:data<=16'd3245;
      82989:data<=16'd2563;
      82990:data<=16'd1351;
      82991:data<=-16'd8105;
      82992:data<=-16'd17214;
      82993:data<=-16'd15661;
      82994:data<=-16'd15001;
      82995:data<=-16'd17948;
      82996:data<=-16'd16886;
      82997:data<=-16'd16357;
      82998:data<=-16'd17112;
      82999:data<=-16'd16120;
      83000:data<=-16'd16348;
      83001:data<=-16'd16407;
      83002:data<=-16'd14795;
      83003:data<=-16'd14243;
      83004:data<=-16'd14590;
      83005:data<=-16'd14292;
      83006:data<=-16'd13806;
      83007:data<=-16'd14284;
      83008:data<=-16'd14343;
      83009:data<=-16'd13280;
      83010:data<=-16'd13673;
      83011:data<=-16'd14167;
      83012:data<=-16'd13254;
      83013:data<=-16'd13687;
      83014:data<=-16'd14436;
      83015:data<=-16'd14038;
      83016:data<=-16'd13955;
      83017:data<=-16'd13758;
      83018:data<=-16'd13367;
      83019:data<=-16'd13188;
      83020:data<=-16'd13323;
      83021:data<=-16'd13887;
      83022:data<=-16'd13274;
      83023:data<=-16'd11929;
      83024:data<=-16'd11377;
      83025:data<=-16'd11549;
      83026:data<=-16'd12740;
      83027:data<=-16'd12928;
      83028:data<=-16'd11849;
      83029:data<=-16'd11570;
      83030:data<=-16'd10345;
      83031:data<=-16'd10733;
      83032:data<=-16'd12410;
      83033:data<=-16'd5674;
      83034:data<=16'd2635;
      83035:data<=-16'd76;
      83036:data<=-16'd4014;
      83037:data<=-16'd2792;
      83038:data<=-16'd3621;
      83039:data<=-16'd4983;
      83040:data<=-16'd4387;
      83041:data<=-16'd4617;
      83042:data<=-16'd4473;
      83043:data<=-16'd4109;
      83044:data<=-16'd5231;
      83045:data<=-16'd5914;
      83046:data<=-16'd5783;
      83047:data<=-16'd5809;
      83048:data<=-16'd5069;
      83049:data<=-16'd4070;
      83050:data<=-16'd4554;
      83051:data<=-16'd5961;
      83052:data<=-16'd6499;
      83053:data<=-16'd6132;
      83054:data<=-16'd5720;
      83055:data<=-16'd5100;
      83056:data<=-16'd4599;
      83057:data<=-16'd5236;
      83058:data<=-16'd6222;
      83059:data<=-16'd6181;
      83060:data<=-16'd5765;
      83061:data<=-16'd5668;
      83062:data<=-16'd5156;
      83063:data<=-16'd5019;
      83064:data<=-16'd6466;
      83065:data<=-16'd7514;
      83066:data<=-16'd7169;
      83067:data<=-16'd6801;
      83068:data<=-16'd5903;
      83069:data<=-16'd5084;
      83070:data<=-16'd5430;
      83071:data<=-16'd5476;
      83072:data<=-16'd5529;
      83073:data<=-16'd4554;
      83074:data<=-16'd3078;
      83075:data<=-16'd8504;
      83076:data<=-16'd16639;
      83077:data<=-16'd16590;
      83078:data<=-16'd14281;
      83079:data<=-16'd14674;
      83080:data<=-16'd13617;
      83081:data<=-16'd13027;
      83082:data<=-16'd11929;
      83083:data<=-16'd9283;
      83084:data<=-16'd8862;
      83085:data<=-16'd6131;
      83086:data<=-16'd1488;
      83087:data<=-16'd1671;
      83088:data<=-16'd1325;
      83089:data<=16'd1334;
      83090:data<=16'd967;
      83091:data<=16'd699;
      83092:data<=16'd1588;
      83093:data<=16'd1158;
      83094:data<=16'd1938;
      83095:data<=16'd3676;
      83096:data<=16'd3917;
      83097:data<=16'd4165;
      83098:data<=16'd4977;
      83099:data<=16'd4273;
      83100:data<=16'd3553;
      83101:data<=16'd5174;
      83102:data<=16'd6002;
      83103:data<=16'd5691;
      83104:data<=16'd6886;
      83105:data<=16'd6619;
      83106:data<=16'd5630;
      83107:data<=16'd7203;
      83108:data<=16'd8175;
      83109:data<=16'd8208;
      83110:data<=16'd8595;
      83111:data<=16'd8254;
      83112:data<=16'd8431;
      83113:data<=16'd9015;
      83114:data<=16'd10093;
      83115:data<=16'd10234;
      83116:data<=16'd8428;
      83117:data<=16'd13643;
      83118:data<=16'd23563;
      83119:data<=16'd24988;
      83120:data<=16'd23763;
      83121:data<=16'd25373;
      83122:data<=16'd24260;
      83123:data<=16'd23499;
      83124:data<=16'd23326;
      83125:data<=16'd21631;
      83126:data<=16'd22298;
      83127:data<=16'd22958;
      83128:data<=16'd22074;
      83129:data<=16'd21678;
      83130:data<=16'd20152;
      83131:data<=16'd19020;
      83132:data<=16'd19129;
      83133:data<=16'd19355;
      83134:data<=16'd19757;
      83135:data<=16'd16847;
      83136:data<=16'd11659;
      83137:data<=16'd9665;
      83138:data<=16'd10534;
      83139:data<=16'd11594;
      83140:data<=16'd11254;
      83141:data<=16'd10878;
      83142:data<=16'd11022;
      83143:data<=16'd9482;
      83144:data<=16'd9341;
      83145:data<=16'd10608;
      83146:data<=16'd9755;
      83147:data<=16'd9774;
      83148:data<=16'd9309;
      83149:data<=16'd7374;
      83150:data<=16'd8031;
      83151:data<=16'd8284;
      83152:data<=16'd8436;
      83153:data<=16'd9508;
      83154:data<=16'd7514;
      83155:data<=16'd6790;
      83156:data<=16'd7050;
      83157:data<=16'd6373;
      83158:data<=16'd9323;
      83159:data<=16'd5250;
      83160:data<=-16'd6549;
      83161:data<=-16'd8337;
      83162:data<=-16'd6067;
      83163:data<=-16'd7844;
      83164:data<=-16'd6296;
      83165:data<=-16'd5115;
      83166:data<=-16'd5968;
      83167:data<=-16'd5049;
      83168:data<=-16'd5470;
      83169:data<=-16'd6097;
      83170:data<=-16'd5856;
      83171:data<=-16'd5959;
      83172:data<=-16'd4993;
      83173:data<=-16'd4949;
      83174:data<=-16'd5463;
      83175:data<=-16'd5189;
      83176:data<=-16'd6496;
      83177:data<=-16'd7538;
      83178:data<=-16'd6946;
      83179:data<=-16'd6420;
      83180:data<=-16'd6349;
      83181:data<=-16'd6827;
      83182:data<=-16'd6672;
      83183:data<=-16'd7373;
      83184:data<=-16'd8748;
      83185:data<=-16'd5911;
      83186:data<=-16'd2053;
      83187:data<=-16'd1210;
      83188:data<=-16'd1447;
      83189:data<=-16'd2886;
      83190:data<=-16'd3124;
      83191:data<=-16'd2402;
      83192:data<=-16'd3435;
      83193:data<=-16'd2666;
      83194:data<=-16'd2475;
      83195:data<=-16'd4413;
      83196:data<=-16'd3788;
      83197:data<=-16'd4124;
      83198:data<=-16'd4273;
      83199:data<=-16'd2649;
      83200:data<=-16'd5190;
      83201:data<=-16'd2382;
      83202:data<=16'd8067;
      83203:data<=16'd10005;
      83204:data<=16'd7300;
      83205:data<=16'd8381;
      83206:data<=16'd7670;
      83207:data<=16'd6217;
      83208:data<=16'd5504;
      83209:data<=16'd4309;
      83210:data<=16'd4461;
      83211:data<=16'd4225;
      83212:data<=16'd3918;
      83213:data<=16'd4087;
      83214:data<=16'd2561;
      83215:data<=16'd1773;
      83216:data<=16'd1858;
      83217:data<=16'd1374;
      83218:data<=16'd1730;
      83219:data<=16'd870;
      83220:data<=-16'd1286;
      83221:data<=-16'd2187;
      83222:data<=-16'd2174;
      83223:data<=-16'd1535;
      83224:data<=-16'd1489;
      83225:data<=-16'd2103;
      83226:data<=-16'd2641;
      83227:data<=-16'd4102;
      83228:data<=-16'd4384;
      83229:data<=-16'd4266;
      83230:data<=-16'd5372;
      83231:data<=-16'd4404;
      83232:data<=-16'd4966;
      83233:data<=-16'd7620;
      83234:data<=-16'd6422;
      83235:data<=-16'd7403;
      83236:data<=-16'd11685;
      83237:data<=-16'd11919;
      83238:data<=-16'd11993;
      83239:data<=-16'd13524;
      83240:data<=-16'd14035;
      83241:data<=-16'd13594;
      83242:data<=-16'd10595;
      83243:data<=-16'd13628;
      83244:data<=-16'd24582;
      83245:data<=-16'd27959;
      83246:data<=-16'd25484;
      83247:data<=-16'd26335;
      83248:data<=-16'd25739;
      83249:data<=-16'd23816;
      83250:data<=-16'd22798;
      83251:data<=-16'd21857;
      83252:data<=-16'd22742;
      83253:data<=-16'd22814;
      83254:data<=-16'd21873;
      83255:data<=-16'd21952;
      83256:data<=-16'd20095;
      83257:data<=-16'd18648;
      83258:data<=-16'd19516;
      83259:data<=-16'd19147;
      83260:data<=-16'd18518;
      83261:data<=-16'd17734;
      83262:data<=-16'd15620;
      83263:data<=-16'd14816;
      83264:data<=-16'd15641;
      83265:data<=-16'd16095;
      83266:data<=-16'd15297;
      83267:data<=-16'd14211;
      83268:data<=-16'd13490;
      83269:data<=-16'd12261;
      83270:data<=-16'd11815;
      83271:data<=-16'd11277;
      83272:data<=-16'd9485;
      83273:data<=-16'd9641;
      83274:data<=-16'd9603;
      83275:data<=-16'd7609;
      83276:data<=-16'd6510;
      83277:data<=-16'd4739;
      83278:data<=-16'd3953;
      83279:data<=-16'd4243;
      83280:data<=-16'd2032;
      83281:data<=-16'd1829;
      83282:data<=-16'd892;
      83283:data<=16'd1983;
      83284:data<=-16'd1202;
      83285:data<=16'd3585;
      83286:data<=16'd20198;
      83287:data<=16'd24230;
      83288:data<=16'd20551;
      83289:data<=16'd23798;
      83290:data<=16'd24263;
      83291:data<=16'd22486;
      83292:data<=16'd22991;
      83293:data<=16'd21322;
      83294:data<=16'd20673;
      83295:data<=16'd22046;
      83296:data<=16'd22306;
      83297:data<=16'd21931;
      83298:data<=16'd20939;
      83299:data<=16'd20293;
      83300:data<=16'd19567;
      83301:data<=16'd19205;
      83302:data<=16'd20657;
      83303:data<=16'd20027;
      83304:data<=16'd18325;
      83305:data<=16'd18694;
      83306:data<=16'd17998;
      83307:data<=16'd17579;
      83308:data<=16'd18537;
      83309:data<=16'd18204;
      83310:data<=16'd17860;
      83311:data<=16'd17376;
      83312:data<=16'd16436;
      83313:data<=16'd16083;
      83314:data<=16'd15891;
      83315:data<=16'd16771;
      83316:data<=16'd16642;
      83317:data<=16'd14836;
      83318:data<=16'd14301;
      83319:data<=16'd13570;
      83320:data<=16'd14088;
      83321:data<=16'd15576;
      83322:data<=16'd13967;
      83323:data<=16'd13784;
      83324:data<=16'd13477;
      83325:data<=16'd11176;
      83326:data<=16'd14122;
      83327:data<=16'd11982;
      83328:data<=16'd429;
      83329:data<=-16'd2961;
      83330:data<=-16'd1201;
      83331:data<=-16'd3045;
      83332:data<=-16'd2027;
      83333:data<=-16'd65;
      83334:data<=16'd130;
      83335:data<=-16'd1190;
      83336:data<=-16'd5717;
      83337:data<=-16'd7624;
      83338:data<=-16'd6255;
      83339:data<=-16'd5571;
      83340:data<=-16'd4314;
      83341:data<=-16'd4346;
      83342:data<=-16'd4360;
      83343:data<=-16'd3218;
      83344:data<=-16'd4570;
      83345:data<=-16'd4020;
      83346:data<=-16'd1099;
      83347:data<=-16'd1111;
      83348:data<=-16'd1206;
      83349:data<=-16'd1343;
      83350:data<=-16'd2463;
      83351:data<=-16'd1284;
      83352:data<=16'd320;
      83353:data<=16'd805;
      83354:data<=16'd654;
      83355:data<=16'd99;
      83356:data<=16'd619;
      83357:data<=16'd975;
      83358:data<=16'd1829;
      83359:data<=16'd3298;
      83360:data<=16'd2582;
      83361:data<=16'd2359;
      83362:data<=16'd2255;
      83363:data<=16'd1284;
      83364:data<=16'd3210;
      83365:data<=16'd3926;
      83366:data<=16'd3445;
      83367:data<=16'd4504;
      83368:data<=16'd1861;
      83369:data<=16'd4601;
      83370:data<=16'd16017;
      83371:data<=16'd18486;
      83372:data<=16'd15232;
      83373:data<=16'd16369;
      83374:data<=16'd15488;
      83375:data<=16'd14478;
      83376:data<=16'd14798;
      83377:data<=16'd12196;
      83378:data<=16'd10810;
      83379:data<=16'd10942;
      83380:data<=16'd10313;
      83381:data<=16'd9932;
      83382:data<=16'd8619;
      83383:data<=16'd7473;
      83384:data<=16'd6643;
      83385:data<=16'd6652;
      83386:data<=16'd9982;
      83387:data<=16'd11630;
      83388:data<=16'd9840;
      83389:data<=16'd8789;
      83390:data<=16'd7673;
      83391:data<=16'd7172;
      83392:data<=16'd6925;
      83393:data<=16'd5203;
      83394:data<=16'd5181;
      83395:data<=16'd4996;
      83396:data<=16'd2977;
      83397:data<=16'd2491;
      83398:data<=16'd1824;
      83399:data<=16'd1165;
      83400:data<=16'd1867;
      83401:data<=16'd851;
      83402:data<=-16'd863;
      83403:data<=-16'd1569;
      83404:data<=-16'd1666;
      83405:data<=-16'd1651;
      83406:data<=-16'd2534;
      83407:data<=-16'd2591;
      83408:data<=-16'd3952;
      83409:data<=-16'd6035;
      83410:data<=-16'd3078;
      83411:data<=-16'd5658;
      83412:data<=-16'd17064;
      83413:data<=-16'd20119;
      83414:data<=-16'd18619;
      83415:data<=-16'd21537;
      83416:data<=-16'd20588;
      83417:data<=-16'd18807;
      83418:data<=-16'd19669;
      83419:data<=-16'd18175;
      83420:data<=-16'd18622;
      83421:data<=-16'd20953;
      83422:data<=-16'd20635;
      83423:data<=-16'd19738;
      83424:data<=-16'd18456;
      83425:data<=-16'd17690;
      83426:data<=-16'd18466;
      83427:data<=-16'd18932;
      83428:data<=-16'd19258;
      83429:data<=-16'd18436;
      83430:data<=-16'd17209;
      83431:data<=-16'd17012;
      83432:data<=-16'd16352;
      83433:data<=-16'd17506;
      83434:data<=-16'd18460;
      83435:data<=-16'd16689;
      83436:data<=-16'd19023;
      83437:data<=-16'd22269;
      83438:data<=-16'd20424;
      83439:data<=-16'd20306;
      83440:data<=-16'd21732;
      83441:data<=-16'd20767;
      83442:data<=-16'd20204;
      83443:data<=-16'd18835;
      83444:data<=-16'd16869;
      83445:data<=-16'd17634;
      83446:data<=-16'd19083;
      83447:data<=-16'd18533;
      83448:data<=-16'd17004;
      83449:data<=-16'd16258;
      83450:data<=-16'd14730;
      83451:data<=-16'd14069;
      83452:data<=-16'd17438;
      83453:data<=-16'd14495;
      83454:data<=-16'd2802;
      83455:data<=16'd1753;
      83456:data<=16'd141;
      83457:data<=16'd1184;
      83458:data<=16'd164;
      83459:data<=-16'd1575;
      83460:data<=-16'd981;
      83461:data<=-16'd1275;
      83462:data<=-16'd767;
      83463:data<=16'd171;
      83464:data<=-16'd425;
      83465:data<=-16'd980;
      83466:data<=-16'd1929;
      83467:data<=-16'd2000;
      83468:data<=-16'd893;
      83469:data<=-16'd1201;
      83470:data<=-16'd1280;
      83471:data<=-16'd578;
      83472:data<=-16'd546;
      83473:data<=-16'd400;
      83474:data<=-16'd61;
      83475:data<=16'd482;
      83476:data<=16'd811;
      83477:data<=16'd1468;
      83478:data<=16'd3058;
      83479:data<=16'd2839;
      83480:data<=16'd2416;
      83481:data<=16'd3169;
      83482:data<=16'd2347;
      83483:data<=16'd3785;
      83484:data<=16'd6241;
      83485:data<=16'd4858;
      83486:data<=16'd6860;
      83487:data<=16'd11433;
      83488:data<=16'd11059;
      83489:data<=16'd10592;
      83490:data<=16'd11890;
      83491:data<=16'd12123;
      83492:data<=16'd11658;
      83493:data<=16'd10818;
      83494:data<=16'd11985;
      83495:data<=16'd9818;
      83496:data<=16'd825;
      83497:data<=-16'd2896;
      83498:data<=-16'd1166;
      83499:data<=-16'd2315;
      83500:data<=-16'd2197;
      83501:data<=-16'd1002;
      83502:data<=-16'd552;
      83503:data<=16'd1424;
      83504:data<=16'd1027;
      83505:data<=-16'd358;
      83506:data<=16'd422;
      83507:data<=16'd290;
      83508:data<=16'd1204;
      83509:data<=16'd3019;
      83510:data<=16'd2684;
      83511:data<=16'd2807;
      83512:data<=16'd2960;
      83513:data<=16'd2387;
      83514:data<=16'd3624;
      83515:data<=16'd5207;
      83516:data<=16'd5133;
      83517:data<=16'd4068;
      83518:data<=16'd3791;
      83519:data<=16'd4581;
      83520:data<=16'd5151;
      83521:data<=16'd6602;
      83522:data<=16'd7495;
      83523:data<=16'd6226;
      83524:data<=16'd6108;
      83525:data<=16'd6153;
      83526:data<=16'd5474;
      83527:data<=16'd6613;
      83528:data<=16'd7315;
      83529:data<=16'd7222;
      83530:data<=16'd7275;
      83531:data<=16'd6476;
      83532:data<=16'd6551;
      83533:data<=16'd6425;
      83534:data<=16'd7124;
      83535:data<=16'd8889;
      83536:data<=16'd4554;
      83537:data<=16'd2100;
      83538:data<=16'd10595;
      83539:data<=16'd16594;
      83540:data<=16'd16170;
      83541:data<=16'd16434;
      83542:data<=16'd15386;
      83543:data<=16'd14536;
      83544:data<=16'd14694;
      83545:data<=16'd13935;
      83546:data<=16'd14882;
      83547:data<=16'd14885;
      83548:data<=16'd13412;
      83549:data<=16'd13731;
      83550:data<=16'd12868;
      83551:data<=16'd11909;
      83552:data<=16'd12792;
      83553:data<=16'd12771;
      83554:data<=16'd12769;
      83555:data<=16'd12225;
      83556:data<=16'd10513;
      83557:data<=16'd10285;
      83558:data<=16'd11036;
      83559:data<=16'd12161;
      83560:data<=16'd12276;
      83561:data<=16'd10467;
      83562:data<=16'd9809;
      83563:data<=16'd9752;
      83564:data<=16'd9837;
      83565:data<=16'd11085;
      83566:data<=16'd10851;
      83567:data<=16'd10314;
      83568:data<=16'd10367;
      83569:data<=16'd9207;
      83570:data<=16'd8765;
      83571:data<=16'd8138;
      83572:data<=16'd7351;
      83573:data<=16'd7979;
      83574:data<=16'd6775;
      83575:data<=16'd5929;
      83576:data<=16'd6357;
      83577:data<=16'd4645;
      83578:data<=16'd4531;
      83579:data<=16'd1797;
      83580:data<=-16'd7997;
      83581:data<=-16'd13133;
      83582:data<=-16'd12029;
      83583:data<=-16'd12387;
      83584:data<=-16'd13352;
      83585:data<=-16'd14233;
      83586:data<=-16'd12333;
      83587:data<=-16'd7209;
      83588:data<=-16'd5736;
      83589:data<=-16'd7157;
      83590:data<=-16'd8017;
      83591:data<=-16'd8645;
      83592:data<=-16'd7834;
      83593:data<=-16'd7292;
      83594:data<=-16'd7614;
      83595:data<=-16'd7570;
      83596:data<=-16'd8778;
      83597:data<=-16'd9242;
      83598:data<=-16'd8222;
      83599:data<=-16'd8470;
      83600:data<=-16'd8546;
      83601:data<=-16'd8291;
      83602:data<=-16'd8887;
      83603:data<=-16'd9103;
      83604:data<=-16'd9309;
      83605:data<=-16'd9605;
      83606:data<=-16'd9347;
      83607:data<=-16'd8915;
      83608:data<=-16'd9294;
      83609:data<=-16'd10887;
      83610:data<=-16'd10912;
      83611:data<=-16'd9498;
      83612:data<=-16'd9209;
      83613:data<=-16'd8307;
      83614:data<=-16'd8698;
      83615:data<=-16'd11276;
      83616:data<=-16'd10778;
      83617:data<=-16'd9541;
      83618:data<=-16'd9724;
      83619:data<=-16'd8595;
      83620:data<=-16'd9485;
      83621:data<=-16'd9218;
      83622:data<=-16'd1921;
      83623:data<=16'd3974;
      83624:data<=16'd3783;
      83625:data<=16'd3579;
      83626:data<=16'd4109;
      83627:data<=16'd2649;
      83628:data<=16'd705;
      83629:data<=16'd808;
      83630:data<=16'd1172;
      83631:data<=16'd694;
      83632:data<=16'd1556;
      83633:data<=16'd746;
      83634:data<=-16'd1788;
      83635:data<=-16'd805;
      83636:data<=-16'd1583;
      83637:data<=-16'd6222;
      83638:data<=-16'd6678;
      83639:data<=-16'd5929;
      83640:data<=-16'd7908;
      83641:data<=-16'd7917;
      83642:data<=-16'd7363;
      83643:data<=-16'd7686;
      83644:data<=-16'd6699;
      83645:data<=-16'd6611;
      83646:data<=-16'd7747;
      83647:data<=-16'd8073;
      83648:data<=-16'd7761;
      83649:data<=-16'd7043;
      83650:data<=-16'd6428;
      83651:data<=-16'd6167;
      83652:data<=-16'd6943;
      83653:data<=-16'd8431;
      83654:data<=-16'd8052;
      83655:data<=-16'd7394;
      83656:data<=-16'd7507;
      83657:data<=-16'd6181;
      83658:data<=-16'd6355;
      83659:data<=-16'd7950;
      83660:data<=-16'd7447;
      83661:data<=-16'd7304;
      83662:data<=-16'd6774;
      83663:data<=-16'd6865;
      83664:data<=-16'd14016;
      83665:data<=-16'd21640;
      83666:data<=-16'd22048;
      83667:data<=-16'd20809;
      83668:data<=-16'd20101;
      83669:data<=-16'd18722;
      83670:data<=-16'd18327;
      83671:data<=-16'd17741;
      83672:data<=-16'd16466;
      83673:data<=-16'd15446;
      83674:data<=-16'd14311;
      83675:data<=-16'd13567;
      83676:data<=-16'd13141;
      83677:data<=-16'd11956;
      83678:data<=-16'd9990;
      83679:data<=-16'd8874;
      83680:data<=-16'd8945;
      83681:data<=-16'd8301;
      83682:data<=-16'd7808;
      83683:data<=-16'd7097;
      83684:data<=-16'd4611;
      83685:data<=-16'd4150;
      83686:data<=-16'd3436;
      83687:data<=16'd1744;
      83688:data<=16'd4162;
      83689:data<=16'd3172;
      83690:data<=16'd4611;
      83691:data<=16'd5460;
      83692:data<=16'd5272;
      83693:data<=16'd5934;
      83694:data<=16'd5780;
      83695:data<=16'd6049;
      83696:data<=16'd6854;
      83697:data<=16'd7743;
      83698:data<=16'd8746;
      83699:data<=16'd7964;
      83700:data<=16'd7447;
      83701:data<=16'd7649;
      83702:data<=16'd7636;
      83703:data<=16'd9703;
      83704:data<=16'd9658;
      83705:data<=16'd9103;
      83706:data<=16'd16609;
      83707:data<=16'd23951;
      83708:data<=16'd24178;
      83709:data<=16'd24486;
      83710:data<=16'd24811;
      83711:data<=16'd23302;
      83712:data<=16'd22600;
      83713:data<=16'd21608;
      83714:data<=16'd20560;
      83715:data<=16'd20697;
      83716:data<=16'd21067;
      83717:data<=16'd20905;
      83718:data<=16'd19835;
      83719:data<=16'd18891;
      83720:data<=16'd18352;
      83721:data<=16'd18657;
      83722:data<=16'd20104;
      83723:data<=16'd19479;
      83724:data<=16'd17992;
      83725:data<=16'd18010;
      83726:data<=16'd16666;
      83727:data<=16'd16358;
      83728:data<=16'd18067;
      83729:data<=16'd17120;
      83730:data<=16'd16014;
      83731:data<=16'd16354;
      83732:data<=16'd15440;
      83733:data<=16'd14994;
      83734:data<=16'd15766;
      83735:data<=16'd16557;
      83736:data<=16'd15121;
      83737:data<=16'd10440;
      83738:data<=16'd7539;
      83739:data<=16'd7206;
      83740:data<=16'd7373;
      83741:data<=16'd9125;
      83742:data<=16'd8614;
      83743:data<=16'd6601;
      83744:data<=16'd7374;
      83745:data<=16'd6540;
      83746:data<=16'd6484;
      83747:data<=16'd8631;
      83748:data<=16'd2099;
      83749:data<=-16'd7790;
      83750:data<=-16'd8587;
      83751:data<=-16'd6968;
      83752:data<=-16'd7494;
      83753:data<=-16'd6049;
      83754:data<=-16'd4728;
      83755:data<=-16'd4924;
      83756:data<=-16'd4546;
      83757:data<=-16'd4191;
      83758:data<=-16'd4247;
      83759:data<=-16'd3339;
      83760:data<=-16'd1976;
      83761:data<=-16'd2046;
      83762:data<=-16'd2776;
      83763:data<=-16'd2968;
      83764:data<=-16'd2968;
      83765:data<=-16'd1626;
      83766:data<=16'd77;
      83767:data<=-16'd397;
      83768:data<=-16'd1037;
      83769:data<=-16'd873;
      83770:data<=-16'd1257;
      83771:data<=-16'd1215;
      83772:data<=-16'd1233;
      83773:data<=-16'd1873;
      83774:data<=-16'd1882;
      83775:data<=-16'd1724;
      83776:data<=-16'd1638;
      83777:data<=-16'd2117;
      83778:data<=-16'd3415;
      83779:data<=-16'd3556;
      83780:data<=-16'd3588;
      83781:data<=-16'd4219;
      83782:data<=-16'd3853;
      83783:data<=-16'd4451;
      83784:data<=-16'd5441;
      83785:data<=-16'd5460;
      83786:data<=-16'd5937;
      83787:data<=-16'd3083;
      83788:data<=16'd687;
      83789:data<=-16'd285;
      83790:data<=16'd3556;
      83791:data<=16'd12548;
      83792:data<=16'd13590;
      83793:data<=16'd11094;
      83794:data<=16'd11903;
      83795:data<=16'd11291;
      83796:data<=16'd9556;
      83797:data<=16'd8164;
      83798:data<=16'd6740;
      83799:data<=16'd6529;
      83800:data<=16'd6244;
      83801:data<=16'd5970;
      83802:data<=16'd5553;
      83803:data<=16'd3750;
      83804:data<=16'd3102;
      83805:data<=16'd3181;
      83806:data<=16'd2390;
      83807:data<=16'd2359;
      83808:data<=16'd1980;
      83809:data<=16'd758;
      83810:data<=-16'd208;
      83811:data<=-16'd889;
      83812:data<=-16'd397;
      83813:data<=16'd129;
      83814:data<=-16'd140;
      83815:data<=-16'd1089;
      83816:data<=-16'd3283;
      83817:data<=-16'd3641;
      83818:data<=-16'd2660;
      83819:data<=-16'd3095;
      83820:data<=-16'd2544;
      83821:data<=-16'd3092;
      83822:data<=-16'd5194;
      83823:data<=-16'd4861;
      83824:data<=-16'd5054;
      83825:data<=-16'd5268;
      83826:data<=-16'd4182;
      83827:data<=-16'd5465;
      83828:data<=-16'd6123;
      83829:data<=-16'd6570;
      83830:data<=-16'd7498;
      83831:data<=-16'd5192;
      83832:data<=-16'd9229;
      83833:data<=-16'd19745;
      83834:data<=-16'd22536;
      83835:data<=-16'd21276;
      83836:data<=-16'd21453;
      83837:data<=-16'd22028;
      83838:data<=-16'd25370;
      83839:data<=-16'd25840;
      83840:data<=-16'd23877;
      83841:data<=-16'd25266;
      83842:data<=-16'd24595;
      83843:data<=-16'd23249;
      83844:data<=-16'd23919;
      83845:data<=-16'd22168;
      83846:data<=-16'd21625;
      83847:data<=-16'd22526;
      83848:data<=-16'd21393;
      83849:data<=-16'd21197;
      83850:data<=-16'd20756;
      83851:data<=-16'd19256;
      83852:data<=-16'd18898;
      83853:data<=-16'd19011;
      83854:data<=-16'd19549;
      83855:data<=-16'd18898;
      83856:data<=-16'd17540;
      83857:data<=-16'd17308;
      83858:data<=-16'd16054;
      83859:data<=-16'd16119;
      83860:data<=-16'd17553;
      83861:data<=-16'd16375;
      83862:data<=-16'd15503;
      83863:data<=-16'd14891;
      83864:data<=-16'd13675;
      83865:data<=-16'd14284;
      83866:data<=-16'd14040;
      83867:data<=-16'd13946;
      83868:data<=-16'd14358;
      83869:data<=-16'd12499;
      83870:data<=-16'd12516;
      83871:data<=-16'd11944;
      83872:data<=-16'd9773;
      83873:data<=-16'd11417;
      83874:data<=-16'd6549;
      83875:data<=16'd5103;
      83876:data<=16'd7570;
      83877:data<=16'd5967;
      83878:data<=16'd7923;
      83879:data<=16'd8199;
      83880:data<=16'd7840;
      83881:data<=16'd8043;
      83882:data<=16'd7656;
      83883:data<=16'd7806;
      83884:data<=16'd8566;
      83885:data<=16'd9509;
      83886:data<=16'd8981;
      83887:data<=16'd10152;
      83888:data<=16'd14924;
      83889:data<=16'd15975;
      83890:data<=16'd15091;
      83891:data<=16'd16859;
      83892:data<=16'd16483;
      83893:data<=16'd15982;
      83894:data<=16'd16788;
      83895:data<=16'd15241;
      83896:data<=16'd14904;
      83897:data<=16'd16078;
      83898:data<=16'd16078;
      83899:data<=16'd16161;
      83900:data<=16'd15666;
      83901:data<=16'd15306;
      83902:data<=16'd15291;
      83903:data<=16'd14948;
      83904:data<=16'd15649;
      83905:data<=16'd14886;
      83906:data<=16'd13623;
      83907:data<=16'd14128;
      83908:data<=16'd12906;
      83909:data<=16'd13063;
      83910:data<=16'd14963;
      83911:data<=16'd13547;
      83912:data<=16'd13345;
      83913:data<=16'd13368;
      83914:data<=16'd11409;
      83915:data<=16'd13267;
      83916:data<=16'd10319;
      83917:data<=-16'd522;
      83918:data<=-16'd3650;
      83919:data<=-16'd1037;
      83920:data<=-16'd2055;
      83921:data<=-16'd1673;
      83922:data<=16'd714;
      83923:data<=16'd1242;
      83924:data<=16'd1259;
      83925:data<=16'd1457;
      83926:data<=16'd875;
      83927:data<=16'd132;
      83928:data<=16'd1415;
      83929:data<=16'd3327;
      83930:data<=16'd2890;
      83931:data<=16'd2206;
      83932:data<=16'd2094;
      83933:data<=16'd1333;
      83934:data<=16'd1765;
      83935:data<=16'd3234;
      83936:data<=16'd3704;
      83937:data<=16'd1917;
      83938:data<=-16'd1733;
      83939:data<=-16'd3683;
      83940:data<=-16'd3218;
      83941:data<=-16'd2179;
      83942:data<=-16'd1237;
      83943:data<=-16'd1673;
      83944:data<=-16'd2046;
      83945:data<=-16'd1783;
      83946:data<=-16'd2146;
      83947:data<=-16'd318;
      83948:data<=16'd1310;
      83949:data<=-16'd252;
      83950:data<=-16'd55;
      83951:data<=16'd215;
      83952:data<=-16'd899;
      83953:data<=16'd1017;
      83954:data<=16'd1952;
      83955:data<=16'd1427;
      83956:data<=16'd2153;
      83957:data<=16'd368;
      83958:data<=16'd3459;
      83959:data<=16'd14436;
      83960:data<=16'd18777;
      83961:data<=16'd16636;
      83962:data<=16'd16813;
      83963:data<=16'd16108;
      83964:data<=16'd14269;
      83965:data<=16'd14286;
      83966:data<=16'd14927;
      83967:data<=16'd15230;
      83968:data<=16'd14654;
      83969:data<=16'd13952;
      83970:data<=16'd13174;
      83971:data<=16'd11814;
      83972:data<=16'd11718;
      83973:data<=16'd11805;
      83974:data<=16'd10774;
      83975:data<=16'd10249;
      83976:data<=16'd9650;
      83977:data<=16'd8969;
      83978:data<=16'd8322;
      83979:data<=16'd6583;
      83980:data<=16'd5439;
      83981:data<=16'd5474;
      83982:data<=16'd5494;
      83983:data<=16'd5253;
      83984:data<=16'd4372;
      83985:data<=16'd3377;
      83986:data<=16'd2338;
      83987:data<=16'd3210;
      83988:data<=16'd7216;
      83989:data<=16'd8381;
      83990:data<=16'd6443;
      83991:data<=16'd5888;
      83992:data<=16'd4381;
      83993:data<=16'd3595;
      83994:data<=16'd4400;
      83995:data<=16'd3253;
      83996:data<=16'd3475;
      83997:data<=16'd2860;
      83998:data<=16'd197;
      83999:data<=16'd1994;
      84000:data<=-16'd1351;
      84001:data<=-16'd12668;
      84002:data<=-16'd15722;
      84003:data<=-16'd14029;
      84004:data<=-16'd15955;
      84005:data<=-16'd15390;
      84006:data<=-16'd14537;
      84007:data<=-16'd15437;
      84008:data<=-16'd14287;
      84009:data<=-16'd14060;
      84010:data<=-16'd15320;
      84011:data<=-16'd15370;
      84012:data<=-16'd14698;
      84013:data<=-16'd13847;
      84014:data<=-16'd13362;
      84015:data<=-16'd13279;
      84016:data<=-16'd14131;
      84017:data<=-16'd15208;
      84018:data<=-16'd14108;
      84019:data<=-16'd13201;
      84020:data<=-16'd13183;
      84021:data<=-16'd11958;
      84022:data<=-16'd12660;
      84023:data<=-16'd14507;
      84024:data<=-16'd13671;
      84025:data<=-16'd12800;
      84026:data<=-16'd12916;
      84027:data<=-16'd12336;
      84028:data<=-16'd12516;
      84029:data<=-16'd13970;
      84030:data<=-16'd13973;
      84031:data<=-16'd12104;
      84032:data<=-16'd11963;
      84033:data<=-16'd12440;
      84034:data<=-16'd11477;
      84035:data<=-16'd12484;
      84036:data<=-16'd12807;
      84037:data<=-16'd12457;
      84038:data<=-16'd17305;
      84039:data<=-16'd18824;
      84040:data<=-16'd15814;
      84041:data<=-16'd18713;
      84042:data<=-16'd15960;
      84043:data<=-16'd3770;
      84044:data<=-16'd341;
      84045:data<=-16'd2591;
      84046:data<=-16'd1014;
      84047:data<=-16'd1698;
      84048:data<=-16'd3806;
      84049:data<=-16'd3591;
      84050:data<=-16'd3397;
      84051:data<=-16'd3151;
      84052:data<=-16'd2455;
      84053:data<=-16'd2426;
      84054:data<=-16'd3899;
      84055:data<=-16'd5319;
      84056:data<=-16'd4519;
      84057:data<=-16'd3653;
      84058:data<=-16'd3369;
      84059:data<=-16'd3090;
      84060:data<=-16'd4593;
      84061:data<=-16'd5350;
      84062:data<=-16'd4211;
      84063:data<=-16'd4156;
      84064:data<=-16'd3873;
      84065:data<=-16'd3142;
      84066:data<=-16'd3809;
      84067:data<=-16'd4355;
      84068:data<=-16'd4228;
      84069:data<=-16'd4015;
      84070:data<=-16'd3755;
      84071:data<=-16'd3254;
      84072:data<=-16'd2541;
      84073:data<=-16'd3089;
      84074:data<=-16'd3483;
      84075:data<=-16'd2390;
      84076:data<=-16'd2070;
      84077:data<=-16'd1460;
      84078:data<=-16'd253;
      84079:data<=16'd320;
      84080:data<=16'd1794;
      84081:data<=16'd1768;
      84082:data<=16'd1394;
      84083:data<=16'd3845;
      84084:data<=16'd652;
      84085:data<=-16'd8141;
      84086:data<=-16'd10862;
      84087:data<=-16'd8146;
      84088:data<=-16'd4390;
      84089:data<=-16'd1145;
      84090:data<=-16'd954;
      84091:data<=-16'd229;
      84092:data<=16'd1635;
      84093:data<=16'd1201;
      84094:data<=16'd1394;
      84095:data<=16'd2362;
      84096:data<=16'd2170;
      84097:data<=16'd3086;
      84098:data<=16'd4487;
      84099:data<=16'd4866;
      84100:data<=16'd4987;
      84101:data<=16'd5151;
      84102:data<=16'd5426;
      84103:data<=16'd5705;
      84104:data<=16'd6667;
      84105:data<=16'd7467;
      84106:data<=16'd6949;
      84107:data<=16'd7075;
      84108:data<=16'd6881;
      84109:data<=16'd6103;
      84110:data<=16'd7539;
      84111:data<=16'd8246;
      84112:data<=16'd7423;
      84113:data<=16'd7928;
      84114:data<=16'd7600;
      84115:data<=16'd7219;
      84116:data<=16'd8420;
      84117:data<=16'd8836;
      84118:data<=16'd8971;
      84119:data<=16'd8805;
      84120:data<=16'd8210;
      84121:data<=16'd8062;
      84122:data<=16'd7791;
      84123:data<=16'd9961;
      84124:data<=16'd11394;
      84125:data<=16'd8549;
      84126:data<=16'd11975;
      84127:data<=16'd21328;
      84128:data<=16'd24386;
      84129:data<=16'd23911;
      84130:data<=16'd23860;
      84131:data<=16'd22375;
      84132:data<=16'd21552;
      84133:data<=16'd20660;
      84134:data<=16'd19849;
      84135:data<=16'd20842;
      84136:data<=16'd21146;
      84137:data<=16'd19716;
      84138:data<=16'd15984;
      84139:data<=16'd11476;
      84140:data<=16'd10223;
      84141:data<=16'd11010;
      84142:data<=16'd12160;
      84143:data<=16'd12505;
      84144:data<=16'd11015;
      84145:data<=16'd10571;
      84146:data<=16'd10128;
      84147:data<=16'd9629;
      84148:data<=16'd11546;
      84149:data<=16'd11071;
      84150:data<=16'd9468;
      84151:data<=16'd10511;
      84152:data<=16'd9276;
      84153:data<=16'd8834;
      84154:data<=16'd11426;
      84155:data<=16'd10781;
      84156:data<=16'd9781;
      84157:data<=16'd10219;
      84158:data<=16'd8990;
      84159:data<=16'd8702;
      84160:data<=16'd9389;
      84161:data<=16'd9956;
      84162:data<=16'd10260;
      84163:data<=16'd9295;
      84164:data<=16'd9239;
      84165:data<=16'd8419;
      84166:data<=16'd7738;
      84167:data<=16'd10840;
      84168:data<=16'd7717;
      84169:data<=-16'd2796;
      84170:data<=-16'd6959;
      84171:data<=-16'd6598;
      84172:data<=-16'd7335;
      84173:data<=-16'd6316;
      84174:data<=-16'd5683;
      84175:data<=-16'd6337;
      84176:data<=-16'd6115;
      84177:data<=-16'd5770;
      84178:data<=-16'd5935;
      84179:data<=-16'd6931;
      84180:data<=-16'd7371;
      84181:data<=-16'd6607;
      84182:data<=-16'd6328;
      84183:data<=-16'd6378;
      84184:data<=-16'd7060;
      84185:data<=-16'd7762;
      84186:data<=-16'd7940;
      84187:data<=-16'd8668;
      84188:data<=-16'd6099;
      84189:data<=-16'd1554;
      84190:data<=-16'd1481;
      84191:data<=-16'd2282;
      84192:data<=-16'd2699;
      84193:data<=-16'd4946;
      84194:data<=-16'd4828;
      84195:data<=-16'd3903;
      84196:data<=-16'd4197;
      84197:data<=-16'd3849;
      84198:data<=-16'd5241;
      84199:data<=-16'd5868;
      84200:data<=-16'd4751;
      84201:data<=-16'd5642;
      84202:data<=-16'd5110;
      84203:data<=-16'd4922;
      84204:data<=-16'd7777;
      84205:data<=-16'd7905;
      84206:data<=-16'd7623;
      84207:data<=-16'd8210;
      84208:data<=-16'd6858;
      84209:data<=-16'd8040;
      84210:data<=-16'd6519;
      84211:data<=16'd1994;
      84212:data<=16'd6035;
      84213:data<=16'd5012;
      84214:data<=16'd5826;
      84215:data<=16'd5909;
      84216:data<=16'd4059;
      84217:data<=16'd1953;
      84218:data<=16'd998;
      84219:data<=16'd1292;
      84220:data<=16'd990;
      84221:data<=16'd1451;
      84222:data<=16'd1278;
      84223:data<=-16'd1791;
      84224:data<=-16'd2816;
      84225:data<=-16'd1290;
      84226:data<=-16'd1049;
      84227:data<=-16'd1111;
      84228:data<=-16'd1389;
      84229:data<=-16'd2789;
      84230:data<=-16'd4165;
      84231:data<=-16'd4447;
      84232:data<=-16'd4147;
      84233:data<=-16'd4397;
      84234:data<=-16'd3896;
      84235:data<=-16'd3920;
      84236:data<=-16'd5673;
      84237:data<=-16'd5071;
      84238:data<=-16'd6012;
      84239:data<=-16'd11227;
      84240:data<=-16'd12000;
      84241:data<=-16'd11095;
      84242:data<=-16'd13643;
      84243:data<=-16'd13191;
      84244:data<=-16'd11828;
      84245:data<=-16'd12255;
      84246:data<=-16'd11035;
      84247:data<=-16'd11329;
      84248:data<=-16'd12468;
      84249:data<=-16'd12058;
      84250:data<=-16'd11899;
      84251:data<=-16'd10144;
      84252:data<=-16'd11899;
      84253:data<=-16'd20862;
      84254:data<=-16'd26497;
      84255:data<=-16'd26248;
      84256:data<=-16'd25529;
      84257:data<=-16'd24004;
      84258:data<=-16'd22360;
      84259:data<=-16'd21276;
      84260:data<=-16'd20945;
      84261:data<=-16'd21820;
      84262:data<=-16'd21073;
      84263:data<=-16'd19637;
      84264:data<=-16'd19246;
      84265:data<=-16'd17805;
      84266:data<=-16'd17224;
      84267:data<=-16'd18410;
      84268:data<=-16'd18210;
      84269:data<=-16'd16844;
      84270:data<=-16'd15973;
      84271:data<=-16'd15808;
      84272:data<=-16'd15247;
      84273:data<=-16'd13781;
      84274:data<=-16'd12986;
      84275:data<=-16'd12587;
      84276:data<=-16'd11956;
      84277:data<=-16'd11624;
      84278:data<=-16'd10678;
      84279:data<=-16'd9186;
      84280:data<=-16'd7771;
      84281:data<=-16'd6751;
      84282:data<=-16'd6291;
      84283:data<=-16'd5498;
      84284:data<=-16'd5338;
      84285:data<=-16'd4570;
      84286:data<=-16'd2027;
      84287:data<=-16'd2029;
      84288:data<=-16'd587;
      84289:data<=16'd5253;
      84290:data<=16'd5968;
      84291:data<=16'd5295;
      84292:data<=16'd8907;
      84293:data<=16'd7768;
      84294:data<=16'd8273;
      84295:data<=16'd17879;
      84296:data<=16'd23058;
      84297:data<=16'd22037;
      84298:data<=16'd23085;
      84299:data<=16'd23322;
      84300:data<=16'd22078;
      84301:data<=16'd21793;
      84302:data<=16'd20952;
      84303:data<=16'd19640;
      84304:data<=16'd19331;
      84305:data<=16'd19980;
      84306:data<=16'd19687;
      84307:data<=16'd18125;
      84308:data<=16'd17062;
      84309:data<=16'd16419;
      84310:data<=16'd17171;
      84311:data<=16'd18900;
      84312:data<=16'd18137;
      84313:data<=16'd16772;
      84314:data<=16'd16551;
      84315:data<=16'd15414;
      84316:data<=16'd15529;
      84317:data<=16'd17058;
      84318:data<=16'd16584;
      84319:data<=16'd15596;
      84320:data<=16'd15421;
      84321:data<=16'd14572;
      84322:data<=16'd13928;
      84323:data<=16'd14725;
      84324:data<=16'd15440;
      84325:data<=16'd14865;
      84326:data<=16'd14340;
      84327:data<=16'd13409;
      84328:data<=16'd11397;
      84329:data<=16'd11837;
      84330:data<=16'd13773;
      84331:data<=16'd12975;
      84332:data<=16'd12023;
      84333:data<=16'd11700;
      84334:data<=16'd10317;
      84335:data<=16'd11267;
      84336:data<=16'd11576;
      84337:data<=16'd4595;
      84338:data<=-16'd4636;
      84339:data<=-16'd9273;
      84340:data<=-16'd10288;
      84341:data<=-16'd9407;
      84342:data<=-16'd7679;
      84343:data<=-16'd6815;
      84344:data<=-16'd6819;
      84345:data<=-16'd6435;
      84346:data<=-16'd5717;
      84347:data<=-16'd5386;
      84348:data<=-16'd4387;
      84349:data<=-16'd2889;
      84350:data<=-16'd3118;
      84351:data<=-16'd3870;
      84352:data<=-16'd3688;
      84353:data<=-16'd3870;
      84354:data<=-16'd2955;
      84355:data<=-16'd758;
      84356:data<=-16'd370;
      84357:data<=-16'd358;
      84358:data<=16'd253;
      84359:data<=-16'd852;
      84360:data<=-16'd1057;
      84361:data<=16'd893;
      84362:data<=16'd1102;
      84363:data<=16'd466;
      84364:data<=16'd892;
      84365:data<=16'd359;
      84366:data<=16'd217;
      84367:data<=16'd2055;
      84368:data<=16'd2814;
      84369:data<=16'd2278;
      84370:data<=16'd2789;
      84371:data<=16'd2776;
      84372:data<=16'd1701;
      84373:data<=16'd1750;
      84374:data<=16'd1510;
      84375:data<=16'd646;
      84376:data<=16'd1436;
      84377:data<=16'd1127;
      84378:data<=16'd955;
      84379:data<=16'd7492;
      84380:data<=16'd14604;
      84381:data<=16'd14401;
      84382:data<=16'd13245;
      84383:data<=16'd14122;
      84384:data<=16'd12903;
      84385:data<=16'd11032;
      84386:data<=16'd9600;
      84387:data<=16'd7682;
      84388:data<=16'd7846;
      84389:data<=16'd10229;
      84390:data<=16'd11138;
      84391:data<=16'd9565;
      84392:data<=16'd7714;
      84393:data<=16'd6874;
      84394:data<=16'd6296;
      84395:data<=16'd5527;
      84396:data<=16'd4996;
      84397:data<=16'd4749;
      84398:data<=16'd3908;
      84399:data<=16'd2165;
      84400:data<=16'd1327;
      84401:data<=16'd1639;
      84402:data<=16'd1580;
      84403:data<=16'd1571;
      84404:data<=16'd607;
      84405:data<=-16'd1721;
      84406:data<=-16'd2231;
      84407:data<=-16'd1888;
      84408:data<=-16'd2476;
      84409:data<=-16'd2279;
      84410:data<=-16'd3093;
      84411:data<=-16'd4949;
      84412:data<=-16'd4760;
      84413:data<=-16'd4399;
      84414:data<=-16'd4620;
      84415:data<=-16'd4093;
      84416:data<=-16'd4275;
      84417:data<=-16'd5307;
      84418:data<=-16'd6542;
      84419:data<=-16'd6460;
      84420:data<=-16'd5896;
      84421:data<=-16'd11521;
      84422:data<=-16'd20183;
      84423:data<=-16'd22268;
      84424:data<=-16'd21399;
      84425:data<=-16'd21713;
      84426:data<=-16'd20521;
      84427:data<=-16'd19603;
      84428:data<=-16'd19608;
      84429:data<=-16'd19396;
      84430:data<=-16'd19701;
      84431:data<=-16'd18907;
      84432:data<=-16'd18145;
      84433:data<=-16'd18387;
      84434:data<=-16'd16833;
      84435:data<=-16'd16487;
      84436:data<=-16'd18284;
      84437:data<=-16'd17250;
      84438:data<=-16'd16639;
      84439:data<=-16'd19394;
      84440:data<=-16'd20137;
      84441:data<=-16'd18824;
      84442:data<=-16'd19168;
      84443:data<=-16'd19748;
      84444:data<=-16'd19147;
      84445:data<=-16'd18568;
      84446:data<=-16'd17945;
      84447:data<=-16'd16783;
      84448:data<=-16'd16574;
      84449:data<=-16'd17273;
      84450:data<=-16'd16697;
      84451:data<=-16'd15465;
      84452:data<=-16'd14687;
      84453:data<=-16'd13896;
      84454:data<=-16'd13967;
      84455:data<=-16'd14515;
      84456:data<=-16'd13996;
      84457:data<=-16'd13121;
      84458:data<=-16'd12944;
      84459:data<=-16'd12894;
      84460:data<=-16'd11858;
      84461:data<=-16'd12155;
      84462:data<=-16'd13791;
      84463:data<=-16'd8197;
      84464:data<=16'd2438;
      84465:data<=16'd5184;
      84466:data<=16'd3394;
      84467:data<=16'd3906;
      84468:data<=16'd2505;
      84469:data<=16'd1309;
      84470:data<=16'd2544;
      84471:data<=16'd2005;
      84472:data<=16'd1309;
      84473:data<=16'd1797;
      84474:data<=16'd1903;
      84475:data<=16'd2361;
      84476:data<=16'd2323;
      84477:data<=16'd2074;
      84478:data<=16'd2831;
      84479:data<=16'd3792;
      84480:data<=16'd4981;
      84481:data<=16'd5388;
      84482:data<=16'd5212;
      84483:data<=16'd5674;
      84484:data<=16'd5063;
      84485:data<=16'd5239;
      84486:data<=16'd7495;
      84487:data<=16'd7876;
      84488:data<=16'd7938;
      84489:data<=16'd10320;
      84490:data<=16'd11714;
      84491:data<=16'd11257;
      84492:data<=16'd11549;
      84493:data<=16'd12715;
      84494:data<=16'd12525;
      84495:data<=16'd11699;
      84496:data<=16'd11750;
      84497:data<=16'd11004;
      84498:data<=16'd11388;
      84499:data<=16'd13280;
      84500:data<=16'd12742;
      84501:data<=16'd12731;
      84502:data<=16'd12968;
      84503:data<=16'd11647;
      84504:data<=16'd13994;
      84505:data<=16'd11344;
      84506:data<=-16'd317;
      84507:data<=-16'd3524;
      84508:data<=-16'd347;
      84509:data<=-16'd2021;
      84510:data<=-16'd1337;
      84511:data<=16'd1207;
      84512:data<=16'd1014;
      84513:data<=16'd1932;
      84514:data<=16'd2649;
      84515:data<=16'd2285;
      84516:data<=16'd2188;
      84517:data<=16'd2716;
      84518:data<=16'd4767;
      84519:data<=16'd4528;
      84520:data<=16'd3102;
      84521:data<=16'd4435;
      84522:data<=16'd4349;
      84523:data<=16'd4253;
      84524:data<=16'd6513;
      84525:data<=16'd6517;
      84526:data<=16'd5996;
      84527:data<=16'd6328;
      84528:data<=16'd5526;
      84529:data<=16'd5982;
      84530:data<=16'd7263;
      84531:data<=16'd7670;
      84532:data<=16'd7611;
      84533:data<=16'd7013;
      84534:data<=16'd6981;
      84535:data<=16'd7006;
      84536:data<=16'd7436;
      84537:data<=16'd8856;
      84538:data<=16'd7999;
      84539:data<=16'd5709;
      84540:data<=16'd3946;
      84541:data<=16'd2761;
      84542:data<=16'd3870;
      84543:data<=16'd4147;
      84544:data<=16'd3436;
      84545:data<=16'd4085;
      84546:data<=16'd2484;
      84547:data<=16'd6026;
      84548:data<=16'd17835;
      84549:data<=16'd21719;
      84550:data<=16'd18541;
      84551:data<=16'd19096;
      84552:data<=16'd18489;
      84553:data<=16'd16428;
      84554:data<=16'd16684;
      84555:data<=16'd16980;
      84556:data<=16'd16913;
      84557:data<=16'd16002;
      84558:data<=16'd15292;
      84559:data<=16'd15097;
      84560:data<=16'd13397;
      84561:data<=16'd13832;
      84562:data<=16'd15456;
      84563:data<=16'd13981;
      84564:data<=16'd13327;
      84565:data<=16'd13306;
      84566:data<=16'd11776;
      84567:data<=16'd12029;
      84568:data<=16'd12725;
      84569:data<=16'd12205;
      84570:data<=16'd11834;
      84571:data<=16'd11189;
      84572:data<=16'd10636;
      84573:data<=16'd9735;
      84574:data<=16'd8454;
      84575:data<=16'd8135;
      84576:data<=16'd7868;
      84577:data<=16'd7614;
      84578:data<=16'd7204;
      84579:data<=16'd6049;
      84580:data<=16'd5156;
      84581:data<=16'd3850;
      84582:data<=16'd3137;
      84583:data<=16'd3347;
      84584:data<=16'd2601;
      84585:data<=16'd3240;
      84586:data<=16'd2817;
      84587:data<=-16'd117;
      84588:data<=16'd858;
      84589:data<=-16'd995;
      84590:data<=-16'd9423;
      84591:data<=-16'd11605;
      84592:data<=-16'd10534;
      84593:data<=-16'd13147;
      84594:data<=-16'd12536;
      84595:data<=-16'd11015;
      84596:data<=-16'd11793;
      84597:data<=-16'd11217;
      84598:data<=-16'd11543;
      84599:data<=-16'd12199;
      84600:data<=-16'd11658;
      84601:data<=-16'd12002;
      84602:data<=-16'd11461;
      84603:data<=-16'd10977;
      84604:data<=-16'd11949;
      84605:data<=-16'd12290;
      84606:data<=-16'd13141;
      84607:data<=-16'd13362;
      84608:data<=-16'd11922;
      84609:data<=-16'd11596;
      84610:data<=-16'd11224;
      84611:data<=-16'd11204;
      84612:data<=-16'd12571;
      84613:data<=-16'd12223;
      84614:data<=-16'd11800;
      84615:data<=-16'd12205;
      84616:data<=-16'd10901;
      84617:data<=-16'd10828;
      84618:data<=-16'd12513;
      84619:data<=-16'd12411;
      84620:data<=-16'd11546;
      84621:data<=-16'd11233;
      84622:data<=-16'd10695;
      84623:data<=-16'd10683;
      84624:data<=-16'd11906;
      84625:data<=-16'd12260;
      84626:data<=-16'd11221;
      84627:data<=-16'd11517;
      84628:data<=-16'd11160;
      84629:data<=-16'd10326;
      84630:data<=-16'd13026;
      84631:data<=-16'd9953;
      84632:data<=16'd1421;
      84633:data<=16'd4589;
      84634:data<=16'd1477;
      84635:data<=16'd3160;
      84636:data<=16'd2500;
      84637:data<=-16'd356;
      84638:data<=16'd839;
      84639:data<=-16'd393;
      84640:data<=-16'd4523;
      84641:data<=-16'd5180;
      84642:data<=-16'd4516;
      84643:data<=-16'd5591;
      84644:data<=-16'd6343;
      84645:data<=-16'd5582;
      84646:data<=-16'd5160;
      84647:data<=-16'd4916;
      84648:data<=-16'd4029;
      84649:data<=-16'd5100;
      84650:data<=-16'd6705;
      84651:data<=-16'd6079;
      84652:data<=-16'd6011;
      84653:data<=-16'd6087;
      84654:data<=-16'd5095;
      84655:data<=-16'd5583;
      84656:data<=-16'd6152;
      84657:data<=-16'd5776;
      84658:data<=-16'd6134;
      84659:data<=-16'd6106;
      84660:data<=-16'd5318;
      84661:data<=-16'd5207;
      84662:data<=-16'd6132;
      84663:data<=-16'd6552;
      84664:data<=-16'd5949;
      84665:data<=-16'd6209;
      84666:data<=-16'd5774;
      84667:data<=-16'd4972;
      84668:data<=-16'd6742;
      84669:data<=-16'd6981;
      84670:data<=-16'd6190;
      84671:data<=-16'd6722;
      84672:data<=-16'd4131;
      84673:data<=-16'd6642;
      84674:data<=-16'd17352;
      84675:data<=-16'd20281;
      84676:data<=-16'd17523;
      84677:data<=-16'd18174;
      84678:data<=-16'd16547;
      84679:data<=-16'd14371;
      84680:data<=-16'd13671;
      84681:data<=-16'd11441;
      84682:data<=-16'd10916;
      84683:data<=-16'd10237;
      84684:data<=-16'd8674;
      84685:data<=-16'd9266;
      84686:data<=-16'd7485;
      84687:data<=-16'd5277;
      84688:data<=-16'd6291;
      84689:data<=-16'd4458;
      84690:data<=-16'd637;
      84691:data<=16'd764;
      84692:data<=16'd1521;
      84693:data<=16'd2358;
      84694:data<=16'd2927;
      84695:data<=16'd3031;
      84696:data<=16'd3139;
      84697:data<=16'd3466;
      84698:data<=16'd2898;
      84699:data<=16'd3454;
      84700:data<=16'd5107;
      84701:data<=16'd5262;
      84702:data<=16'd5359;
      84703:data<=16'd5256;
      84704:data<=16'd5042;
      84705:data<=16'd6351;
      84706:data<=16'd6790;
      84707:data<=16'd6382;
      84708:data<=16'd6416;
      84709:data<=16'd6432;
      84710:data<=16'd7241;
      84711:data<=16'd7121;
      84712:data<=16'd7213;
      84713:data<=16'd8113;
      84714:data<=16'd6360;
      84715:data<=16'd10088;
      84716:data<=16'd20673;
      84717:data<=16'd23605;
      84718:data<=16'd21755;
      84719:data<=16'd22962;
      84720:data<=16'd22149;
      84721:data<=16'd20838;
      84722:data<=16'd20442;
      84723:data<=16'd19091;
      84724:data<=16'd19904;
      84725:data<=16'd20381;
      84726:data<=16'd19005;
      84727:data<=16'd18924;
      84728:data<=16'd18215;
      84729:data<=16'd17124;
      84730:data<=16'd17170;
      84731:data<=16'd17183;
      84732:data<=16'd17478;
      84733:data<=16'd16683;
      84734:data<=16'd15277;
      84735:data<=16'd15015;
      84736:data<=16'd14219;
      84737:data<=16'd14427;
      84738:data<=16'd15723;
      84739:data<=16'd14116;
      84740:data<=16'd10739;
      84741:data<=16'd8526;
      84742:data<=16'd8426;
      84743:data<=16'd9491;
      84744:data<=16'd9708;
      84745:data<=16'd9855;
      84746:data<=16'd9530;
      84747:data<=16'd8387;
      84748:data<=16'd8254;
      84749:data<=16'd8181;
      84750:data<=16'd8739;
      84751:data<=16'd9360;
      84752:data<=16'd7985;
      84753:data<=16'd8244;
      84754:data<=16'd8096;
      84755:data<=16'd6537;
      84756:data<=16'd9477;
      84757:data<=16'd7174;
      84758:data<=-16'd4037;
      84759:data<=-16'd8100;
      84760:data<=-16'd6969;
      84761:data<=-16'd7971;
      84762:data<=-16'd5592;
      84763:data<=-16'd3741;
      84764:data<=-16'd4728;
      84765:data<=-16'd4276;
      84766:data<=-16'd4992;
      84767:data<=-16'd5039;
      84768:data<=-16'd2866;
      84769:data<=-16'd2576;
      84770:data<=-16'd2549;
      84771:data<=-16'd2408;
      84772:data<=-16'd3080;
      84773:data<=-16'd2641;
      84774:data<=-16'd2892;
      84775:data<=-16'd3307;
      84776:data<=-16'd2384;
      84777:data<=-16'd2616;
      84778:data<=-16'd2864;
      84779:data<=-16'd2541;
      84780:data<=-16'd3689;
      84781:data<=-16'd5068;
      84782:data<=-16'd5762;
      84783:data<=-16'd5629;
      84784:data<=-16'd5137;
      84785:data<=-16'd5589;
      84786:data<=-16'd5879;
      84787:data<=-16'd6393;
      84788:data<=-16'd7483;
      84789:data<=-16'd6326;
      84790:data<=-16'd3482;
      84791:data<=-16'd1812;
      84792:data<=-16'd2190;
      84793:data<=-16'd3444;
      84794:data<=-16'd4061;
      84795:data<=-16'd4940;
      84796:data<=-16'd5090;
      84797:data<=-16'd4567;
      84798:data<=-16'd6172;
      84799:data<=-16'd3556;
      84800:data<=16'd5497;
      84801:data<=16'd9341;
      84802:data<=16'd7262;
      84803:data<=16'd6768;
      84804:data<=16'd6651;
      84805:data<=16'd5594;
      84806:data<=16'd3990;
      84807:data<=16'd2508;
      84808:data<=16'd2696;
      84809:data<=16'd2588;
      84810:data<=16'd2262;
      84811:data<=16'd2452;
      84812:data<=16'd851;
      84813:data<=-16'd493;
      84814:data<=-16'd165;
      84815:data<=-16'd132;
      84816:data<=16'd161;
      84817:data<=-16'd261;
      84818:data<=-16'd2112;
      84819:data<=-16'd3192;
      84820:data<=-16'd3301;
      84821:data<=-16'd3245;
      84822:data<=-16'd3206;
      84823:data<=-16'd2673;
      84824:data<=-16'd2444;
      84825:data<=-16'd4017;
      84826:data<=-16'd4720;
      84827:data<=-16'd4404;
      84828:data<=-16'd4951;
      84829:data<=-16'd4091;
      84830:data<=-16'd4282;
      84831:data<=-16'd6488;
      84832:data<=-16'd6357;
      84833:data<=-16'd6545;
      84834:data<=-16'd6731;
      84835:data<=-16'd4827;
      84836:data<=-16'd5999;
      84837:data<=-16'd7564;
      84838:data<=-16'd6901;
      84839:data<=-16'd7862;
      84840:data<=-16'd8583;
      84841:data<=-16'd12833;
      84842:data<=-16'd22315;
      84843:data<=-16'd26605;
      84844:data<=-16'd26040;
      84845:data<=-16'd25569;
      84846:data<=-16'd23808;
      84847:data<=-16'd22748;
      84848:data<=-16'd21717;
      84849:data<=-16'd20912;
      84850:data<=-16'd22469;
      84851:data<=-16'd21704;
      84852:data<=-16'd19488;
      84853:data<=-16'd19123;
      84854:data<=-16'd17888;
      84855:data<=-16'd17584;
      84856:data<=-16'd18466;
      84857:data<=-16'd17776;
      84858:data<=-16'd17098;
      84859:data<=-16'd16110;
      84860:data<=-16'd15091;
      84861:data<=-16'd15173;
      84862:data<=-16'd14715;
      84863:data<=-16'd14540;
      84864:data<=-16'd14592;
      84865:data<=-16'd14286;
      84866:data<=-16'd14313;
      84867:data<=-16'd13026;
      84868:data<=-16'd12373;
      84869:data<=-16'd13251;
      84870:data<=-16'd12463;
      84871:data<=-16'd11888;
      84872:data<=-16'd11588;
      84873:data<=-16'd10313;
      84874:data<=-16'd10379;
      84875:data<=-16'd9885;
      84876:data<=-16'd8895;
      84877:data<=-16'd8552;
      84878:data<=-16'd6816;
      84879:data<=-16'd6607;
      84880:data<=-16'd6155;
      84881:data<=-16'd3401;
      84882:data<=-16'd4211;
      84883:data<=-16'd1566;
      84884:data<=16'd9027;
      84885:data<=16'd13796;
      84886:data<=16'd12511;
      84887:data<=16'd13941;
      84888:data<=16'd14612;
      84889:data<=16'd13611;
      84890:data<=16'd14936;
      84891:data<=16'd17350;
      84892:data<=16'd17616;
      84893:data<=16'd16760;
      84894:data<=16'd17608;
      84895:data<=16'd17653;
      84896:data<=16'd16302;
      84897:data<=16'd16452;
      84898:data<=16'd15661;
      84899:data<=16'd14871;
      84900:data<=16'd16631;
      84901:data<=16'd16836;
      84902:data<=16'd15998;
      84903:data<=16'd15945;
      84904:data<=16'd14707;
      84905:data<=16'd14668;
      84906:data<=16'd16158;
      84907:data<=16'd16563;
      84908:data<=16'd16271;
      84909:data<=16'd15161;
      84910:data<=16'd14298;
      84911:data<=16'd14390;
      84912:data<=16'd14436;
      84913:data<=16'd15003;
      84914:data<=16'd14753;
      84915:data<=16'd14298;
      84916:data<=16'd14953;
      84917:data<=16'd13623;
      84918:data<=16'd12916;
      84919:data<=16'd14264;
      84920:data<=16'd13221;
      84921:data<=16'd13267;
      84922:data<=16'd13872;
      84923:data<=16'd11341;
      84924:data<=16'd12616;
      84925:data<=16'd12895;
      84926:data<=16'd3824;
      84927:data<=-16'd2387;
      84928:data<=-16'd1551;
      84929:data<=-16'd2165;
      84930:data<=-16'd1798;
      84931:data<=16'd767;
      84932:data<=16'd1281;
      84933:data<=16'd778;
      84934:data<=16'd499;
      84935:data<=16'd455;
      84936:data<=16'd723;
      84937:data<=16'd1052;
      84938:data<=16'd2390;
      84939:data<=16'd3266;
      84940:data<=16'd1506;
      84941:data<=-16'd1485;
      84942:data<=-16'd3165;
      84943:data<=-16'd2014;
      84944:data<=-16'd76;
      84945:data<=16'd309;
      84946:data<=16'd719;
      84947:data<=16'd772;
      84948:data<=-16'd88;
      84949:data<=16'd717;
      84950:data<=16'd1892;
      84951:data<=16'd1645;
      84952:data<=16'd1760;
      84953:data<=16'd1847;
      84954:data<=16'd1457;
      84955:data<=16'd1851;
      84956:data<=16'd2372;
      84957:data<=16'd2367;
      84958:data<=16'd2557;
      84959:data<=16'd2977;
      84960:data<=16'd2608;
      84961:data<=16'd2032;
      84962:data<=16'd3028;
      84963:data<=16'd4073;
      84964:data<=16'd4294;
      84965:data<=16'd4484;
      84966:data<=16'd2690;
      84967:data<=16'd3768;
      84968:data<=16'd13347;
      84969:data<=16'd20732;
      84970:data<=16'd19308;
      84971:data<=16'd17666;
      84972:data<=16'd17370;
      84973:data<=16'd15920;
      84974:data<=16'd15491;
      84975:data<=16'd14722;
      84976:data<=16'd13653;
      84977:data<=16'd13809;
      84978:data<=16'd12706;
      84979:data<=16'd11555;
      84980:data<=16'd11611;
      84981:data<=16'd9627;
      84982:data<=16'd7377;
      84983:data<=16'd7679;
      84984:data<=16'd7709;
      84985:data<=16'd6623;
      84986:data<=16'd6328;
      84987:data<=16'd5859;
      84988:data<=16'd3871;
      84989:data<=16'd2497;
      84990:data<=16'd3959;
      84991:data<=16'd6463;
      84992:data<=16'd7236;
      84993:data<=16'd5979;
      84994:data<=16'd4052;
      84995:data<=16'd3071;
      84996:data<=16'd3080;
      84997:data<=16'd3058;
      84998:data<=16'd2948;
      84999:data<=16'd2494;
      85000:data<=16'd1178;
      85001:data<=-16'd94;
      85002:data<=-16'd375;
      85003:data<=-16'd669;
      85004:data<=-16'd1280;
      85005:data<=-16'd735;
      85006:data<=-16'd1061;
      85007:data<=-16'd3394;
      85008:data<=-16'd3087;
      85009:data<=-16'd3630;
      85010:data<=-16'd11433;
      85011:data<=-16'd17653;
      85012:data<=-16'd17423;
      85013:data<=-16'd18265;
      85014:data<=-16'd18841;
      85015:data<=-16'd16803;
      85016:data<=-16'd16224;
      85017:data<=-16'd15811;
      85018:data<=-16'd15696;
      85019:data<=-16'd17361;
      85020:data<=-16'd17196;
      85021:data<=-16'd15993;
      85022:data<=-16'd15561;
      85023:data<=-16'd14380;
      85024:data<=-16'd14361;
      85025:data<=-16'd15614;
      85026:data<=-16'd15716;
      85027:data<=-16'd15339;
      85028:data<=-16'd14888;
      85029:data<=-16'd14066;
      85030:data<=-16'd13198;
      85031:data<=-16'd13244;
      85032:data<=-16'd14499;
      85033:data<=-16'd14566;
      85034:data<=-16'd13653;
      85035:data<=-16'd13022;
      85036:data<=-16'd11617;
      85037:data<=-16'd12222;
      85038:data<=-16'd14242;
      85039:data<=-16'd13209;
      85040:data<=-16'd13596;
      85041:data<=-16'd16662;
      85042:data<=-16'd16402;
      85043:data<=-16'd15333;
      85044:data<=-16'd16146;
      85045:data<=-16'd15420;
      85046:data<=-16'd14190;
      85047:data<=-16'd14515;
      85048:data<=-16'd14051;
      85049:data<=-16'd12380;
      85050:data<=-16'd13176;
      85051:data<=-16'd13775;
      85052:data<=-16'd6619;
      85053:data<=16'd2109;
      85054:data<=16'd3488;
      85055:data<=16'd3145;
      85056:data<=16'd2763;
      85057:data<=-16'd100;
      85058:data<=-16'd365;
      85059:data<=16'd805;
      85060:data<=16'd526;
      85061:data<=16'd1327;
      85062:data<=16'd738;
      85063:data<=-16'd861;
      85064:data<=-16'd294;
      85065:data<=-16'd640;
      85066:data<=-16'd1284;
      85067:data<=-16'd368;
      85068:data<=-16'd646;
      85069:data<=-16'd1532;
      85070:data<=-16'd1838;
      85071:data<=-16'd2053;
      85072:data<=-16'd1756;
      85073:data<=-16'd1579;
      85074:data<=-16'd1354;
      85075:data<=-16'd945;
      85076:data<=-16'd1025;
      85077:data<=-16'd836;
      85078:data<=-16'd422;
      85079:data<=-16'd9;
      85080:data<=16'd335;
      85081:data<=16'd766;
      85082:data<=16'd2488;
      85083:data<=16'd3410;
      85084:data<=16'd2899;
      85085:data<=16'd3168;
      85086:data<=16'd2422;
      85087:data<=16'd2522;
      85088:data<=16'd4987;
      85089:data<=16'd5049;
      85090:data<=16'd5465;
      85091:data<=16'd8009;
      85092:data<=16'd8605;
      85093:data<=16'd9094;
      85094:data<=16'd5483;
      85095:data<=-16'd3704;
      85096:data<=-16'd6607;
      85097:data<=-16'd4256;
      85098:data<=-16'd4140;
      85099:data<=-16'd3269;
      85100:data<=-16'd2043;
      85101:data<=-16'd1571;
      85102:data<=-16'd905;
      85103:data<=-16'd1286;
      85104:data<=-16'd1245;
      85105:data<=-16'd1387;
      85106:data<=-16'd1080;
      85107:data<=16'd1692;
      85108:data<=16'd2005;
      85109:data<=16'd957;
      85110:data<=16'd2062;
      85111:data<=16'd1680;
      85112:data<=16'd2190;
      85113:data<=16'd4200;
      85114:data<=16'd3811;
      85115:data<=16'd4194;
      85116:data<=16'd4769;
      85117:data<=16'd3698;
      85118:data<=16'd4179;
      85119:data<=16'd4975;
      85120:data<=16'd5303;
      85121:data<=16'd5598;
      85122:data<=16'd5046;
      85123:data<=16'd4819;
      85124:data<=16'd3962;
      85125:data<=16'd4184;
      85126:data<=16'd6564;
      85127:data<=16'd6475;
      85128:data<=16'd6222;
      85129:data<=16'd6833;
      85130:data<=16'd5457;
      85131:data<=16'd6346;
      85132:data<=16'd7759;
      85133:data<=16'd7210;
      85134:data<=16'd7262;
      85135:data<=16'd5594;
      85136:data<=16'd9456;
      85137:data<=16'd20682;
      85138:data<=16'd23730;
      85139:data<=16'd21387;
      85140:data<=16'd20988;
      85141:data<=16'd16601;
      85142:data<=16'd13609;
      85143:data<=16'd14566;
      85144:data<=16'd14114;
      85145:data<=16'd15001;
      85146:data<=16'd15329;
      85147:data<=16'd13858;
      85148:data<=16'd13517;
      85149:data<=16'd11775;
      85150:data<=16'd11706;
      85151:data<=16'd13923;
      85152:data<=16'd12831;
      85153:data<=16'd11803;
      85154:data<=16'd11812;
      85155:data<=16'd10766;
      85156:data<=16'd11597;
      85157:data<=16'd12114;
      85158:data<=16'd10968;
      85159:data<=16'd10804;
      85160:data<=16'd10674;
      85161:data<=16'd10308;
      85162:data<=16'd10006;
      85163:data<=16'd10217;
      85164:data<=16'd10951;
      85165:data<=16'd10202;
      85166:data<=16'd9559;
      85167:data<=16'd9288;
      85168:data<=16'd8428;
      85169:data<=16'd9406;
      85170:data<=16'd9608;
      85171:data<=16'd8120;
      85172:data<=16'd7840;
      85173:data<=16'd7042;
      85174:data<=16'd7289;
      85175:data<=16'd7465;
      85176:data<=16'd5560;
      85177:data<=16'd6813;
      85178:data<=16'd3287;
      85179:data<=-16'd8211;
      85180:data<=-16'd11265;
      85181:data<=-16'd9398;
      85182:data<=-16'd12276;
      85183:data<=-16'd12060;
      85184:data<=-16'd10511;
      85185:data<=-16'd11418;
      85186:data<=-16'd11215;
      85187:data<=-16'd11756;
      85188:data<=-16'd12460;
      85189:data<=-16'd12680;
      85190:data<=-16'd12234;
      85191:data<=-16'd8746;
      85192:data<=-16'd7259;
      85193:data<=-16'd7975;
      85194:data<=-16'd7257;
      85195:data<=-16'd8663;
      85196:data<=-16'd9242;
      85197:data<=-16'd7808;
      85198:data<=-16'd8419;
      85199:data<=-16'd7605;
      85200:data<=-16'd7585;
      85201:data<=-16'd10392;
      85202:data<=-16'd10199;
      85203:data<=-16'd9453;
      85204:data<=-16'd9556;
      85205:data<=-16'd8543;
      85206:data<=-16'd9486;
      85207:data<=-16'd10537;
      85208:data<=-16'd10404;
      85209:data<=-16'd10818;
      85210:data<=-16'd10451;
      85211:data<=-16'd10317;
      85212:data<=-16'd10053;
      85213:data<=-16'd9694;
      85214:data<=-16'd10569;
      85215:data<=-16'd9950;
      85216:data<=-16'd9776;
      85217:data<=-16'd9749;
      85218:data<=-16'd8214;
      85219:data<=-16'd10998;
      85220:data<=-16'd9186;
      85221:data<=16'd2626;
      85222:data<=16'd6669;
      85223:data<=16'd4062;
      85224:data<=16'd5128;
      85225:data<=16'd3078;
      85226:data<=16'd472;
      85227:data<=16'd1441;
      85228:data<=16'd1078;
      85229:data<=16'd1210;
      85230:data<=16'd1633;
      85231:data<=16'd569;
      85232:data<=-16'd256;
      85233:data<=-16'd1506;
      85234:data<=-16'd1377;
      85235:data<=-16'd426;
      85236:data<=-16'd930;
      85237:data<=-16'd1030;
      85238:data<=-16'd2487;
      85239:data<=-16'd3877;
      85240:data<=-16'd2892;
      85241:data<=-16'd4833;
      85242:data<=-16'd7309;
      85243:data<=-16'd6473;
      85244:data<=-16'd6852;
      85245:data<=-16'd7818;
      85246:data<=-16'd7545;
      85247:data<=-16'd7388;
      85248:data<=-16'd7080;
      85249:data<=-16'd7103;
      85250:data<=-16'd7071;
      85251:data<=-16'd7321;
      85252:data<=-16'd7694;
      85253:data<=-16'd6731;
      85254:data<=-16'd7210;
      85255:data<=-16'd7962;
      85256:data<=-16'd7259;
      85257:data<=-16'd8399;
      85258:data<=-16'd8116;
      85259:data<=-16'd7206;
      85260:data<=-16'd8216;
      85261:data<=-16'd5457;
      85262:data<=-16'd8332;
      85263:data<=-16'd21235;
      85264:data<=-16'd25358;
      85265:data<=-16'd21969;
      85266:data<=-16'd22395;
      85267:data<=-16'd20932;
      85268:data<=-16'd18891;
      85269:data<=-16'd19682;
      85270:data<=-16'd19277;
      85271:data<=-16'd18679;
      85272:data<=-16'd18295;
      85273:data<=-16'd17901;
      85274:data<=-16'd17491;
      85275:data<=-16'd15567;
      85276:data<=-16'd15085;
      85277:data<=-16'd15048;
      85278:data<=-16'd13186;
      85279:data<=-16'd12907;
      85280:data<=-16'd12443;
      85281:data<=-16'd10909;
      85282:data<=-16'd10346;
      85283:data<=-16'd8708;
      85284:data<=-16'd7752;
      85285:data<=-16'd7746;
      85286:data<=-16'd6936;
      85287:data<=-16'd7468;
      85288:data<=-16'd6131;
      85289:data<=-16'd3503;
      85290:data<=-16'd3935;
      85291:data<=-16'd2038;
      85292:data<=16'd1231;
      85293:data<=16'd972;
      85294:data<=16'd1811;
      85295:data<=16'd3891;
      85296:data<=16'd4373;
      85297:data<=16'd4285;
      85298:data<=16'd4199;
      85299:data<=16'd4576;
      85300:data<=16'd4528;
      85301:data<=16'd6178;
      85302:data<=16'd8069;
      85303:data<=16'd4913;
      85304:data<=16'd8190;
      85305:data<=16'd20466;
      85306:data<=16'd23434;
      85307:data<=16'd20980;
      85308:data<=16'd22711;
      85309:data<=16'd21106;
      85310:data<=16'd19341;
      85311:data<=16'd20280;
      85312:data<=16'd18956;
      85313:data<=16'd19215;
      85314:data<=16'd20548;
      85315:data<=16'd19919;
      85316:data<=16'd19769;
      85317:data<=16'd18742;
      85318:data<=16'd17747;
      85319:data<=16'd18398;
      85320:data<=16'd18239;
      85321:data<=16'd17785;
      85322:data<=16'd17324;
      85323:data<=16'd16877;
      85324:data<=16'd16906;
      85325:data<=16'd16407;
      85326:data<=16'd16923;
      85327:data<=16'd17479;
      85328:data<=16'd16645;
      85329:data<=16'd16603;
      85330:data<=16'd15531;
      85331:data<=16'd14302;
      85332:data<=16'd15620;
      85333:data<=16'd15867;
      85334:data<=16'd15006;
      85335:data<=16'd14298;
      85336:data<=16'd13317;
      85337:data<=16'd13706;
      85338:data<=16'd13330;
      85339:data<=16'd13103;
      85340:data<=16'd14017;
      85341:data<=16'd11189;
      85342:data<=16'd8358;
      85343:data<=16'd7553;
      85344:data<=16'd6589;
      85345:data<=16'd9432;
      85346:data<=16'd6664;
      85347:data<=-16'd5307;
      85348:data<=-16'd8942;
      85349:data<=-16'd6613;
      85350:data<=-16'd7609;
      85351:data<=-16'd5629;
      85352:data<=-16'd3808;
      85353:data<=-16'd4681;
      85354:data<=-16'd4052;
      85355:data<=-16'd4640;
      85356:data<=-16'd4821;
      85357:data<=-16'd3287;
      85358:data<=-16'd2987;
      85359:data<=-16'd2443;
      85360:data<=-16'd2540;
      85361:data<=-16'd2884;
      85362:data<=-16'd1965;
      85363:data<=-16'd1926;
      85364:data<=-16'd972;
      85365:data<=-16'd434;
      85366:data<=-16'd1803;
      85367:data<=-16'd813;
      85368:data<=-16'd381;
      85369:data<=-16'd996;
      85370:data<=16'd933;
      85371:data<=16'd1145;
      85372:data<=16'd493;
      85373:data<=16'd1192;
      85374:data<=16'd482;
      85375:data<=16'd352;
      85376:data<=16'd314;
      85377:data<=-16'd80;
      85378:data<=16'd784;
      85379:data<=16'd27;
      85380:data<=16'd0;
      85381:data<=16'd1099;
      85382:data<=-16'd517;
      85383:data<=-16'd1419;
      85384:data<=-16'd1912;
      85385:data<=-16'd1855;
      85386:data<=-16'd329;
      85387:data<=-16'd2843;
      85388:data<=-16'd422;
      85389:data<=16'd10038;
      85390:data<=16'd12131;
      85391:data<=16'd10980;
      85392:data<=16'd14868;
      85393:data<=16'd14293;
      85394:data<=16'd12040;
      85395:data<=16'd11700;
      85396:data<=16'd9940;
      85397:data<=16'd9723;
      85398:data<=16'd9533;
      85399:data<=16'd8719;
      85400:data<=16'd9028;
      85401:data<=16'd7241;
      85402:data<=16'd5591;
      85403:data<=16'd5673;
      85404:data<=16'd5206;
      85405:data<=16'd5409;
      85406:data<=16'd5147;
      85407:data<=16'd3983;
      85408:data<=16'd2896;
      85409:data<=16'd1563;
      85410:data<=16'd1750;
      85411:data<=16'd1718;
      85412:data<=16'd873;
      85413:data<=16'd1001;
      85414:data<=-16'd459;
      85415:data<=-16'd1121;
      85416:data<=-16'd179;
      85417:data<=-16'd1337;
      85418:data<=-16'd1027;
      85419:data<=-16'd681;
      85420:data<=-16'd2945;
      85421:data<=-16'd3181;
      85422:data<=-16'd3500;
      85423:data<=-16'd4117;
      85424:data<=-16'd3175;
      85425:data<=-16'd4203;
      85426:data<=-16'd4598;
      85427:data<=-16'd5309;
      85428:data<=-16'd7051;
      85429:data<=-16'd4331;
      85430:data<=-16'd7300;
      85431:data<=-16'd18359;
      85432:data<=-16'd22092;
      85433:data<=-16'd21334;
      85434:data<=-16'd21951;
      85435:data<=-16'd20365;
      85436:data<=-16'd19669;
      85437:data<=-16'd19193;
      85438:data<=-16'd18569;
      85439:data<=-16'd19992;
      85440:data<=-16'd19055;
      85441:data<=-16'd18798;
      85442:data<=-16'd21695;
      85443:data<=-16'd21531;
      85444:data<=-16'd20530;
      85445:data<=-16'd21079;
      85446:data<=-16'd20512;
      85447:data<=-16'd19937;
      85448:data<=-16'd19258;
      85449:data<=-16'd18600;
      85450:data<=-16'd18351;
      85451:data<=-16'd17681;
      85452:data<=-16'd18066;
      85453:data<=-16'd17652;
      85454:data<=-16'd15899;
      85455:data<=-16'd15819;
      85456:data<=-16'd15138;
      85457:data<=-16'd14269;
      85458:data<=-16'd15177;
      85459:data<=-16'd14828;
      85460:data<=-16'd14230;
      85461:data<=-16'd14055;
      85462:data<=-16'd12781;
      85463:data<=-16'd12578;
      85464:data<=-16'd12747;
      85465:data<=-16'd12384;
      85466:data<=-16'd11964;
      85467:data<=-16'd10492;
      85468:data<=-16'd10346;
      85469:data<=-16'd10381;
      85470:data<=-16'd9535;
      85471:data<=-16'd11218;
      85472:data<=-16'd7435;
      85473:data<=16'd3903;
      85474:data<=16'd8160;
      85475:data<=16'd6203;
      85476:data<=16'd7016;
      85477:data<=16'd7268;
      85478:data<=16'd6630;
      85479:data<=16'd7122;
      85480:data<=16'd6922;
      85481:data<=16'd6693;
      85482:data<=16'd7277;
      85483:data<=16'd8560;
      85484:data<=16'd9273;
      85485:data<=16'd8754;
      85486:data<=16'd8671;
      85487:data<=16'd7961;
      85488:data<=16'd7917;
      85489:data<=16'd10157;
      85490:data<=16'd10210;
      85491:data<=16'd10495;
      85492:data<=16'd13969;
      85493:data<=16'd14357;
      85494:data<=16'd13206;
      85495:data<=16'd14650;
      85496:data<=16'd14913;
      85497:data<=16'd13961;
      85498:data<=16'd13577;
      85499:data<=16'd12969;
      85500:data<=16'd12502;
      85501:data<=16'd12847;
      85502:data<=16'd14040;
      85503:data<=16'd13823;
      85504:data<=16'd12618;
      85505:data<=16'd12807;
      85506:data<=16'd11800;
      85507:data<=16'd11379;
      85508:data<=16'd13069;
      85509:data<=16'd12052;
      85510:data<=16'd11744;
      85511:data<=16'd12721;
      85512:data<=16'd10854;
      85513:data<=16'd11925;
      85514:data<=16'd10677;
      85515:data<=16'd572;
      85516:data<=-16'd4452;
      85517:data<=-16'd2746;
      85518:data<=-16'd3664;
      85519:data<=-16'd3278;
      85520:data<=-16'd1243;
      85521:data<=-16'd1007;
      85522:data<=-16'd1093;
      85523:data<=-16'd1454;
      85524:data<=-16'd1034;
      85525:data<=-16'd431;
      85526:data<=-16'd132;
      85527:data<=16'd1783;
      85528:data<=16'd2272;
      85529:data<=16'd1512;
      85530:data<=16'd2068;
      85531:data<=16'd1363;
      85532:data<=16'd1497;
      85533:data<=16'd3369;
      85534:data<=16'd3351;
      85535:data<=16'd3216;
      85536:data<=16'd3221;
      85537:data<=16'd2826;
      85538:data<=16'd3827;
      85539:data<=16'd4485;
      85540:data<=16'd5086;
      85541:data<=16'd5030;
      85542:data<=16'd1989;
      85543:data<=16'd143;
      85544:data<=16'd623;
      85545:data<=16'd1168;
      85546:data<=16'd2308;
      85547:data<=16'd2300;
      85548:data<=16'd1953;
      85549:data<=16'd2308;
      85550:data<=16'd1783;
      85551:data<=16'd2748;
      85552:data<=16'd3827;
      85553:data<=16'd3712;
      85554:data<=16'd4821;
      85555:data<=16'd3660;
      85556:data<=16'd5100;
      85557:data<=16'd15183;
      85558:data<=16'd21384;
      85559:data<=16'd19923;
      85560:data<=16'd19415;
      85561:data<=16'd18365;
      85562:data<=16'd16525;
      85563:data<=16'd16863;
      85564:data<=16'd17613;
      85565:data<=16'd17705;
      85566:data<=16'd16521;
      85567:data<=16'd15512;
      85568:data<=16'd15482;
      85569:data<=16'd14311;
      85570:data<=16'd14126;
      85571:data<=16'd14879;
      85572:data<=16'd14055;
      85573:data<=16'd13775;
      85574:data<=16'd13430;
      85575:data<=16'd12328;
      85576:data<=16'd12141;
      85577:data<=16'd11295;
      85578:data<=16'd10408;
      85579:data<=16'd10188;
      85580:data<=16'd9226;
      85581:data<=16'd8805;
      85582:data<=16'd7985;
      85583:data<=16'd5952;
      85584:data<=16'd4795;
      85585:data<=16'd4356;
      85586:data<=16'd4514;
      85587:data<=16'd4402;
      85588:data<=16'd3495;
      85589:data<=16'd2940;
      85590:data<=16'd1171;
      85591:data<=16'd526;
      85592:data<=16'd2934;
      85593:data<=16'd3670;
      85594:data<=16'd3780;
      85595:data<=16'd3410;
      85596:data<=16'd614;
      85597:data<=16'd1068;
      85598:data<=-16'd591;
      85599:data<=-16'd10470;
      85600:data<=-16'd15864;
      85601:data<=-16'd15045;
      85602:data<=-16'd16578;
      85603:data<=-16'd16725;
      85604:data<=-16'd15346;
      85605:data<=-16'd15840;
      85606:data<=-16'd15358;
      85607:data<=-16'd15010;
      85608:data<=-16'd16116;
      85609:data<=-16'd16111;
      85610:data<=-16'd15191;
      85611:data<=-16'd14483;
      85612:data<=-16'd14114;
      85613:data<=-16'd13969;
      85614:data<=-16'd14236;
      85615:data<=-16'd14991;
      85616:data<=-16'd14777;
      85617:data<=-16'd14164;
      85618:data<=-16'd14176;
      85619:data<=-16'd13336;
      85620:data<=-16'd12986;
      85621:data<=-16'd14076;
      85622:data<=-16'd14075;
      85623:data<=-16'd13524;
      85624:data<=-16'd13286;
      85625:data<=-16'd12258;
      85626:data<=-16'd12049;
      85627:data<=-16'd13367;
      85628:data<=-16'd14181;
      85629:data<=-16'd13899;
      85630:data<=-16'd13054;
      85631:data<=-16'd12120;
      85632:data<=-16'd11913;
      85633:data<=-16'd12812;
      85634:data<=-16'd13018;
      85635:data<=-16'd11606;
      85636:data<=-16'd11527;
      85637:data<=-16'd11765;
      85638:data<=-16'd10202;
      85639:data<=-16'd11458;
      85640:data<=-16'd11148;
      85641:data<=-16'd2100;
      85642:data<=16'd3412;
      85643:data<=-16'd9;
      85644:data<=-16'd523;
      85645:data<=16'd256;
      85646:data<=-16'd2188;
      85647:data<=-16'd2362;
      85648:data<=-16'd1776;
      85649:data<=-16'd2065;
      85650:data<=-16'd1148;
      85651:data<=-16'd1754;
      85652:data<=-16'd3236;
      85653:data<=-16'd3336;
      85654:data<=-16'd3145;
      85655:data<=-16'd2617;
      85656:data<=-16'd2722;
      85657:data<=-16'd3269;
      85658:data<=-16'd3322;
      85659:data<=-16'd4275;
      85660:data<=-16'd4654;
      85661:data<=-16'd4262;
      85662:data<=-16'd4616;
      85663:data<=-16'd3971;
      85664:data<=-16'd4137;
      85665:data<=-16'd6017;
      85666:data<=-16'd6111;
      85667:data<=-16'd5683;
      85668:data<=-16'd5541;
      85669:data<=-16'd4464;
      85670:data<=-16'd4739;
      85671:data<=-16'd5952;
      85672:data<=-16'd5991;
      85673:data<=-16'd5547;
      85674:data<=-16'd5254;
      85675:data<=-16'd5285;
      85676:data<=-16'd5518;
      85677:data<=-16'd5689;
      85678:data<=-16'd4934;
      85679:data<=-16'd3630;
      85680:data<=-16'd3844;
      85681:data<=-16'd3635;
      85682:data<=-16'd4323;
      85683:data<=-16'd10944;
      85684:data<=-16'd16857;
      85685:data<=-16'd16298;
      85686:data<=-16'd14983;
      85687:data<=-16'd14794;
      85688:data<=-16'd14430;
      85689:data<=-16'd13129;
      85690:data<=-16'd10851;
      85691:data<=-16'd10716;
      85692:data<=-16'd9265;
      85693:data<=-16'd4977;
      85694:data<=-16'd4617;
      85695:data<=-16'd4763;
      85696:data<=-16'd2137;
      85697:data<=-16'd1865;
      85698:data<=-16'd1574;
      85699:data<=-16'd634;
      85700:data<=-16'd1718;
      85701:data<=-16'd861;
      85702:data<=16'd1292;
      85703:data<=16'd1767;
      85704:data<=16'd1949;
      85705:data<=16'd1789;
      85706:data<=16'd1970;
      85707:data<=16'd2572;
      85708:data<=16'd2966;
      85709:data<=16'd4040;
      85710:data<=16'd4043;
      85711:data<=16'd3577;
      85712:data<=16'd4109;
      85713:data<=16'd3415;
      85714:data<=16'd3698;
      85715:data<=16'd5770;
      85716:data<=16'd6241;
      85717:data<=16'd6558;
      85718:data<=16'd6748;
      85719:data<=16'd5821;
      85720:data<=16'd5968;
      85721:data<=16'd6693;
      85722:data<=16'd7489;
      85723:data<=16'd7374;
      85724:data<=16'd7394;
      85725:data<=16'd13899;
      85726:data<=16'd22309;
      85727:data<=16'd23837;
      85728:data<=16'd22980;
      85729:data<=16'd22656;
      85730:data<=16'd21325;
      85731:data<=16'd20701;
      85732:data<=16'd19826;
      85733:data<=16'd19567;
      85734:data<=16'd21161;
      85735:data<=16'd20947;
      85736:data<=16'd19473;
      85737:data<=16'd18735;
      85738:data<=16'd17672;
      85739:data<=16'd17249;
      85740:data<=16'd17893;
      85741:data<=16'd18407;
      85742:data<=16'd16775;
      85743:data<=16'd12592;
      85744:data<=16'd10505;
      85745:data<=16'd11491;
      85746:data<=16'd11991;
      85747:data<=16'd11928;
      85748:data<=16'd11348;
      85749:data<=16'd10466;
      85750:data<=16'd10395;
      85751:data<=16'd10395;
      85752:data<=16'd11047;
      85753:data<=16'd11544;
      85754:data<=16'd10481;
      85755:data<=16'd10222;
      85756:data<=16'd9922;
      85757:data<=16'd8531;
      85758:data<=16'd9031;
      85759:data<=16'd10072;
      85760:data<=16'd9629;
      85761:data<=16'd9104;
      85762:data<=16'd8658;
      85763:data<=16'd8252;
      85764:data<=16'd8073;
      85765:data<=16'd9065;
      85766:data<=16'd9445;
      85767:data<=16'd3318;
      85768:data<=-16'd5098;
      85769:data<=-16'd6499;
      85770:data<=-16'd4259;
      85771:data<=-16'd3571;
      85772:data<=-16'd3118;
      85773:data<=-16'd2695;
      85774:data<=-16'd2632;
      85775:data<=-16'd2914;
      85776:data<=-16'd3113;
      85777:data<=-16'd2767;
      85778:data<=-16'd2921;
      85779:data<=-16'd2874;
      85780:data<=-16'd2822;
      85781:data<=-16'd3830;
      85782:data<=-16'd3767;
      85783:data<=-16'd3889;
      85784:data<=-16'd5730;
      85785:data<=-16'd6044;
      85786:data<=-16'd5597;
      85787:data<=-16'd5805;
      85788:data<=-16'd5168;
      85789:data<=-16'd5195;
      85790:data<=-16'd6278;
      85791:data<=-16'd6848;
      85792:data<=-16'd5882;
      85793:data<=-16'd2937;
      85794:data<=-16'd1513;
      85795:data<=-16'd2802;
      85796:data<=-16'd3836;
      85797:data<=-16'd4561;
      85798:data<=-16'd4487;
      85799:data<=-16'd3753;
      85800:data<=-16'd3900;
      85801:data<=-16'd3626;
      85802:data<=-16'd4099;
      85803:data<=-16'd5250;
      85804:data<=-16'd4951;
      85805:data<=-16'd5880;
      85806:data<=-16'd5897;
      85807:data<=-16'd4266;
      85808:data<=-16'd6078;
      85809:data<=-16'd3336;
      85810:data<=16'd6053;
      85811:data<=16'd8091;
      85812:data<=16'd5732;
      85813:data<=16'd6896;
      85814:data<=16'd5609;
      85815:data<=16'd3231;
      85816:data<=16'd3650;
      85817:data<=16'd3500;
      85818:data<=16'd3357;
      85819:data<=16'd3703;
      85820:data<=16'd2485;
      85821:data<=16'd758;
      85822:data<=16'd133;
      85823:data<=16'd469;
      85824:data<=16'd55;
      85825:data<=-16'd617;
      85826:data<=-16'd68;
      85827:data<=-16'd987;
      85828:data<=-16'd3106;
      85829:data<=-16'd3298;
      85830:data<=-16'd3225;
      85831:data<=-16'd3362;
      85832:data<=-16'd2754;
      85833:data<=-16'd3457;
      85834:data<=-16'd4775;
      85835:data<=-16'd4504;
      85836:data<=-16'd3891;
      85837:data<=-16'd3782;
      85838:data<=-16'd3271;
      85839:data<=-16'd3485;
      85840:data<=-16'd5062;
      85841:data<=-16'd5385;
      85842:data<=-16'd5783;
      85843:data<=-16'd8745;
      85844:data<=-16'd9770;
      85845:data<=-16'd8980;
      85846:data<=-16'd10520;
      85847:data<=-16'd10825;
      85848:data<=-16'd9997;
      85849:data<=-16'd10091;
      85850:data<=-16'd8431;
      85851:data<=-16'd11611;
      85852:data<=-16'd21288;
      85853:data<=-16'd24692;
      85854:data<=-16'd22193;
      85855:data<=-16'd21755;
      85856:data<=-16'd21088;
      85857:data<=-16'd19754;
      85858:data<=-16'd19782;
      85859:data<=-16'd20158;
      85860:data<=-16'd20274;
      85861:data<=-16'd19415;
      85862:data<=-16'd18298;
      85863:data<=-16'd17411;
      85864:data<=-16'd16718;
      85865:data<=-16'd17587;
      85866:data<=-16'd17562;
      85867:data<=-16'd16076;
      85868:data<=-16'd16249;
      85869:data<=-16'd15491;
      85870:data<=-16'd13905;
      85871:data<=-16'd14643;
      85872:data<=-16'd14471;
      85873:data<=-16'd13211;
      85874:data<=-16'd12927;
      85875:data<=-16'd11923;
      85876:data<=-16'd11295;
      85877:data<=-16'd11307;
      85878:data<=-16'd10477;
      85879:data<=-16'd9868;
      85880:data<=-16'd9092;
      85881:data<=-16'd8366;
      85882:data<=-16'd8423;
      85883:data<=-16'd7244;
      85884:data<=-16'd4933;
      85885:data<=-16'd3656;
      85886:data<=-16'd3748;
      85887:data<=-16'd3489;
      85888:data<=-16'd2704;
      85889:data<=-16'd2690;
      85890:data<=-16'd817;
      85891:data<=16'd749;
      85892:data<=-16'd883;
      85893:data<=16'd5348;
      85894:data<=16'd17584;
      85895:data<=16'd19490;
      85896:data<=16'd17523;
      85897:data<=16'd19711;
      85898:data<=16'd18700;
      85899:data<=16'd17417;
      85900:data<=16'd18013;
      85901:data<=16'd16383;
      85902:data<=16'd16686;
      85903:data<=16'd18433;
      85904:data<=16'd17832;
      85905:data<=16'd17224;
      85906:data<=16'd16651;
      85907:data<=16'd16010;
      85908:data<=16'd16349;
      85909:data<=16'd16977;
      85910:data<=16'd17650;
      85911:data<=16'd17091;
      85912:data<=16'd15914;
      85913:data<=16'd15484;
      85914:data<=16'd14994;
      85915:data<=16'd15656;
      85916:data<=16'd16271;
      85917:data<=16'd15180;
      85918:data<=16'd15050;
      85919:data<=16'd14712;
      85920:data<=16'd13529;
      85921:data<=16'd14345;
      85922:data<=16'd15291;
      85923:data<=16'd14822;
      85924:data<=16'd13966;
      85925:data<=16'd13000;
      85926:data<=16'd12515;
      85927:data<=16'd12592;
      85928:data<=16'd13908;
      85929:data<=16'd14428;
      85930:data<=16'd12466;
      85931:data<=16'd12301;
      85932:data<=16'd12495;
      85933:data<=16'd11909;
      85934:data<=16'd14342;
      85935:data<=16'd10954;
      85936:data<=16'd466;
      85937:data<=-16'd2270;
      85938:data<=16'd55;
      85939:data<=-16'd740;
      85940:data<=-16'd6;
      85941:data<=16'd1547;
      85942:data<=16'd840;
      85943:data<=-16'd1152;
      85944:data<=-16'd3671;
      85945:data<=-16'd4059;
      85946:data<=-16'd2731;
      85947:data<=-16'd1838;
      85948:data<=-16'd1306;
      85949:data<=-16'd1756;
      85950:data<=-16'd1804;
      85951:data<=-16'd1307;
      85952:data<=-16'd1366;
      85953:data<=-16'd202;
      85954:data<=16'd537;
      85955:data<=16'd190;
      85956:data<=16'd890;
      85957:data<=16'd619;
      85958:data<=16'd534;
      85959:data<=16'd1997;
      85960:data<=16'd1706;
      85961:data<=16'd1206;
      85962:data<=16'd1539;
      85963:data<=16'd814;
      85964:data<=16'd908;
      85965:data<=16'd2091;
      85966:data<=16'd2934;
      85967:data<=16'd2980;
      85968:data<=16'd2419;
      85969:data<=16'd2732;
      85970:data<=16'd2779;
      85971:data<=16'd3016;
      85972:data<=16'd4508;
      85973:data<=16'd3891;
      85974:data<=16'd3683;
      85975:data<=16'd4537;
      85976:data<=16'd2291;
      85977:data<=16'd5504;
      85978:data<=16'd14818;
      85979:data<=16'd16604;
      85980:data<=16'd14236;
      85981:data<=16'd14604;
      85982:data<=16'd13594;
      85983:data<=16'd12258;
      85984:data<=16'd11126;
      85985:data<=16'd9259;
      85986:data<=16'd9357;
      85987:data<=16'd9007;
      85988:data<=16'd7379;
      85989:data<=16'd7262;
      85990:data<=16'd6696;
      85991:data<=16'd5022;
      85992:data<=16'd4225;
      85993:data<=16'd5418;
      85994:data<=16'd8161;
      85995:data<=16'd8878;
      85996:data<=16'd6907;
      85997:data<=16'd4977;
      85998:data<=16'd3902;
      85999:data<=16'd3950;
      86000:data<=16'd4141;
      86001:data<=16'd3656;
      86002:data<=16'd2811;
      86003:data<=16'd1180;
      86004:data<=16'd652;
      86005:data<=16'd1089;
      86006:data<=16'd133;
      86007:data<=16'd42;
      86008:data<=16'd106;
      86009:data<=-16'd1671;
      86010:data<=-16'd2220;
      86011:data<=-16'd2334;
      86012:data<=-16'd3136;
      86013:data<=-16'd2907;
      86014:data<=-16'd3025;
      86015:data<=-16'd3556;
      86016:data<=-16'd4971;
      86017:data<=-16'd6087;
      86018:data<=-16'd3852;
      86019:data<=-16'd6649;
      86020:data<=-16'd16337;
      86021:data<=-16'd19778;
      86022:data<=-16'd18604;
      86023:data<=-16'd19619;
      86024:data<=-16'd18662;
      86025:data<=-16'd17285;
      86026:data<=-16'd17578;
      86027:data<=-16'd17529;
      86028:data<=-16'd18578;
      86029:data<=-16'd18956;
      86030:data<=-16'd17814;
      86031:data<=-16'd17713;
      86032:data<=-16'd17302;
      86033:data<=-16'd16630;
      86034:data<=-16'd16888;
      86035:data<=-16'd17042;
      86036:data<=-16'd16973;
      86037:data<=-16'd16475;
      86038:data<=-16'd15729;
      86039:data<=-16'd14783;
      86040:data<=-16'd14410;
      86041:data<=-16'd15617;
      86042:data<=-16'd15400;
      86043:data<=-16'd15562;
      86044:data<=-16'd18794;
      86045:data<=-16'd18760;
      86046:data<=-16'd17170;
      86047:data<=-16'd18904;
      86048:data<=-16'd18534;
      86049:data<=-16'd17014;
      86050:data<=-16'd16888;
      86051:data<=-16'd15176;
      86052:data<=-16'd14754;
      86053:data<=-16'd15702;
      86054:data<=-16'd15379;
      86055:data<=-16'd14994;
      86056:data<=-16'd13869;
      86057:data<=-16'd13577;
      86058:data<=-16'd13605;
      86059:data<=-16'd12786;
      86060:data<=-16'd14775;
      86061:data<=-16'd11586;
      86062:data<=-16'd784;
      86063:data<=16'd2397;
      86064:data<=16'd287;
      86065:data<=16'd1381;
      86066:data<=16'd162;
      86067:data<=-16'd1054;
      86068:data<=-16'd133;
      86069:data<=-16'd946;
      86070:data<=-16'd553;
      86071:data<=-16'd45;
      86072:data<=-16'd1504;
      86073:data<=-16'd1554;
      86074:data<=-16'd1224;
      86075:data<=-16'd1395;
      86076:data<=-16'd1298;
      86077:data<=-16'd1216;
      86078:data<=-16'd227;
      86079:data<=-16'd70;
      86080:data<=-16'd767;
      86081:data<=-16'd143;
      86082:data<=16'd9;
      86083:data<=16'd79;
      86084:data<=16'd1401;
      86085:data<=16'd2153;
      86086:data<=16'd2215;
      86087:data<=16'd2259;
      86088:data<=16'd2387;
      86089:data<=16'd2340;
      86090:data<=16'd2924;
      86091:data<=16'd4895;
      86092:data<=16'd4934;
      86093:data<=16'd4899;
      86094:data<=16'd8153;
      86095:data<=16'd8849;
      86096:data<=16'd8167;
      86097:data<=16'd10290;
      86098:data<=16'd10229;
      86099:data<=16'd9627;
      86100:data<=16'd9881;
      86101:data<=16'd8436;
      86102:data<=16'd9664;
      86103:data<=16'd7997;
      86104:data<=-16'd857;
      86105:data<=-16'd4193;
      86106:data<=-16'd2118;
      86107:data<=-16'd2878;
      86108:data<=-16'd2963;
      86109:data<=-16'd1601;
      86110:data<=-16'd411;
      86111:data<=16'd663;
      86112:data<=16'd103;
      86113:data<=-16'd130;
      86114:data<=16'd402;
      86115:data<=16'd1017;
      86116:data<=16'd2826;
      86117:data<=16'd3172;
      86118:data<=16'd2343;
      86119:data<=16'd2561;
      86120:data<=16'd2200;
      86121:data<=16'd2732;
      86122:data<=16'd4528;
      86123:data<=16'd4957;
      86124:data<=16'd4842;
      86125:data<=16'd4626;
      86126:data<=16'd4387;
      86127:data<=16'd4755;
      86128:data<=16'd5483;
      86129:data<=16'd6660;
      86130:data<=16'd6407;
      86131:data<=16'd5445;
      86132:data<=16'd6144;
      86133:data<=16'd5923;
      86134:data<=16'd5979;
      86135:data<=16'd7982;
      86136:data<=16'd8067;
      86137:data<=16'd7504;
      86138:data<=16'd7705;
      86139:data<=16'd7312;
      86140:data<=16'd7909;
      86141:data<=16'd8202;
      86142:data<=16'd8341;
      86143:data<=16'd7712;
      86144:data<=16'd3110;
      86145:data<=16'd4501;
      86146:data<=16'd14945;
      86147:data<=16'd18873;
      86148:data<=16'd16600;
      86149:data<=16'd17127;
      86150:data<=16'd16774;
      86151:data<=16'd15423;
      86152:data<=16'd15556;
      86153:data<=16'd15584;
      86154:data<=16'd15855;
      86155:data<=16'd15317;
      86156:data<=16'd14082;
      86157:data<=16'd13705;
      86158:data<=16'd12974;
      86159:data<=16'd13226;
      86160:data<=16'd14360;
      86161:data<=16'd13579;
      86162:data<=16'd12965;
      86163:data<=16'd13015;
      86164:data<=16'd11585;
      86165:data<=16'd10968;
      86166:data<=16'd11973;
      86167:data<=16'd11899;
      86168:data<=16'd11075;
      86169:data<=16'd10862;
      86170:data<=16'd10176;
      86171:data<=16'd9700;
      86172:data<=16'd10831;
      86173:data<=16'd11013;
      86174:data<=16'd9747;
      86175:data<=16'd9326;
      86176:data<=16'd8701;
      86177:data<=16'd8232;
      86178:data<=16'd8241;
      86179:data<=16'd6704;
      86180:data<=16'd6135;
      86181:data<=16'd6384;
      86182:data<=16'd5051;
      86183:data<=16'd5401;
      86184:data<=16'd4849;
      86185:data<=16'd1988;
      86186:data<=16'd2663;
      86187:data<=16'd105;
      86188:data<=-16'd9213;
      86189:data<=-16'd13115;
      86190:data<=-16'd12120;
      86191:data<=-16'd13392;
      86192:data<=-16'd13846;
      86193:data<=-16'd12334;
      86194:data<=-16'd9700;
      86195:data<=-16'd7492;
      86196:data<=-16'd8476;
      86197:data<=-16'd9304;
      86198:data<=-16'd8795;
      86199:data<=-16'd9503;
      86200:data<=-16'd9659;
      86201:data<=-16'd9125;
      86202:data<=-16'd9118;
      86203:data<=-16'd9509;
      86204:data<=-16'd10660;
      86205:data<=-16'd10605;
      86206:data<=-16'd9694;
      86207:data<=-16'd9747;
      86208:data<=-16'd9168;
      86209:data<=-16'd9389;
      86210:data<=-16'd10625;
      86211:data<=-16'd10134;
      86212:data<=-16'd10202;
      86213:data<=-16'd10583;
      86214:data<=-16'd9204;
      86215:data<=-16'd9348;
      86216:data<=-16'd10581;
      86217:data<=-16'd10272;
      86218:data<=-16'd9943;
      86219:data<=-16'd9852;
      86220:data<=-16'd9113;
      86221:data<=-16'd8654;
      86222:data<=-16'd9771;
      86223:data<=-16'd10781;
      86224:data<=-16'd9852;
      86225:data<=-16'd10002;
      86226:data<=-16'd10213;
      86227:data<=-16'd8639;
      86228:data<=-16'd10220;
      86229:data<=-16'd9323;
      86230:data<=-16'd349;
      86231:data<=16'd4034;
      86232:data<=16'd1965;
      86233:data<=16'd2775;
      86234:data<=16'd2681;
      86235:data<=16'd734;
      86236:data<=16'd1048;
      86237:data<=16'd482;
      86238:data<=-16'd423;
      86239:data<=16'd294;
      86240:data<=-16'd215;
      86241:data<=-16'd1469;
      86242:data<=-16'd1704;
      86243:data<=-16'd2384;
      86244:data<=-16'd4625;
      86245:data<=-16'd6097;
      86246:data<=-16'd5281;
      86247:data<=-16'd5756;
      86248:data<=-16'd7645;
      86249:data<=-16'd7204;
      86250:data<=-16'd6240;
      86251:data<=-16'd6304;
      86252:data<=-16'd5839;
      86253:data<=-16'd5858;
      86254:data<=-16'd6727;
      86255:data<=-16'd7262;
      86256:data<=-16'd7272;
      86257:data<=-16'd6839;
      86258:data<=-16'd6237;
      86259:data<=-16'd6247;
      86260:data<=-16'd7689;
      86261:data<=-16'd8514;
      86262:data<=-16'd7233;
      86263:data<=-16'd6643;
      86264:data<=-16'd6370;
      86265:data<=-16'd5990;
      86266:data<=-16'd7682;
      86267:data<=-16'd7790;
      86268:data<=-16'd6479;
      86269:data<=-16'd7141;
      86270:data<=-16'd5796;
      86271:data<=-16'd7042;
      86272:data<=-16'd15902;
      86273:data<=-16'd21123;
      86274:data<=-16'd20048;
      86275:data<=-16'd19660;
      86276:data<=-16'd18847;
      86277:data<=-16'd17978;
      86278:data<=-16'd17432;
      86279:data<=-16'd15446;
      86280:data<=-16'd14795;
      86281:data<=-16'd14404;
      86282:data<=-16'd12757;
      86283:data<=-16'd12493;
      86284:data<=-16'd11450;
      86285:data<=-16'd9189;
      86286:data<=-16'd8636;
      86287:data<=-16'd8103;
      86288:data<=-16'd7194;
      86289:data<=-16'd7022;
      86290:data<=-16'd6012;
      86291:data<=-16'd4220;
      86292:data<=-16'd3005;
      86293:data<=-16'd1906;
      86294:data<=16'd481;
      86295:data<=16'd2943;
      86296:data<=16'd2945;
      86297:data<=16'd2949;
      86298:data<=16'd4918;
      86299:data<=16'd5542;
      86300:data<=16'd4993;
      86301:data<=16'd5407;
      86302:data<=16'd5274;
      86303:data<=16'd5118;
      86304:data<=16'd6743;
      86305:data<=16'd7953;
      86306:data<=16'd7233;
      86307:data<=16'd6989;
      86308:data<=16'd7586;
      86309:data<=16'd7468;
      86310:data<=16'd8627;
      86311:data<=16'd10134;
      86312:data<=16'd8352;
      86313:data<=16'd9307;
      86314:data<=16'd17138;
      86315:data<=16'd22848;
      86316:data<=16'd23205;
      86317:data<=16'd23212;
      86318:data<=16'd22641;
      86319:data<=16'd21640;
      86320:data<=16'd21452;
      86321:data<=16'd20186;
      86322:data<=16'd19469;
      86323:data<=16'd20692;
      86324:data<=16'd20941;
      86325:data<=16'd20436;
      86326:data<=16'd20072;
      86327:data<=16'd18860;
      86328:data<=16'd18707;
      86329:data<=16'd20051;
      86330:data<=16'd20263;
      86331:data<=16'd19390;
      86332:data<=16'd18383;
      86333:data<=16'd17552;
      86334:data<=16'd17766;
      86335:data<=16'd18240;
      86336:data<=16'd17893;
      86337:data<=16'd17312;
      86338:data<=16'd16768;
      86339:data<=16'd16143;
      86340:data<=16'd15487;
      86341:data<=16'd15182;
      86342:data<=16'd15716;
      86343:data<=16'd15438;
      86344:data<=16'd12844;
      86345:data<=16'd9967;
      86346:data<=16'd8849;
      86347:data<=16'd9401;
      86348:data<=16'd10693;
      86349:data<=16'd10781;
      86350:data<=16'd9558;
      86351:data<=16'd9174;
      86352:data<=16'd9001;
      86353:data<=16'd8740;
      86354:data<=16'd10434;
      86355:data<=16'd9720;
      86356:data<=16'd2014;
      86357:data<=-16'd5157;
      86358:data<=-16'd5589;
      86359:data<=-16'd3879;
      86360:data<=-16'd2933;
      86361:data<=-16'd2278;
      86362:data<=-16'd2588;
      86363:data<=-16'd2799;
      86364:data<=-16'd2529;
      86365:data<=-16'd2446;
      86366:data<=-16'd1521;
      86367:data<=-16'd470;
      86368:data<=-16'd519;
      86369:data<=-16'd419;
      86370:data<=-16'd23;
      86371:data<=-16'd393;
      86372:data<=-16'd690;
      86373:data<=16'd355;
      86374:data<=16'd1425;
      86375:data<=16'd907;
      86376:data<=16'd253;
      86377:data<=16'd314;
      86378:data<=16'd65;
      86379:data<=16'd14;
      86380:data<=-16'd39;
      86381:data<=-16'd672;
      86382:data<=-16'd378;
      86383:data<=16'd256;
      86384:data<=-16'd566;
      86385:data<=-16'd1785;
      86386:data<=-16'd2393;
      86387:data<=-16'd2660;
      86388:data<=-16'd2719;
      86389:data<=-16'd3010;
      86390:data<=-16'd3586;
      86391:data<=-16'd3827;
      86392:data<=-16'd4120;
      86393:data<=-16'd5039;
      86394:data<=-16'd4276;
      86395:data<=-16'd1064;
      86396:data<=-16'd329;
      86397:data<=-16'd1330;
      86398:data<=16'd3284;
      86399:data<=16'd9956;
      86400:data<=16'd10370;
      86401:data<=16'd8395;
      86402:data<=16'd8945;
      86403:data<=16'd8658;
      86404:data<=16'd6563;
      86405:data<=16'd5495;
      86406:data<=16'd5238;
      86407:data<=16'd4664;
      86408:data<=16'd4399;
      86409:data<=16'd4002;
      86410:data<=16'd2590;
      86411:data<=16'd1394;
      86412:data<=16'd1019;
      86413:data<=16'd502;
      86414:data<=16'd411;
      86415:data<=16'd840;
      86416:data<=-16'd41;
      86417:data<=-16'd1538;
      86418:data<=-16'd1754;
      86419:data<=-16'd1970;
      86420:data<=-16'd2645;
      86421:data<=-16'd2181;
      86422:data<=-16'd2196;
      86423:data<=-16'd4084;
      86424:data<=-16'd5178;
      86425:data<=-16'd4907;
      86426:data<=-16'd4660;
      86427:data<=-16'd4038;
      86428:data<=-16'd4592;
      86429:data<=-16'd6974;
      86430:data<=-16'd7527;
      86431:data<=-16'd6381;
      86432:data<=-16'd6528;
      86433:data<=-16'd6730;
      86434:data<=-16'd6619;
      86435:data<=-16'd7652;
      86436:data<=-16'd8429;
      86437:data<=-16'd8486;
      86438:data<=-16'd8132;
      86439:data<=-16'd7773;
      86440:data<=-16'd12248;
      86441:data<=-16'd20789;
      86442:data<=-16'd23497;
      86443:data<=-16'd20768;
      86444:data<=-16'd21361;
      86445:data<=-16'd23824;
      86446:data<=-16'd23588;
      86447:data<=-16'd22571;
      86448:data<=-16'd22072;
      86449:data<=-16'd21185;
      86450:data<=-16'd20033;
      86451:data<=-16'd19176;
      86452:data<=-16'd18701;
      86453:data<=-16'd18322;
      86454:data<=-16'd18359;
      86455:data<=-16'd18554;
      86456:data<=-16'd17901;
      86457:data<=-16'd17156;
      86458:data<=-16'd16621;
      86459:data<=-16'd15559;
      86460:data<=-16'd15493;
      86461:data<=-16'd16563;
      86462:data<=-16'd16157;
      86463:data<=-16'd14897;
      86464:data<=-16'd14519;
      86465:data<=-16'd13602;
      86466:data<=-16'd12727;
      86467:data<=-16'd13738;
      86468:data<=-16'd14110;
      86469:data<=-16'd12874;
      86470:data<=-16'd12217;
      86471:data<=-16'd11392;
      86472:data<=-16'd10916;
      86473:data<=-16'd12002;
      86474:data<=-16'd12038;
      86475:data<=-16'd11191;
      86476:data<=-16'd10721;
      86477:data<=-16'd9996;
      86478:data<=-16'd10128;
      86479:data<=-16'd9283;
      86480:data<=-16'd8123;
      86481:data<=-16'd9268;
      86482:data<=-16'd4269;
      86483:data<=16'd5855;
      86484:data<=16'd7389;
      86485:data<=16'd5668;
      86486:data<=16'd8217;
      86487:data<=16'd8160;
      86488:data<=16'd7370;
      86489:data<=16'd8499;
      86490:data<=16'd7521;
      86491:data<=16'd7641;
      86492:data<=16'd9386;
      86493:data<=16'd9462;
      86494:data<=16'd10143;
      86495:data<=16'd11035;
      86496:data<=16'd10543;
      86497:data<=16'd10784;
      86498:data<=16'd12163;
      86499:data<=16'd13012;
      86500:data<=16'd12207;
      86501:data<=16'd11185;
      86502:data<=16'd11132;
      86503:data<=16'd10768;
      86504:data<=16'd11119;
      86505:data<=16'd12176;
      86506:data<=16'd11771;
      86507:data<=16'd11383;
      86508:data<=16'd11317;
      86509:data<=16'd10329;
      86510:data<=16'd10454;
      86511:data<=16'd11862;
      86512:data<=16'd12078;
      86513:data<=16'd11021;
      86514:data<=16'd10411;
      86515:data<=16'd10282;
      86516:data<=16'd10439;
      86517:data<=16'd12032;
      86518:data<=16'd12358;
      86519:data<=16'd10393;
      86520:data<=16'd10492;
      86521:data<=16'd10299;
      86522:data<=16'd9618;
      86523:data<=16'd12434;
      86524:data<=16'd8943;
      86525:data<=-16'd1527;
      86526:data<=-16'd3576;
      86527:data<=-16'd975;
      86528:data<=-16'd2188;
      86529:data<=-16'd1262;
      86530:data<=16'd996;
      86531:data<=16'd963;
      86532:data<=16'd898;
      86533:data<=16'd846;
      86534:data<=16'd1083;
      86535:data<=16'd1764;
      86536:data<=16'd2416;
      86537:data<=16'd3324;
      86538:data<=16'd3124;
      86539:data<=16'd2651;
      86540:data<=16'd2781;
      86541:data<=16'd2713;
      86542:data<=16'd3839;
      86543:data<=16'd4541;
      86544:data<=16'd3247;
      86545:data<=16'd2191;
      86546:data<=16'd1354;
      86547:data<=16'd1632;
      86548:data<=16'd2907;
      86549:data<=16'd2594;
      86550:data<=16'd2928;
      86551:data<=16'd3915;
      86552:data<=16'd2896;
      86553:data<=16'd2394;
      86554:data<=16'd3383;
      86555:data<=16'd4191;
      86556:data<=16'd4243;
      86557:data<=16'd3883;
      86558:data<=16'd3882;
      86559:data<=16'd3007;
      86560:data<=16'd3278;
      86561:data<=16'd5510;
      86562:data<=16'd4676;
      86563:data<=16'd4193;
      86564:data<=16'd5151;
      86565:data<=16'd2460;
      86566:data<=16'd6510;
      86567:data<=16'd17801;
      86568:data<=16'd19469;
      86569:data<=16'd16219;
      86570:data<=16'd16941;
      86571:data<=16'd15898;
      86572:data<=16'd14880;
      86573:data<=16'd15666;
      86574:data<=16'd15057;
      86575:data<=16'd14816;
      86576:data<=16'd14281;
      86577:data<=16'd13073;
      86578:data<=16'd12936;
      86579:data<=16'd12111;
      86580:data<=16'd10983;
      86581:data<=16'd10490;
      86582:data<=16'd9818;
      86583:data<=16'd9753;
      86584:data<=16'd9583;
      86585:data<=16'd8296;
      86586:data<=16'd6405;
      86587:data<=16'd4787;
      86588:data<=16'd4393;
      86589:data<=16'd4199;
      86590:data<=16'd4017;
      86591:data<=16'd3668;
      86592:data<=16'd1265;
      86593:data<=-16'd466;
      86594:data<=16'd638;
      86595:data<=16'd1956;
      86596:data<=16'd2655;
      86597:data<=16'd2008;
      86598:data<=16'd396;
      86599:data<=-16'd353;
      86600:data<=-16'd1071;
      86601:data<=-16'd1174;
      86602:data<=-16'd1225;
      86603:data<=-16'd2218;
      86604:data<=-16'd2038;
      86605:data<=-16'd3389;
      86606:data<=-16'd4725;
      86607:data<=-16'd2062;
      86608:data<=-16'd5749;
      86609:data<=-16'd15820;
      86610:data<=-16'd18431;
      86611:data<=-16'd17341;
      86612:data<=-16'd18384;
      86613:data<=-16'd17455;
      86614:data<=-16'd16637;
      86615:data<=-16'd16745;
      86616:data<=-16'd16307;
      86617:data<=-16'd16901;
      86618:data<=-16'd16703;
      86619:data<=-16'd15920;
      86620:data<=-16'd16190;
      86621:data<=-16'd15458;
      86622:data<=-16'd14478;
      86623:data<=-16'd14845;
      86624:data<=-16'd15602;
      86625:data<=-16'd15796;
      86626:data<=-16'd15294;
      86627:data<=-16'd14780;
      86628:data<=-16'd13799;
      86629:data<=-16'd13782;
      86630:data<=-16'd15664;
      86631:data<=-16'd15179;
      86632:data<=-16'd13647;
      86633:data<=-16'd14064;
      86634:data<=-16'd13142;
      86635:data<=-16'd12962;
      86636:data<=-16'd14424;
      86637:data<=-16'd13374;
      86638:data<=-16'd12736;
      86639:data<=-16'd13230;
      86640:data<=-16'd12477;
      86641:data<=-16'd12760;
      86642:data<=-16'd13203;
      86643:data<=-16'd12995;
      86644:data<=-16'd12945;
      86645:data<=-16'd12921;
      86646:data<=-16'd14324;
      86647:data<=-16'd13746;
      86648:data<=-16'd12736;
      86649:data<=-16'd15920;
      86650:data<=-16'd11796;
      86651:data<=-16'd663;
      86652:data<=16'd1383;
      86653:data<=-16'd241;
      86654:data<=16'd758;
      86655:data<=-16'd1494;
      86656:data<=-16'd2196;
      86657:data<=-16'd368;
      86658:data<=-16'd946;
      86659:data<=-16'd1045;
      86660:data<=-16'd1442;
      86661:data<=-16'd2955;
      86662:data<=-16'd2557;
      86663:data<=-16'd2177;
      86664:data<=-16'd2232;
      86665:data<=-16'd1623;
      86666:data<=-16'd1983;
      86667:data<=-16'd2846;
      86668:data<=-16'd3149;
      86669:data<=-16'd3048;
      86670:data<=-16'd3116;
      86671:data<=-16'd3353;
      86672:data<=-16'd3046;
      86673:data<=-16'd3523;
      86674:data<=-16'd4411;
      86675:data<=-16'd4108;
      86676:data<=-16'd4040;
      86677:data<=-16'd4065;
      86678:data<=-16'd3968;
      86679:data<=-16'd4156;
      86680:data<=-16'd3162;
      86681:data<=-16'd2584;
      86682:data<=-16'd2652;
      86683:data<=-16'd1835;
      86684:data<=-16'd2061;
      86685:data<=-16'd1415;
      86686:data<=16'd467;
      86687:data<=16'd397;
      86688:data<=16'd1071;
      86689:data<=16'd1348;
      86690:data<=16'd629;
      86691:data<=16'd3037;
      86692:data<=16'd567;
      86693:data<=-16'd8056;
      86694:data<=-16'd9767;
      86695:data<=-16'd6940;
      86696:data<=-16'd6476;
      86697:data<=-16'd5529;
      86698:data<=-16'd4223;
      86699:data<=-16'd2429;
      86700:data<=-16'd1125;
      86701:data<=-16'd2196;
      86702:data<=-16'd1686;
      86703:data<=-16'd602;
      86704:data<=-16'd525;
      86705:data<=16'd1864;
      86706:data<=16'd2719;
      86707:data<=16'd930;
      86708:data<=16'd1422;
      86709:data<=16'd2155;
      86710:data<=16'd2140;
      86711:data<=16'd3372;
      86712:data<=16'd4112;
      86713:data<=16'd4305;
      86714:data<=16'd4579;
      86715:data<=16'd4132;
      86716:data<=16'd4034;
      86717:data<=16'd5344;
      86718:data<=16'd6813;
      86719:data<=16'd6630;
      86720:data<=16'd6203;
      86721:data<=16'd6670;
      86722:data<=16'd6120;
      86723:data<=16'd6411;
      86724:data<=16'd8288;
      86725:data<=16'd8254;
      86726:data<=16'd7767;
      86727:data<=16'd7882;
      86728:data<=16'd7451;
      86729:data<=16'd8319;
      86730:data<=16'd9216;
      86731:data<=16'd9520;
      86732:data<=16'd9561;
      86733:data<=16'd7712;
      86734:data<=16'd10877;
      86735:data<=16'd20083;
      86736:data<=16'd23325;
      86737:data<=16'd21963;
      86738:data<=16'd22503;
      86739:data<=16'd21655;
      86740:data<=16'd20325;
      86741:data<=16'd19685;
      86742:data<=16'd18911;
      86743:data<=16'd20125;
      86744:data<=16'd20002;
      86745:data<=16'd17294;
      86746:data<=16'd15916;
      86747:data<=16'd14856;
      86748:data<=16'd14707;
      86749:data<=16'd16161;
      86750:data<=16'd15887;
      86751:data<=16'd15065;
      86752:data<=16'd14794;
      86753:data<=16'd13982;
      86754:data<=16'd14093;
      86755:data<=16'd14352;
      86756:data<=16'd13808;
      86757:data<=16'd13584;
      86758:data<=16'd13045;
      86759:data<=16'd12111;
      86760:data<=16'd11840;
      86761:data<=16'd12631;
      86762:data<=16'd13044;
      86763:data<=16'd11650;
      86764:data<=16'd10977;
      86765:data<=16'd11380;
      86766:data<=16'd10668;
      86767:data<=16'd10740;
      86768:data<=16'd11414;
      86769:data<=16'd10851;
      86770:data<=16'd10634;
      86771:data<=16'd10657;
      86772:data<=16'd10204;
      86773:data<=16'd9661;
      86774:data<=16'd10135;
      86775:data<=16'd11634;
      86776:data<=16'd7491;
      86777:data<=-16'd1735;
      86778:data<=-16'd4921;
      86779:data<=-16'd3732;
      86780:data<=-16'd4611;
      86781:data<=-16'd4454;
      86782:data<=-16'd3795;
      86783:data<=-16'd4269;
      86784:data<=-16'd3946;
      86785:data<=-16'd4288;
      86786:data<=-16'd5303;
      86787:data<=-16'd5665;
      86788:data<=-16'd6162;
      86789:data<=-16'd6216;
      86790:data<=-16'd5702;
      86791:data<=-16'd5523;
      86792:data<=-16'd6423;
      86793:data<=-16'd8031;
      86794:data<=-16'd8090;
      86795:data<=-16'd6968;
      86796:data<=-16'd5761;
      86797:data<=-16'd4564;
      86798:data<=-16'd5557;
      86799:data<=-16'd7210;
      86800:data<=-16'd6805;
      86801:data<=-16'd6529;
      86802:data<=-16'd6557;
      86803:data<=-16'd6152;
      86804:data<=-16'd6561;
      86805:data<=-16'd7274;
      86806:data<=-16'd7811;
      86807:data<=-16'd7762;
      86808:data<=-16'd7424;
      86809:data<=-16'd7460;
      86810:data<=-16'd6843;
      86811:data<=-16'd7686;
      86812:data<=-16'd9818;
      86813:data<=-16'd9241;
      86814:data<=-16'd8608;
      86815:data<=-16'd8496;
      86816:data<=-16'd7504;
      86817:data<=-16'd9330;
      86818:data<=-16'd7488;
      86819:data<=16'd1709;
      86820:data<=16'd5530;
      86821:data<=16'd3706;
      86822:data<=16'd4364;
      86823:data<=16'd3617;
      86824:data<=16'd1459;
      86825:data<=16'd1515;
      86826:data<=16'd1136;
      86827:data<=16'd491;
      86828:data<=16'd696;
      86829:data<=-16'd121;
      86830:data<=-16'd1606;
      86831:data<=-16'd2347;
      86832:data<=-16'd2384;
      86833:data<=-16'd2293;
      86834:data<=-16'd1621;
      86835:data<=-16'd734;
      86836:data<=-16'd2052;
      86837:data<=-16'd4064;
      86838:data<=-16'd3900;
      86839:data<=-16'd3805;
      86840:data<=-16'd4237;
      86841:data<=-16'd3413;
      86842:data<=-16'd3806;
      86843:data<=-16'd5800;
      86844:data<=-16'd6043;
      86845:data<=-16'd5914;
      86846:data<=-16'd7432;
      86847:data<=-16'd7835;
      86848:data<=-16'd7503;
      86849:data<=-16'd8849;
      86850:data<=-16'd9100;
      86851:data<=-16'd7982;
      86852:data<=-16'd8305;
      86853:data<=-16'd7973;
      86854:data<=-16'd7204;
      86855:data<=-16'd8282;
      86856:data<=-16'd8493;
      86857:data<=-16'd8269;
      86858:data<=-16'd8466;
      86859:data<=-16'd6607;
      86860:data<=-16'd8856;
      86861:data<=-16'd18163;
      86862:data<=-16'd23134;
      86863:data<=-16'd21208;
      86864:data<=-16'd20447;
      86865:data<=-16'd20316;
      86866:data<=-16'd18628;
      86867:data<=-16'd18356;
      86868:data<=-16'd19108;
      86869:data<=-16'd18671;
      86870:data<=-16'd17794;
      86871:data<=-16'd17097;
      86872:data<=-16'd16073;
      86873:data<=-16'd15653;
      86874:data<=-16'd16587;
      86875:data<=-16'd17001;
      86876:data<=-16'd16001;
      86877:data<=-16'd15024;
      86878:data<=-16'd14358;
      86879:data<=-16'd13761;
      86880:data<=-16'd13204;
      86881:data<=-16'd12311;
      86882:data<=-16'd11486;
      86883:data<=-16'd10675;
      86884:data<=-16'd10113;
      86885:data<=-16'd10314;
      86886:data<=-16'd9132;
      86887:data<=-16'd6784;
      86888:data<=-16'd6155;
      86889:data<=-16'd5726;
      86890:data<=-16'd4619;
      86891:data<=-16'd4349;
      86892:data<=-16'd3263;
      86893:data<=-16'd1522;
      86894:data<=-16'd1221;
      86895:data<=-16'd817;
      86896:data<=16'd579;
      86897:data<=16'd1236;
      86898:data<=16'd1466;
      86899:data<=16'd3371;
      86900:data<=16'd4714;
      86901:data<=16'd3005;
      86902:data<=16'd5280;
      86903:data<=16'd13714;
      86904:data<=16'd17822;
      86905:data<=16'd17327;
      86906:data<=16'd18539;
      86907:data<=16'd18319;
      86908:data<=16'd17091;
      86909:data<=16'd17176;
      86910:data<=16'd15676;
      86911:data<=16'd15411;
      86912:data<=16'd17337;
      86913:data<=16'd16650;
      86914:data<=16'd15383;
      86915:data<=16'd15544;
      86916:data<=16'd14897;
      86917:data<=16'd14913;
      86918:data<=16'd16149;
      86919:data<=16'd16084;
      86920:data<=16'd14932;
      86921:data<=16'd14375;
      86922:data<=16'd14076;
      86923:data<=16'd13708;
      86924:data<=16'd14408;
      86925:data<=16'd14939;
      86926:data<=16'd13849;
      86927:data<=16'd13383;
      86928:data<=16'd13394;
      86929:data<=16'd12513;
      86930:data<=16'd12824;
      86931:data<=16'd13638;
      86932:data<=16'd13157;
      86933:data<=16'd13097;
      86934:data<=16'd13171;
      86935:data<=16'd12225;
      86936:data<=16'd12236;
      86937:data<=16'd13436;
      86938:data<=16'd13229;
      86939:data<=16'd12281;
      86940:data<=16'd12396;
      86941:data<=16'd11197;
      86942:data<=16'd10170;
      86943:data<=16'd12800;
      86944:data<=16'd11247;
      86945:data<=16'd1859;
      86946:data<=-16'd4334;
      86947:data<=-16'd4582;
      86948:data<=-16'd4505;
      86949:data<=-16'd3359;
      86950:data<=-16'd1835;
      86951:data<=-16'd2123;
      86952:data<=-16'd1979;
      86953:data<=-16'd1410;
      86954:data<=-16'd1858;
      86955:data<=-16'd1533;
      86956:data<=-16'd190;
      86957:data<=16'd0;
      86958:data<=-16'd179;
      86959:data<=16'd505;
      86960:data<=16'd176;
      86961:data<=-16'd205;
      86962:data<=16'd1149;
      86963:data<=16'd1513;
      86964:data<=16'd1118;
      86965:data<=16'd1597;
      86966:data<=16'd1149;
      86967:data<=16'd1330;
      86968:data<=16'd2849;
      86969:data<=16'd2905;
      86970:data<=16'd2704;
      86971:data<=16'd2796;
      86972:data<=16'd2302;
      86973:data<=16'd2992;
      86974:data<=16'd3809;
      86975:data<=16'd3653;
      86976:data<=16'd4012;
      86977:data<=16'd3952;
      86978:data<=16'd3215;
      86979:data<=16'd2928;
      86980:data<=16'd2663;
      86981:data<=16'd2337;
      86982:data<=16'd2012;
      86983:data<=16'd2046;
      86984:data<=16'd1944;
      86985:data<=16'd290;
      86986:data<=16'd984;
      86987:data<=16'd7241;
      86988:data<=16'd12407;
      86989:data<=16'd11884;
      86990:data<=16'd10416;
      86991:data<=16'd10514;
      86992:data<=16'd9743;
      86993:data<=16'd7815;
      86994:data<=16'd6296;
      86995:data<=16'd6105;
      86996:data<=16'd7048;
      86997:data<=16'd7515;
      86998:data<=16'd6863;
      86999:data<=16'd5363;
      87000:data<=16'd3334;
      87001:data<=16'd2766;
      87002:data<=16'd3334;
      87003:data<=16'd2952;
      87004:data<=16'd2813;
      87005:data<=16'd1986;
      87006:data<=-16'd370;
      87007:data<=-16'd549;
      87008:data<=-16'd58;
      87009:data<=-16'd1111;
      87010:data<=-16'd635;
      87011:data<=-16'd907;
      87012:data<=-16'd3234;
      87013:data<=-16'd3284;
      87014:data<=-16'd2983;
      87015:data<=-16'd4115;
      87016:data<=-16'd3668;
      87017:data<=-16'd3298;
      87018:data<=-16'd4673;
      87019:data<=-16'd5450;
      87020:data<=-16'd5184;
      87021:data<=-16'd4971;
      87022:data<=-16'd5049;
      87023:data<=-16'd5081;
      87024:data<=-16'd5504;
      87025:data<=-16'd7031;
      87026:data<=-16'd7671;
      87027:data<=-16'd6202;
      87028:data<=-16'd6902;
      87029:data<=-16'd13279;
      87030:data<=-16'd20463;
      87031:data<=-16'd22178;
      87032:data<=-16'd20877;
      87033:data<=-16'd20744;
      87034:data<=-16'd20143;
      87035:data<=-16'd18628;
      87036:data<=-16'd18393;
      87037:data<=-16'd19138;
      87038:data<=-16'd19250;
      87039:data<=-16'd18369;
      87040:data<=-16'd17752;
      87041:data<=-16'd17528;
      87042:data<=-16'd16719;
      87043:data<=-16'd16819;
      87044:data<=-16'd17644;
      87045:data<=-16'd17261;
      87046:data<=-16'd17468;
      87047:data<=-16'd18087;
      87048:data<=-16'd16957;
      87049:data<=-16'd16551;
      87050:data<=-16'd17332;
      87051:data<=-16'd16710;
      87052:data<=-16'd16095;
      87053:data<=-16'd16093;
      87054:data<=-16'd14973;
      87055:data<=-16'd14483;
      87056:data<=-16'd15244;
      87057:data<=-16'd14606;
      87058:data<=-16'd13661;
      87059:data<=-16'd13890;
      87060:data<=-16'd13097;
      87061:data<=-16'd12366;
      87062:data<=-16'd13488;
      87063:data<=-16'd13687;
      87064:data<=-16'd12592;
      87065:data<=-16'd12125;
      87066:data<=-16'd11765;
      87067:data<=-16'd11242;
      87068:data<=-16'd11044;
      87069:data<=-16'd11949;
      87070:data<=-16'd11749;
      87071:data<=-16'd5368;
      87072:data<=16'd2728;
      87073:data<=16'd4150;
      87074:data<=16'd2264;
      87075:data<=16'd1839;
      87076:data<=16'd1512;
      87077:data<=16'd1275;
      87078:data<=16'd1289;
      87079:data<=16'd1413;
      87080:data<=16'd2074;
      87081:data<=16'd2130;
      87082:data<=16'd1968;
      87083:data<=16'd2493;
      87084:data<=16'd2760;
      87085:data<=16'd2790;
      87086:data<=16'd3137;
      87087:data<=16'd4091;
      87088:data<=16'd4936;
      87089:data<=16'd4673;
      87090:data<=16'd4974;
      87091:data<=16'd5629;
      87092:data<=16'd5025;
      87093:data<=16'd5636;
      87094:data<=16'd7021;
      87095:data<=16'd6551;
      87096:data<=16'd7062;
      87097:data<=16'd8812;
      87098:data<=16'd8526;
      87099:data<=16'd8246;
      87100:data<=16'd9679;
      87101:data<=16'd10279;
      87102:data<=16'd9981;
      87103:data<=16'd9959;
      87104:data<=16'd9379;
      87105:data<=16'd9401;
      87106:data<=16'd10985;
      87107:data<=16'd11230;
      87108:data<=16'd10580;
      87109:data<=16'd11056;
      87110:data<=16'd9966;
      87111:data<=16'd9479;
      87112:data<=16'd11585;
      87113:data<=16'd7409;
      87114:data<=-16'd1782;
      87115:data<=-16'd3671;
      87116:data<=-16'd1415;
      87117:data<=-16'd2091;
      87118:data<=-16'd1425;
      87119:data<=16'd717;
      87120:data<=16'd719;
      87121:data<=16'd552;
      87122:data<=16'd995;
      87123:data<=16'd704;
      87124:data<=16'd1071;
      87125:data<=16'd2728;
      87126:data<=16'd3381;
      87127:data<=16'd2899;
      87128:data<=16'd3133;
      87129:data<=16'd3028;
      87130:data<=16'd2830;
      87131:data<=16'd4546;
      87132:data<=16'd5562;
      87133:data<=16'd4766;
      87134:data<=16'd4828;
      87135:data<=16'd4931;
      87136:data<=16'd4755;
      87137:data<=16'd5806;
      87138:data<=16'd6667;
      87139:data<=16'd6595;
      87140:data<=16'd6683;
      87141:data<=16'd6974;
      87142:data<=16'd6498;
      87143:data<=16'd6015;
      87144:data<=16'd7550;
      87145:data<=16'd8320;
      87146:data<=16'd6485;
      87147:data<=16'd5635;
      87148:data<=16'd4855;
      87149:data<=16'd4373;
      87150:data<=16'd6748;
      87151:data<=16'd6975;
      87152:data<=16'd5836;
      87153:data<=16'd6536;
      87154:data<=16'd5074;
      87155:data<=16'd8945;
      87156:data<=16'd20084;
      87157:data<=16'd22316;
      87158:data<=16'd18319;
      87159:data<=16'd19202;
      87160:data<=16'd18936;
      87161:data<=16'd16791;
      87162:data<=16'd17256;
      87163:data<=16'd17575;
      87164:data<=16'd17214;
      87165:data<=16'd16980;
      87166:data<=16'd16069;
      87167:data<=16'd14625;
      87168:data<=16'd14339;
      87169:data<=16'd16146;
      87170:data<=16'd16136;
      87171:data<=16'd14437;
      87172:data<=16'd14512;
      87173:data<=16'd13415;
      87174:data<=16'd12760;
      87175:data<=16'd14795;
      87176:data<=16'd14055;
      87177:data<=16'd12322;
      87178:data<=16'd12536;
      87179:data<=16'd11627;
      87180:data<=16'd11188;
      87181:data<=16'd11260;
      87182:data<=16'd10029;
      87183:data<=16'd9285;
      87184:data<=16'd8678;
      87185:data<=16'd8194;
      87186:data<=16'd7542;
      87187:data<=16'd5912;
      87188:data<=16'd5398;
      87189:data<=16'd4936;
      87190:data<=16'd4097;
      87191:data<=16'd4184;
      87192:data<=16'd3427;
      87193:data<=16'd2984;
      87194:data<=16'd1691;
      87195:data<=-16'd461;
      87196:data<=16'd1595;
      87197:data<=-16'd452;
      87198:data<=-16'd9768;
      87199:data<=-16'd12713;
      87200:data<=-16'd11932;
      87201:data<=-16'd13932;
      87202:data<=-16'd12904;
      87203:data<=-16'd11590;
      87204:data<=-16'd12041;
      87205:data<=-16'd11556;
      87206:data<=-16'd12713;
      87207:data<=-16'd13344;
      87208:data<=-16'd12249;
      87209:data<=-16'd12480;
      87210:data<=-16'd12428;
      87211:data<=-16'd12157;
      87212:data<=-16'd12378;
      87213:data<=-16'd12357;
      87214:data<=-16'd12935;
      87215:data<=-16'd12780;
      87216:data<=-16'd11990;
      87217:data<=-16'd11544;
      87218:data<=-16'd11279;
      87219:data<=-16'd12601;
      87220:data<=-16'd12953;
      87221:data<=-16'd11627;
      87222:data<=-16'd11637;
      87223:data<=-16'd10760;
      87224:data<=-16'd10339;
      87225:data<=-16'd11963;
      87226:data<=-16'd11670;
      87227:data<=-16'd11362;
      87228:data<=-16'd11395;
      87229:data<=-16'd10055;
      87230:data<=-16'd10687;
      87231:data<=-16'd11667;
      87232:data<=-16'd11926;
      87233:data<=-16'd12366;
      87234:data<=-16'd11150;
      87235:data<=-16'd11207;
      87236:data<=-16'd10593;
      87237:data<=-16'd8986;
      87238:data<=-16'd12437;
      87239:data<=-16'd9644;
      87240:data<=16'd1792;
      87241:data<=16'd4267;
      87242:data<=16'd2190;
      87243:data<=16'd2939;
      87244:data<=16'd440;
      87245:data<=-16'd197;
      87246:data<=16'd887;
      87247:data<=-16'd1472;
      87248:data<=-16'd1865;
      87249:data<=-16'd1780;
      87250:data<=-16'd3674;
      87251:data<=-16'd3632;
      87252:data<=-16'd3063;
      87253:data<=-16'd3034;
      87254:data<=-16'd3093;
      87255:data<=-16'd3247;
      87256:data<=-16'd3184;
      87257:data<=-16'd4676;
      87258:data<=-16'd5241;
      87259:data<=-16'd4165;
      87260:data<=-16'd4802;
      87261:data<=-16'd4252;
      87262:data<=-16'd3909;
      87263:data<=-16'd6390;
      87264:data<=-16'd6076;
      87265:data<=-16'd4493;
      87266:data<=-16'd4952;
      87267:data<=-16'd4834;
      87268:data<=-16'd5513;
      87269:data<=-16'd6576;
      87270:data<=-16'd6270;
      87271:data<=-16'd6135;
      87272:data<=-16'd5891;
      87273:data<=-16'd5997;
      87274:data<=-16'd6079;
      87275:data<=-16'd6020;
      87276:data<=-16'd7183;
      87277:data<=-16'd6693;
      87278:data<=-16'd6288;
      87279:data<=-16'd7009;
      87280:data<=-16'd4270;
      87281:data<=-16'd6692;
      87282:data<=-16'd16645;
      87283:data<=-16'd19294;
      87284:data<=-16'd16443;
      87285:data<=-16'd16328;
      87286:data<=-16'd15317;
      87287:data<=-16'd13696;
      87288:data<=-16'd12515;
      87289:data<=-16'd10977;
      87290:data<=-16'd10370;
      87291:data<=-16'd9726;
      87292:data<=-16'd9564;
      87293:data<=-16'd8678;
      87294:data<=-16'd6034;
      87295:data<=-16'd5665;
      87296:data<=-16'd5042;
      87297:data<=-16'd2558;
      87298:data<=-16'd2643;
      87299:data<=-16'd2150;
      87300:data<=16'd71;
      87301:data<=16'd458;
      87302:data<=16'd826;
      87303:data<=16'd1392;
      87304:data<=16'd1372;
      87305:data<=16'd1594;
      87306:data<=16'd2076;
      87307:data<=16'd3486;
      87308:data<=16'd3823;
      87309:data<=16'd3607;
      87310:data<=16'd4767;
      87311:data<=16'd3982;
      87312:data<=16'd4096;
      87313:data<=16'd6830;
      87314:data<=16'd6457;
      87315:data<=16'd5823;
      87316:data<=16'd6252;
      87317:data<=16'd5171;
      87318:data<=16'd6407;
      87319:data<=16'd7680;
      87320:data<=16'd7638;
      87321:data<=16'd8396;
      87322:data<=16'd6378;
      87323:data<=16'd8893;
      87324:data<=16'd18766;
      87325:data<=16'd22192;
      87326:data<=16'd20889;
      87327:data<=16'd21546;
      87328:data<=16'd20168;
      87329:data<=16'd19017;
      87330:data<=16'd18607;
      87331:data<=16'd17843;
      87332:data<=16'd19465;
      87333:data<=16'd19494;
      87334:data<=16'd17975;
      87335:data<=16'd18114;
      87336:data<=16'd17100;
      87337:data<=16'd17088;
      87338:data<=16'd18352;
      87339:data<=16'd17197;
      87340:data<=16'd16318;
      87341:data<=16'd16048;
      87342:data<=16'd15268;
      87343:data<=16'd15412;
      87344:data<=16'd15353;
      87345:data<=16'd15170;
      87346:data<=16'd14283;
      87347:data<=16'd12337;
      87348:data<=16'd11696;
      87349:data<=16'd11080;
      87350:data<=16'd11171;
      87351:data<=16'd12627;
      87352:data<=16'd11579;
      87353:data<=16'd10704;
      87354:data<=16'd11195;
      87355:data<=16'd9626;
      87356:data<=16'd9498;
      87357:data<=16'd10904;
      87358:data<=16'd10589;
      87359:data<=16'd10132;
      87360:data<=16'd9360;
      87361:data<=16'd8940;
      87362:data<=16'd9118;
      87363:data<=16'd9151;
      87364:data<=16'd10545;
      87365:data<=16'd7068;
      87366:data<=-16'd2141;
      87367:data<=-16'd5451;
      87368:data<=-16'd4152;
      87369:data<=-16'd4015;
      87370:data<=-16'd2541;
      87371:data<=-16'd2040;
      87372:data<=-16'd2638;
      87373:data<=-16'd2046;
      87374:data<=-16'd2538;
      87375:data<=-16'd2153;
      87376:data<=-16'd503;
      87377:data<=-16'd472;
      87378:data<=-16'd731;
      87379:data<=-16'd1216;
      87380:data<=-16'd1459;
      87381:data<=-16'd799;
      87382:data<=-16'd1227;
      87383:data<=-16'd1466;
      87384:data<=-16'd1465;
      87385:data<=-16'd2050;
      87386:data<=-16'd1331;
      87387:data<=-16'd1744;
      87388:data<=-16'd3756;
      87389:data<=-16'd4065;
      87390:data<=-16'd4074;
      87391:data<=-16'd4329;
      87392:data<=-16'd4235;
      87393:data<=-16'd4555;
      87394:data<=-16'd4955;
      87395:data<=-16'd6123;
      87396:data<=-16'd6275;
      87397:data<=-16'd4593;
      87398:data<=-16'd4117;
      87399:data<=-16'd3633;
      87400:data<=-16'd4065;
      87401:data<=-16'd6469;
      87402:data<=-16'd6213;
      87403:data<=-16'd5714;
      87404:data<=-16'd5941;
      87405:data<=-16'd4602;
      87406:data<=-16'd6862;
      87407:data<=-16'd5967;
      87408:data<=16'd3545;
      87409:data<=16'd6983;
      87410:data<=16'd4669;
      87411:data<=16'd5858;
      87412:data<=16'd4451;
      87413:data<=16'd1688;
      87414:data<=16'd2068;
      87415:data<=16'd1445;
      87416:data<=16'd694;
      87417:data<=16'd889;
      87418:data<=16'd638;
      87419:data<=-16'd227;
      87420:data<=-16'd2406;
      87421:data<=-16'd2726;
      87422:data<=-16'd1718;
      87423:data<=-16'd2622;
      87424:data<=-16'd2268;
      87425:data<=-16'd2628;
      87426:data<=-16'd5347;
      87427:data<=-16'd5077;
      87428:data<=-16'd4501;
      87429:data<=-16'd5677;
      87430:data<=-16'd5012;
      87431:data<=-16'd5397;
      87432:data<=-16'd7219;
      87433:data<=-16'd7007;
      87434:data<=-16'd6537;
      87435:data<=-16'd6901;
      87436:data<=-16'd6957;
      87437:data<=-16'd6966;
      87438:data<=-16'd7755;
      87439:data<=-16'd8493;
      87440:data<=-16'd8064;
      87441:data<=-16'd8381;
      87442:data<=-16'd8513;
      87443:data<=-16'd7257;
      87444:data<=-16'd8510;
      87445:data<=-16'd9993;
      87446:data<=-16'd9406;
      87447:data<=-16'd10458;
      87448:data<=-16'd10530;
      87449:data<=-16'd12322;
      87450:data<=-16'd21156;
      87451:data<=-16'd26292;
      87452:data<=-16'd24139;
      87453:data<=-16'd23566;
      87454:data<=-16'd23175;
      87455:data<=-16'd21218;
      87456:data<=-16'd21168;
      87457:data<=-16'd22037;
      87458:data<=-16'd21754;
      87459:data<=-16'd20271;
      87460:data<=-16'd19635;
      87461:data<=-16'd19473;
      87462:data<=-16'd18049;
      87463:data<=-16'd18730;
      87464:data<=-16'd19901;
      87465:data<=-16'd17758;
      87466:data<=-16'd16883;
      87467:data<=-16'd17064;
      87468:data<=-16'd15509;
      87469:data<=-16'd15805;
      87470:data<=-16'd16633;
      87471:data<=-16'd15440;
      87472:data<=-16'd14871;
      87473:data<=-16'd14895;
      87474:data<=-16'd14107;
      87475:data<=-16'd13561;
      87476:data<=-16'd14169;
      87477:data<=-16'd14081;
      87478:data<=-16'd12408;
      87479:data<=-16'd12135;
      87480:data<=-16'd12336;
      87481:data<=-16'd10971;
      87482:data<=-16'd10396;
      87483:data<=-16'd9744;
      87484:data<=-16'd8784;
      87485:data<=-16'd8937;
      87486:data<=-16'd8006;
      87487:data<=-16'd7157;
      87488:data<=-16'd6076;
      87489:data<=-16'd3921;
      87490:data<=-16'd4943;
      87491:data<=-16'd2258;
      87492:data<=16'd7536;
      87493:data<=16'd10981;
      87494:data<=16'd9824;
      87495:data<=16'd12275;
      87496:data<=16'd12357;
      87497:data<=16'd11659;
      87498:data<=16'd13458;
      87499:data<=16'd13197;
      87500:data<=16'd13279;
      87501:data<=16'd14675;
      87502:data<=16'd14430;
      87503:data<=16'd14199;
      87504:data<=16'd13502;
      87505:data<=16'd12602;
      87506:data<=16'd13670;
      87507:data<=16'd14440;
      87508:data<=16'd14169;
      87509:data<=16'd14157;
      87510:data<=16'd13819;
      87511:data<=16'd13221;
      87512:data<=16'd13012;
      87513:data<=16'd13740;
      87514:data<=16'd14468;
      87515:data<=16'd13785;
      87516:data<=16'd13151;
      87517:data<=16'd12969;
      87518:data<=16'd12302;
      87519:data<=16'd12430;
      87520:data<=16'd13397;
      87521:data<=16'd13732;
      87522:data<=16'd13562;
      87523:data<=16'd13241;
      87524:data<=16'd12480;
      87525:data<=16'd12196;
      87526:data<=16'd13379;
      87527:data<=16'd13776;
      87528:data<=16'd12657;
      87529:data<=16'd12634;
      87530:data<=16'd12242;
      87531:data<=16'd11837;
      87532:data<=16'd14310;
      87533:data<=16'd12289;
      87534:data<=16'd3078;
      87535:data<=-16'd1550;
      87536:data<=-16'd159;
      87537:data<=-16'd299;
      87538:data<=-16'd2;
      87539:data<=16'd2058;
      87540:data<=16'd2030;
      87541:data<=16'd1072;
      87542:data<=16'd1519;
      87543:data<=16'd1967;
      87544:data<=16'd2288;
      87545:data<=16'd3704;
      87546:data<=16'd4411;
      87547:data<=16'd2928;
      87548:data<=16'd1478;
      87549:data<=16'd1334;
      87550:data<=16'd1912;
      87551:data<=16'd2951;
      87552:data<=16'd3459;
      87553:data<=16'd3489;
      87554:data<=16'd3711;
      87555:data<=16'd3315;
      87556:data<=16'd3052;
      87557:data<=16'd3974;
      87558:data<=16'd4757;
      87559:data<=16'd4728;
      87560:data<=16'd4337;
      87561:data<=16'd3955;
      87562:data<=16'd3997;
      87563:data<=16'd4629;
      87564:data<=16'd5667;
      87565:data<=16'd5956;
      87566:data<=16'd5565;
      87567:data<=16'd5582;
      87568:data<=16'd5033;
      87569:data<=16'd5283;
      87570:data<=16'd7330;
      87571:data<=16'd7109;
      87572:data<=16'd6216;
      87573:data<=16'd6969;
      87574:data<=16'd5062;
      87575:data<=16'd6484;
      87576:data<=16'd16181;
      87577:data<=16'd21153;
      87578:data<=16'd18618;
      87579:data<=16'd18395;
      87580:data<=16'd18377;
      87581:data<=16'd16452;
      87582:data<=16'd16321;
      87583:data<=16'd16128;
      87584:data<=16'd15120;
      87585:data<=16'd14428;
      87586:data<=16'd13377;
      87587:data<=16'd12810;
      87588:data<=16'd11620;
      87589:data<=16'd9347;
      87590:data<=16'd8708;
      87591:data<=16'd8696;
      87592:data<=16'd8076;
      87593:data<=16'd7964;
      87594:data<=16'd6766;
      87595:data<=16'd4323;
      87596:data<=16'd3662;
      87597:data<=16'd4751;
      87598:data<=16'd5269;
      87599:data<=16'd5071;
      87600:data<=16'd4407;
      87601:data<=16'd2740;
      87602:data<=16'd1706;
      87603:data<=16'd1739;
      87604:data<=16'd957;
      87605:data<=16'd948;
      87606:data<=16'd1465;
      87607:data<=-16'd614;
      87608:data<=-16'd2541;
      87609:data<=-16'd2303;
      87610:data<=-16'd2209;
      87611:data<=-16'd2184;
      87612:data<=-16'd2438;
      87613:data<=-16'd3465;
      87614:data<=-16'd4604;
      87615:data<=-16'd5068;
      87616:data<=-16'd3691;
      87617:data<=-16'd5382;
      87618:data<=-16'd13221;
      87619:data<=-16'd18651;
      87620:data<=-16'd18816;
      87621:data<=-16'd18766;
      87622:data<=-16'd18565;
      87623:data<=-16'd18134;
      87624:data<=-16'd17699;
      87625:data<=-16'd17221;
      87626:data<=-16'd18421;
      87627:data<=-16'd18944;
      87628:data<=-16'd17813;
      87629:data<=-16'd17456;
      87630:data<=-16'd16565;
      87631:data<=-16'd15756;
      87632:data<=-16'd16917;
      87633:data<=-16'd17640;
      87634:data<=-16'd16897;
      87635:data<=-16'd16198;
      87636:data<=-16'd15764;
      87637:data<=-16'd14663;
      87638:data<=-16'd14484;
      87639:data<=-16'd16334;
      87640:data<=-16'd15957;
      87641:data<=-16'd14248;
      87642:data<=-16'd14713;
      87643:data<=-16'd13467;
      87644:data<=-16'd12693;
      87645:data<=-16'd14916;
      87646:data<=-16'd13932;
      87647:data<=-16'd13007;
      87648:data<=-16'd15221;
      87649:data<=-16'd14490;
      87650:data<=-16'd13402;
      87651:data<=-16'd14666;
      87652:data<=-16'd14737;
      87653:data<=-16'd13964;
      87654:data<=-16'd13047;
      87655:data<=-16'd12797;
      87656:data<=-16'd12665;
      87657:data<=-16'd12138;
      87658:data<=-16'd14331;
      87659:data<=-16'd13041;
      87660:data<=-16'd4058;
      87661:data<=16'd1535;
      87662:data<=16'd1478;
      87663:data<=16'd1231;
      87664:data<=-16'd47;
      87665:data<=-16'd435;
      87666:data<=16'd326;
      87667:data<=16'd191;
      87668:data<=16'd981;
      87669:data<=16'd860;
      87670:data<=-16'd826;
      87671:data<=-16'd1077;
      87672:data<=-16'd1096;
      87673:data<=-16'd1336;
      87674:data<=-16'd840;
      87675:data<=-16'd799;
      87676:data<=-16'd1498;
      87677:data<=-16'd2202;
      87678:data<=-16'd1985;
      87679:data<=-16'd1712;
      87680:data<=-16'd2202;
      87681:data<=-16'd1676;
      87682:data<=-16'd1137;
      87683:data<=-16'd1575;
      87684:data<=-16'd1183;
      87685:data<=-16'd823;
      87686:data<=-16'd892;
      87687:data<=-16'd792;
      87688:data<=-16'd476;
      87689:data<=16'd1460;
      87690:data<=16'd2681;
      87691:data<=16'd1777;
      87692:data<=16'd1944;
      87693:data<=16'd2073;
      87694:data<=16'd2194;
      87695:data<=16'd3940;
      87696:data<=16'd4029;
      87697:data<=16'd4323;
      87698:data<=16'd6707;
      87699:data<=16'd6680;
      87700:data<=16'd6798;
      87701:data<=16'd7692;
      87702:data<=16'd2385;
      87703:data<=-16'd4372;
      87704:data<=-16'd4739;
      87705:data<=-16'd3538;
      87706:data<=-16'd3996;
      87707:data<=-16'd2801;
      87708:data<=-16'd917;
      87709:data<=-16'd926;
      87710:data<=-16'd1051;
      87711:data<=-16'd353;
      87712:data<=-16'd370;
      87713:data<=16'd329;
      87714:data<=16'd2376;
      87715:data<=16'd2751;
      87716:data<=16'd2293;
      87717:data<=16'd3074;
      87718:data<=16'd3116;
      87719:data<=16'd2892;
      87720:data<=16'd4326;
      87721:data<=16'd5556;
      87722:data<=16'd5441;
      87723:data<=16'd5200;
      87724:data<=16'd5253;
      87725:data<=16'd5363;
      87726:data<=16'd6058;
      87727:data<=16'd7329;
      87728:data<=16'd7348;
      87729:data<=16'd6796;
      87730:data<=16'd7523;
      87731:data<=16'd7306;
      87732:data<=16'd6995;
      87733:data<=16'd8928;
      87734:data<=16'd9270;
      87735:data<=16'd8475;
      87736:data<=16'd9326;
      87737:data<=16'd8831;
      87738:data<=16'd8762;
      87739:data<=16'd10210;
      87740:data<=16'd9555;
      87741:data<=16'd9661;
      87742:data<=16'd9706;
      87743:data<=16'd8395;
      87744:data<=16'd14201;
      87745:data<=16'd22786;
      87746:data<=16'd23384;
      87747:data<=16'd21323;
      87748:data<=16'd20615;
      87749:data<=16'd18882;
      87750:data<=16'd17904;
      87751:data<=16'd18155;
      87752:data<=16'd18688;
      87753:data<=16'd18386;
      87754:data<=16'd17277;
      87755:data<=16'd17141;
      87756:data<=16'd16108;
      87757:data<=16'd15332;
      87758:data<=16'd17009;
      87759:data<=16'd16683;
      87760:data<=16'd15379;
      87761:data<=16'd15634;
      87762:data<=16'd14219;
      87763:data<=16'd13523;
      87764:data<=16'd14794;
      87765:data<=16'd14633;
      87766:data<=16'd13937;
      87767:data<=16'd12862;
      87768:data<=16'd11638;
      87769:data<=16'd11743;
      87770:data<=16'd11946;
      87771:data<=16'd12137;
      87772:data<=16'd11703;
      87773:data<=16'd11107;
      87774:data<=16'd11706;
      87775:data<=16'd10452;
      87776:data<=16'd9450;
      87777:data<=16'd11207;
      87778:data<=16'd10933;
      87779:data<=16'd9978;
      87780:data<=16'd9952;
      87781:data<=16'd8898;
      87782:data<=16'd8933;
      87783:data<=16'd7865;
      87784:data<=16'd6672;
      87785:data<=16'd7724;
      87786:data<=16'd2015;
      87787:data<=-16'd6986;
      87788:data<=-16'd8211;
      87789:data<=-16'd8202;
      87790:data<=-16'd10026;
      87791:data<=-16'd9409;
      87792:data<=-16'd9069;
      87793:data<=-16'd9407;
      87794:data<=-16'd9549;
      87795:data<=-16'd10302;
      87796:data<=-16'd10971;
      87797:data<=-16'd11303;
      87798:data<=-16'd9852;
      87799:data<=-16'd8290;
      87800:data<=-16'd8836;
      87801:data<=-16'd8798;
      87802:data<=-16'd9203;
      87803:data<=-16'd10307;
      87804:data<=-16'd9709;
      87805:data<=-16'd9723;
      87806:data<=-16'd9545;
      87807:data<=-16'd8950;
      87808:data<=-16'd10566;
      87809:data<=-16'd10857;
      87810:data<=-16'd10035;
      87811:data<=-16'd10454;
      87812:data<=-16'd9635;
      87813:data<=-16'd9706;
      87814:data<=-16'd11063;
      87815:data<=-16'd11059;
      87816:data<=-16'd11083;
      87817:data<=-16'd10434;
      87818:data<=-16'd9934;
      87819:data<=-16'd10574;
      87820:data<=-16'd10337;
      87821:data<=-16'd11436;
      87822:data<=-16'd11975;
      87823:data<=-16'd10520;
      87824:data<=-16'd11515;
      87825:data<=-16'd10564;
      87826:data<=-16'd9451;
      87827:data<=-16'd13217;
      87828:data<=-16'd8959;
      87829:data<=16'd1119;
      87830:data<=16'd1815;
      87831:data<=16'd617;
      87832:data<=16'd1670;
      87833:data<=-16'd866;
      87834:data<=-16'd1900;
      87835:data<=-16'd1142;
      87836:data<=-16'd1788;
      87837:data<=-16'd1246;
      87838:data<=-16'd1254;
      87839:data<=-16'd2766;
      87840:data<=-16'd3565;
      87841:data<=-16'd3526;
      87842:data<=-16'd3215;
      87843:data<=-16'd3742;
      87844:data<=-16'd3741;
      87845:data<=-16'd3501;
      87846:data<=-16'd5253;
      87847:data<=-16'd5418;
      87848:data<=-16'd5072;
      87849:data<=-16'd7327;
      87850:data<=-16'd7221;
      87851:data<=-16'd6905;
      87852:data<=-16'd9641;
      87853:data<=-16'd9697;
      87854:data<=-16'd8601;
      87855:data<=-16'd9197;
      87856:data<=-16'd8605;
      87857:data<=-16'd8557;
      87858:data<=-16'd9777;
      87859:data<=-16'd10263;
      87860:data<=-16'd9799;
      87861:data<=-16'd8619;
      87862:data<=-16'd8331;
      87863:data<=-16'd8311;
      87864:data<=-16'd8731;
      87865:data<=-16'd10445;
      87866:data<=-16'd9599;
      87867:data<=-16'd9083;
      87868:data<=-16'd10091;
      87869:data<=-16'd7027;
      87870:data<=-16'd10290;
      87871:data<=-16'd21924;
      87872:data<=-16'd23975;
      87873:data<=-16'd20513;
      87874:data<=-16'd21419;
      87875:data<=-16'd20148;
      87876:data<=-16'd19334;
      87877:data<=-16'd21220;
      87878:data<=-16'd20210;
      87879:data<=-16'd18598;
      87880:data<=-16'd17870;
      87881:data<=-16'd17315;
      87882:data<=-16'd17070;
      87883:data<=-16'd15320;
      87884:data<=-16'd14462;
      87885:data<=-16'd14472;
      87886:data<=-16'd13048;
      87887:data<=-16'd13092;
      87888:data<=-16'd12865;
      87889:data<=-16'd10323;
      87890:data<=-16'd9009;
      87891:data<=-16'd8573;
      87892:data<=-16'd7747;
      87893:data<=-16'd6987;
      87894:data<=-16'd6122;
      87895:data<=-16'd5133;
      87896:data<=-16'd3566;
      87897:data<=-16'd2793;
      87898:data<=-16'd1801;
      87899:data<=16'd789;
      87900:data<=16'd836;
      87901:data<=16'd550;
      87902:data<=16'd2798;
      87903:data<=16'd2922;
      87904:data<=16'd2939;
      87905:data<=16'd3970;
      87906:data<=16'd3142;
      87907:data<=16'd3736;
      87908:data<=16'd4974;
      87909:data<=16'd5726;
      87910:data<=16'd6273;
      87911:data<=16'd4008;
      87912:data<=16'd7655;
      87913:data<=16'd17825;
      87914:data<=16'd19964;
      87915:data<=16'd18252;
      87916:data<=16'd19549;
      87917:data<=16'd18851;
      87918:data<=16'd18613;
      87919:data<=16'd18434;
      87920:data<=16'd17206;
      87921:data<=16'd18997;
      87922:data<=16'd19387;
      87923:data<=16'd18230;
      87924:data<=16'd18713;
      87925:data<=16'd16948;
      87926:data<=16'd16175;
      87927:data<=16'd18039;
      87928:data<=16'd17743;
      87929:data<=16'd17174;
      87930:data<=16'd16722;
      87931:data<=16'd15649;
      87932:data<=16'd15973;
      87933:data<=16'd16325;
      87934:data<=16'd16521;
      87935:data<=16'd16060;
      87936:data<=16'd14725;
      87937:data<=16'd14989;
      87938:data<=16'd14468;
      87939:data<=16'd13443;
      87940:data<=16'd14624;
      87941:data<=16'd14537;
      87942:data<=16'd13902;
      87943:data<=16'd14184;
      87944:data<=16'd13207;
      87945:data<=16'd13352;
      87946:data<=16'd14466;
      87947:data<=16'd14354;
      87948:data<=16'd13248;
      87949:data<=16'd10919;
      87950:data<=16'd10182;
      87951:data<=16'd10339;
      87952:data<=16'd10067;
      87953:data<=16'd12098;
      87954:data<=16'd8502;
      87955:data<=-16'd1553;
      87956:data<=-16'd4091;
      87957:data<=-16'd2074;
      87958:data<=-16'd2520;
      87959:data<=-16'd1350;
      87960:data<=-16'd1021;
      87961:data<=-16'd1732;
      87962:data<=-16'd943;
      87963:data<=-16'd1914;
      87964:data<=-16'd1821;
      87965:data<=16'd525;
      87966:data<=16'd896;
      87967:data<=16'd1002;
      87968:data<=16'd1051;
      87969:data<=16'd23;
      87970:data<=16'd720;
      87971:data<=16'd2466;
      87972:data<=16'd3028;
      87973:data<=16'd2520;
      87974:data<=16'd2035;
      87975:data<=16'd2287;
      87976:data<=16'd2682;
      87977:data<=16'd3526;
      87978:data<=16'd4167;
      87979:data<=16'd3768;
      87980:data<=16'd3882;
      87981:data<=16'd3779;
      87982:data<=16'd3181;
      87983:data<=16'd3159;
      87984:data<=16'd2564;
      87985:data<=16'd2376;
      87986:data<=16'd2082;
      87987:data<=16'd861;
      87988:data<=16'd1633;
      87989:data<=16'd1327;
      87990:data<=-16'd905;
      87991:data<=-16'd611;
      87992:data<=-16'd1133;
      87993:data<=-16'd1633;
      87994:data<=-16'd481;
      87995:data<=-16'd3089;
      87996:data<=-16'd1410;
      87997:data<=16'd7694;
      87998:data<=16'd10299;
      87999:data<=16'd8869;
      88000:data<=16'd10574;
      88001:data<=16'd9814;
      88002:data<=16'd7844;
      88003:data<=16'd7330;
      88004:data<=16'd6440;
      88005:data<=16'd6150;
      88006:data<=16'd5695;
      88007:data<=16'd5183;
      88008:data<=16'd4546;
      88009:data<=16'd2349;
      88010:data<=16'd1648;
      88011:data<=16'd1804;
      88012:data<=16'd857;
      88013:data<=16'd1334;
      88014:data<=16'd758;
      88015:data<=-16'd1368;
      88016:data<=-16'd1365;
      88017:data<=-16'd1604;
      88018:data<=-16'd2372;
      88019:data<=-16'd1826;
      88020:data<=-16'd2523;
      88021:data<=-16'd4297;
      88022:data<=-16'd5002;
      88023:data<=-16'd4817;
      88024:data<=-16'd4925;
      88025:data<=-16'd5307;
      88026:data<=-16'd4686;
      88027:data<=-16'd5071;
      88028:data<=-16'd6628;
      88029:data<=-16'd6269;
      88030:data<=-16'd6307;
      88031:data<=-16'd6875;
      88032:data<=-16'd5964;
      88033:data<=-16'd6804;
      88034:data<=-16'd8111;
      88035:data<=-16'd8417;
      88036:data<=-16'd9065;
      88037:data<=-16'd7336;
      88038:data<=-16'd9175;
      88039:data<=-16'd18566;
      88040:data<=-16'd23073;
      88041:data<=-16'd20927;
      88042:data<=-16'd20662;
      88043:data<=-16'd20286;
      88044:data<=-16'd18850;
      88045:data<=-16'd19208;
      88046:data<=-16'd19840;
      88047:data<=-16'd19516;
      88048:data<=-16'd19203;
      88049:data<=-16'd19817;
      88050:data<=-16'd19613;
      88051:data<=-16'd18151;
      88052:data<=-16'd18756;
      88053:data<=-16'd19735;
      88054:data<=-16'd18748;
      88055:data<=-16'd18262;
      88056:data<=-16'd17515;
      88057:data<=-16'd16214;
      88058:data<=-16'd16528;
      88059:data<=-16'd16985;
      88060:data<=-16'd16510;
      88061:data<=-16'd15731;
      88062:data<=-16'd14684;
      88063:data<=-16'd13684;
      88064:data<=-16'd13248;
      88065:data<=-16'd13963;
      88066:data<=-16'd14063;
      88067:data<=-16'd12924;
      88068:data<=-16'd12803;
      88069:data<=-16'd12310;
      88070:data<=-16'd11858;
      88071:data<=-16'd13112;
      88072:data<=-16'd12498;
      88073:data<=-16'd11429;
      88074:data<=-16'd11737;
      88075:data<=-16'd10228;
      88076:data<=-16'd9589;
      88077:data<=-16'd9864;
      88078:data<=-16'd9385;
      88079:data<=-16'd11053;
      88080:data<=-16'd7397;
      88081:data<=16'd2754;
      88082:data<=16'd5741;
      88083:data<=16'd4128;
      88084:data<=16'd5438;
      88085:data<=16'd5262;
      88086:data<=16'd5042;
      88087:data<=16'd6047;
      88088:data<=16'd5230;
      88089:data<=16'd5800;
      88090:data<=16'd7802;
      88091:data<=16'd7674;
      88092:data<=16'd6837;
      88093:data<=16'd6816;
      88094:data<=16'd7001;
      88095:data<=16'd7319;
      88096:data<=16'd8479;
      88097:data<=16'd9300;
      88098:data<=16'd8898;
      88099:data<=16'd10193;
      88100:data<=16'd11740;
      88101:data<=16'd10689;
      88102:data<=16'd11100;
      88103:data<=16'd12515;
      88104:data<=16'd11688;
      88105:data<=16'd11673;
      88106:data<=16'd11981;
      88107:data<=16'd10608;
      88108:data<=16'd10611;
      88109:data<=16'd12267;
      88110:data<=16'd12839;
      88111:data<=16'd12111;
      88112:data<=16'd11838;
      88113:data<=16'd11761;
      88114:data<=16'd11264;
      88115:data<=16'd12609;
      88116:data<=16'd13333;
      88117:data<=16'd11327;
      88118:data<=16'd11697;
      88119:data<=16'd11908;
      88120:data<=16'd10155;
      88121:data<=16'd12605;
      88122:data<=16'd11226;
      88123:data<=16'd1530;
      88124:data<=-16'd2243;
      88125:data<=-16'd238;
      88126:data<=-16'd1328;
      88127:data<=-16'd1224;
      88128:data<=16'd884;
      88129:data<=16'd1149;
      88130:data<=16'd1118;
      88131:data<=16'd1202;
      88132:data<=16'd914;
      88133:data<=16'd1874;
      88134:data<=16'd3953;
      88135:data<=16'd4754;
      88136:data<=16'd4258;
      88137:data<=16'd4273;
      88138:data<=16'd3892;
      88139:data<=16'd3926;
      88140:data<=16'd5627;
      88141:data<=16'd5824;
      88142:data<=16'd5470;
      88143:data<=16'd6352;
      88144:data<=16'd5560;
      88145:data<=16'd5189;
      88146:data<=16'd6678;
      88147:data<=16'd6992;
      88148:data<=16'd7122;
      88149:data<=16'd6721;
      88150:data<=16'd4817;
      88151:data<=16'd4112;
      88152:data<=16'd4769;
      88153:data<=16'd5744;
      88154:data<=16'd5776;
      88155:data<=16'd4822;
      88156:data<=16'd5195;
      88157:data<=16'd5009;
      88158:data<=16'd4931;
      88159:data<=16'd7180;
      88160:data<=16'd7092;
      88161:data<=16'd6655;
      88162:data<=16'd7783;
      88163:data<=16'd5244;
      88164:data<=16'd7304;
      88165:data<=16'd17387;
      88166:data<=16'd21147;
      88167:data<=16'd18989;
      88168:data<=16'd19077;
      88169:data<=16'd18299;
      88170:data<=16'd17086;
      88171:data<=16'd17926;
      88172:data<=16'd18352;
      88173:data<=16'd17434;
      88174:data<=16'd16128;
      88175:data<=16'd15477;
      88176:data<=16'd15018;
      88177:data<=16'd14589;
      88178:data<=16'd15124;
      88179:data<=16'd14957;
      88180:data<=16'd14140;
      88181:data<=16'd13903;
      88182:data<=16'd13039;
      88183:data<=16'd12410;
      88184:data<=16'd11799;
      88185:data<=16'd10619;
      88186:data<=16'd10850;
      88187:data<=16'd10375;
      88188:data<=16'd8619;
      88189:data<=16'd7987;
      88190:data<=16'd6434;
      88191:data<=16'd4686;
      88192:data<=16'd4206;
      88193:data<=16'd3031;
      88194:data<=16'd2843;
      88195:data<=16'd3313;
      88196:data<=16'd2224;
      88197:data<=16'd948;
      88198:data<=-16'd393;
      88199:data<=-16'd124;
      88200:data<=16'd1729;
      88201:data<=16'd1322;
      88202:data<=16'd240;
      88203:data<=-16'd1199;
      88204:data<=-16'd2713;
      88205:data<=-16'd760;
      88206:data<=-16'd2854;
      88207:data<=-16'd11782;
      88208:data<=-16'd16170;
      88209:data<=-16'd16096;
      88210:data<=-16'd16557;
      88211:data<=-16'd15810;
      88212:data<=-16'd15850;
      88213:data<=-16'd16340;
      88214:data<=-16'd15535;
      88215:data<=-16'd16167;
      88216:data<=-16'd16883;
      88217:data<=-16'd16371;
      88218:data<=-16'd16333;
      88219:data<=-16'd15637;
      88220:data<=-16'd14428;
      88221:data<=-16'd14810;
      88222:data<=-16'd16254;
      88223:data<=-16'd16231;
      88224:data<=-16'd14912;
      88225:data<=-16'd14680;
      88226:data<=-16'd14154;
      88227:data<=-16'd13784;
      88228:data<=-16'd15675;
      88229:data<=-16'd15415;
      88230:data<=-16'd13430;
      88231:data<=-16'd13700;
      88232:data<=-16'd12922;
      88233:data<=-16'd12434;
      88234:data<=-16'd14478;
      88235:data<=-16'd14612;
      88236:data<=-16'd13887;
      88237:data<=-16'd13837;
      88238:data<=-16'd12821;
      88239:data<=-16'd12680;
      88240:data<=-16'd13383;
      88241:data<=-16'd13976;
      88242:data<=-16'd13678;
      88243:data<=-16'd12075;
      88244:data<=-16'd12105;
      88245:data<=-16'd11517;
      88246:data<=-16'd10383;
      88247:data<=-16'd13289;
      88248:data<=-16'd11294;
      88249:data<=-16'd2394;
      88250:data<=16'd235;
      88251:data<=-16'd1277;
      88252:data<=-16'd1110;
      88253:data<=-16'd2328;
      88254:data<=-16'd2315;
      88255:data<=-16'd1603;
      88256:data<=-16'd2620;
      88257:data<=-16'd1924;
      88258:data<=-16'd1489;
      88259:data<=-16'd2961;
      88260:data<=-16'd3365;
      88261:data<=-16'd3479;
      88262:data<=-16'd3536;
      88263:data<=-16'd2802;
      88264:data<=-16'd2657;
      88265:data<=-16'd3712;
      88266:data<=-16'd4899;
      88267:data<=-16'd4460;
      88268:data<=-16'd4081;
      88269:data<=-16'd4775;
      88270:data<=-16'd3976;
      88271:data<=-16'd4223;
      88272:data<=-16'd6096;
      88273:data<=-16'd5494;
      88274:data<=-16'd5231;
      88275:data<=-16'd5921;
      88276:data<=-16'd4611;
      88277:data<=-16'd4676;
      88278:data<=-16'd6088;
      88279:data<=-16'd6147;
      88280:data<=-16'd6138;
      88281:data<=-16'd5651;
      88282:data<=-16'd5056;
      88283:data<=-16'd5074;
      88284:data<=-16'd4739;
      88285:data<=-16'd4871;
      88286:data<=-16'd4496;
      88287:data<=-16'd4041;
      88288:data<=-16'd4962;
      88289:data<=-16'd3768;
      88290:data<=-16'd3679;
      88291:data<=-16'd9658;
      88292:data<=-16'd14001;
      88293:data<=-16'd13095;
      88294:data<=-16'd12602;
      88295:data<=-16'd12605;
      88296:data<=-16'd10997;
      88297:data<=-16'd9081;
      88298:data<=-16'd8116;
      88299:data<=-16'd7142;
      88300:data<=-16'd5260;
      88301:data<=-16'd4625;
      88302:data<=-16'd4589;
      88303:data<=-16'd2472;
      88304:data<=-16'd1262;
      88305:data<=-16'd1994;
      88306:data<=-16'd1404;
      88307:data<=-16'd787;
      88308:data<=-16'd1231;
      88309:data<=-16'd5;
      88310:data<=16'd2008;
      88311:data<=16'd1862;
      88312:data<=16'd1375;
      88313:data<=16'd2249;
      88314:data<=16'd1961;
      88315:data<=16'd1876;
      88316:data<=16'd4258;
      88317:data<=16'd4849;
      88318:data<=16'd3814;
      88319:data<=16'd4589;
      88320:data<=16'd4563;
      88321:data<=16'd4722;
      88322:data<=16'd6663;
      88323:data<=16'd6366;
      88324:data<=16'd5548;
      88325:data<=16'd6382;
      88326:data<=16'd6253;
      88327:data<=16'd6516;
      88328:data<=16'd7482;
      88329:data<=16'd7941;
      88330:data<=16'd8592;
      88331:data<=16'd7533;
      88332:data<=16'd8029;
      88333:data<=16'd14929;
      88334:data<=16'd21323;
      88335:data<=16'd21796;
      88336:data<=16'd20618;
      88337:data<=16'd20319;
      88338:data<=16'd19826;
      88339:data<=16'd18762;
      88340:data<=16'd18762;
      88341:data<=16'd19690;
      88342:data<=16'd18976;
      88343:data<=16'd18480;
      88344:data<=16'd19053;
      88345:data<=16'd17541;
      88346:data<=16'd16495;
      88347:data<=16'd17767;
      88348:data<=16'd17573;
      88349:data<=16'd16054;
      88350:data<=16'd14596;
      88351:data<=16'd12794;
      88352:data<=16'd12251;
      88353:data<=16'd13076;
      88354:data<=16'd13318;
      88355:data<=16'd12610;
      88356:data<=16'd12010;
      88357:data<=16'd11829;
      88358:data<=16'd11188;
      88359:data<=16'd11171;
      88360:data<=16'd12025;
      88361:data<=16'd11385;
      88362:data<=16'd10681;
      88363:data<=16'd10904;
      88364:data<=16'd10093;
      88365:data<=16'd10141;
      88366:data<=16'd11106;
      88367:data<=16'd10660;
      88368:data<=16'd10348;
      88369:data<=16'd9676;
      88370:data<=16'd8304;
      88371:data<=16'd8504;
      88372:data<=16'd8831;
      88373:data<=16'd9036;
      88374:data<=16'd8088;
      88375:data<=16'd1444;
      88376:data<=-16'd5524;
      88377:data<=-16'd5553;
      88378:data<=-16'd3627;
      88379:data<=-16'd3554;
      88380:data<=-16'd3416;
      88381:data<=-16'd3686;
      88382:data<=-16'd4034;
      88383:data<=-16'd3465;
      88384:data<=-16'd3550;
      88385:data<=-16'd4449;
      88386:data<=-16'd4557;
      88387:data<=-16'd4126;
      88388:data<=-16'd3856;
      88389:data<=-16'd3601;
      88390:data<=-16'd4511;
      88391:data<=-16'd6187;
      88392:data<=-16'd6144;
      88393:data<=-16'd5747;
      88394:data<=-16'd6208;
      88395:data<=-16'd5732;
      88396:data<=-16'd5937;
      88397:data<=-16'd7336;
      88398:data<=-16'd7348;
      88399:data<=-16'd6998;
      88400:data<=-16'd6492;
      88401:data<=-16'd4916;
      88402:data<=-16'd4720;
      88403:data<=-16'd6056;
      88404:data<=-16'd6902;
      88405:data<=-16'd6825;
      88406:data<=-16'd6234;
      88407:data<=-16'd6228;
      88408:data<=-16'd6122;
      88409:data<=-16'd6261;
      88410:data<=-16'd7952;
      88411:data<=-16'd7823;
      88412:data<=-16'd6608;
      88413:data<=-16'd7359;
      88414:data<=-16'd6464;
      88415:data<=-16'd6586;
      88416:data<=-16'd8739;
      88417:data<=-16'd2913;
      88418:data<=16'd5236;
      88419:data<=16'd4555;
      88420:data<=16'd3230;
      88421:data<=16'd4234;
      88422:data<=16'd1939;
      88423:data<=16'd646;
      88424:data<=16'd1563;
      88425:data<=16'd1111;
      88426:data<=16'd1095;
      88427:data<=16'd1327;
      88428:data<=-16'd58;
      88429:data<=-16'd1309;
      88430:data<=-16'd1162;
      88431:data<=-16'd866;
      88432:data<=-16'd1177;
      88433:data<=-16'd1269;
      88434:data<=-16'd2158;
      88435:data<=-16'd3967;
      88436:data<=-16'd3826;
      88437:data<=-16'd3284;
      88438:data<=-16'd3927;
      88439:data<=-16'd3462;
      88440:data<=-16'd3820;
      88441:data<=-16'd5397;
      88442:data<=-16'd5268;
      88443:data<=-16'd5197;
      88444:data<=-16'd5413;
      88445:data<=-16'd4795;
      88446:data<=-16'd5371;
      88447:data<=-16'd6619;
      88448:data<=-16'd7171;
      88449:data<=-16'd7265;
      88450:data<=-16'd7708;
      88451:data<=-16'd8818;
      88452:data<=-16'd8514;
      88453:data<=-16'd8640;
      88454:data<=-16'd10348;
      88455:data<=-16'd9486;
      88456:data<=-16'd9313;
      88457:data<=-16'd10260;
      88458:data<=-16'd8026;
      88459:data<=-16'd12196;
      88460:data<=-16'd22152;
      88461:data<=-16'd23246;
      88462:data<=-16'd20582;
      88463:data<=-16'd20996;
      88464:data<=-16'd19397;
      88465:data<=-16'd18776;
      88466:data<=-16'd20095;
      88467:data<=-16'd19144;
      88468:data<=-16'd18163;
      88469:data<=-16'd17872;
      88470:data<=-16'd17014;
      88471:data<=-16'd16472;
      88472:data<=-16'd16478;
      88473:data<=-16'd16565;
      88474:data<=-16'd15477;
      88475:data<=-16'd14472;
      88476:data<=-16'd14522;
      88477:data<=-16'd13347;
      88478:data<=-16'd12627;
      88479:data<=-16'd13244;
      88480:data<=-16'd12703;
      88481:data<=-16'd12204;
      88482:data<=-16'd11928;
      88483:data<=-16'd11144;
      88484:data<=-16'd10627;
      88485:data<=-16'd9568;
      88486:data<=-16'd9057;
      88487:data<=-16'd8617;
      88488:data<=-16'd6848;
      88489:data<=-16'd6639;
      88490:data<=-16'd6338;
      88491:data<=-16'd4209;
      88492:data<=-16'd3659;
      88493:data<=-16'd3216;
      88494:data<=-16'd2112;
      88495:data<=-16'd1912;
      88496:data<=-16'd1108;
      88497:data<=-16'd67;
      88498:data<=16'd1814;
      88499:data<=16'd2887;
      88500:data<=16'd1662;
      88501:data<=16'd6977;
      88502:data<=16'd16428;
      88503:data<=16'd18315;
      88504:data<=16'd17979;
      88505:data<=16'd18729;
      88506:data<=16'd16874;
      88507:data<=16'd16965;
      88508:data<=16'd17243;
      88509:data<=16'd15747;
      88510:data<=16'd17462;
      88511:data<=16'd18383;
      88512:data<=16'd16901;
      88513:data<=16'd17114;
      88514:data<=16'd16284;
      88515:data<=16'd15306;
      88516:data<=16'd16772;
      88517:data<=16'd17139;
      88518:data<=16'd16274;
      88519:data<=16'd15970;
      88520:data<=16'd15487;
      88521:data<=16'd15001;
      88522:data<=16'd15361;
      88523:data<=16'd16110;
      88524:data<=16'd15330;
      88525:data<=16'd14214;
      88526:data<=16'd14531;
      88527:data<=16'd13929;
      88528:data<=16'd13879;
      88529:data<=16'd15643;
      88530:data<=16'd15068;
      88531:data<=16'd13790;
      88532:data<=16'd13913;
      88533:data<=16'd13019;
      88534:data<=16'd13147;
      88535:data<=16'd14534;
      88536:data<=16'd14270;
      88537:data<=16'd13474;
      88538:data<=16'd13197;
      88539:data<=16'd13066;
      88540:data<=16'd12242;
      88541:data<=16'd12229;
      88542:data<=16'd14239;
      88543:data<=16'd10704;
      88544:data<=16'd2314;
      88545:data<=16'd576;
      88546:data<=16'd2062;
      88547:data<=16'd1542;
      88548:data<=16'd3287;
      88549:data<=16'd3835;
      88550:data<=16'd2616;
      88551:data<=16'd3612;
      88552:data<=16'd2990;
      88553:data<=16'd2265;
      88554:data<=16'd4291;
      88555:data<=16'd4666;
      88556:data<=16'd4194;
      88557:data<=16'd4511;
      88558:data<=16'd4099;
      88559:data<=16'd4340;
      88560:data<=16'd5115;
      88561:data<=16'd5473;
      88562:data<=16'd5325;
      88563:data<=16'd4702;
      88564:data<=16'd5289;
      88565:data<=16'd6119;
      88566:data<=16'd6109;
      88567:data<=16'd6370;
      88568:data<=16'd5891;
      88569:data<=16'd5676;
      88570:data<=16'd6147;
      88571:data<=16'd5262;
      88572:data<=16'd5541;
      88573:data<=16'd7166;
      88574:data<=16'd7036;
      88575:data<=16'd6552;
      88576:data<=16'd6185;
      88577:data<=16'd5398;
      88578:data<=16'd5724;
      88579:data<=16'd7224;
      88580:data<=16'd8064;
      88581:data<=16'd6789;
      88582:data<=16'd6231;
      88583:data<=16'd6602;
      88584:data<=16'd4469;
      88585:data<=16'd6798;
      88586:data<=16'd14598;
      88587:data<=16'd15505;
      88588:data<=16'd12763;
      88589:data<=16'd13762;
      88590:data<=16'd12710;
      88591:data<=16'd10182;
      88592:data<=16'd9254;
      88593:data<=16'd8085;
      88594:data<=16'd7884;
      88595:data<=16'd7890;
      88596:data<=16'd7194;
      88597:data<=16'd6398;
      88598:data<=16'd4476;
      88599:data<=16'd3603;
      88600:data<=16'd3656;
      88601:data<=16'd2799;
      88602:data<=16'd3045;
      88603:data<=16'd2599;
      88604:data<=16'd652;
      88605:data<=16'd17;
      88606:data<=-16'd705;
      88607:data<=-16'd1395;
      88608:data<=-16'd972;
      88609:data<=-16'd1398;
      88610:data<=-16'd2582;
      88611:data<=-16'd3548;
      88612:data<=-16'd3606;
      88613:data<=-16'd3523;
      88614:data<=-16'd4350;
      88615:data<=-16'd4181;
      88616:data<=-16'd4628;
      88617:data<=-16'd6335;
      88618:data<=-16'd6018;
      88619:data<=-16'd6314;
      88620:data<=-16'd7062;
      88621:data<=-16'd5799;
      88622:data<=-16'd6771;
      88623:data<=-16'd8526;
      88624:data<=-16'd8592;
      88625:data<=-16'd8862;
      88626:data<=-16'd7602;
      88627:data<=-16'd9724;
      88628:data<=-16'd17346;
      88629:data<=-16'd20403;
      88630:data<=-16'd19378;
      88631:data<=-16'd19328;
      88632:data<=-16'd18034;
      88633:data<=-16'd17123;
      88634:data<=-16'd17352;
      88635:data<=-16'd17845;
      88636:data<=-16'd19112;
      88637:data<=-16'd18437;
      88638:data<=-16'd17268;
      88639:data<=-16'd17330;
      88640:data<=-16'd16078;
      88641:data<=-16'd16046;
      88642:data<=-16'd17358;
      88643:data<=-16'd16725;
      88644:data<=-16'd16343;
      88645:data<=-16'd16076;
      88646:data<=-16'd14690;
      88647:data<=-16'd14692;
      88648:data<=-16'd15427;
      88649:data<=-16'd15282;
      88650:data<=-16'd15038;
      88651:data<=-16'd14596;
      88652:data<=-16'd13452;
      88653:data<=-16'd13001;
      88654:data<=-16'd14368;
      88655:data<=-16'd14650;
      88656:data<=-16'd13039;
      88657:data<=-16'd12759;
      88658:data<=-16'd12587;
      88659:data<=-16'd11835;
      88660:data<=-16'd12472;
      88661:data<=-16'd12348;
      88662:data<=-16'd11632;
      88663:data<=-16'd11900;
      88664:data<=-16'd11218;
      88665:data<=-16'd10308;
      88666:data<=-16'd9885;
      88667:data<=-16'd10536;
      88668:data<=-16'd12419;
      88669:data<=-16'd8589;
      88670:data<=16'd3;
      88671:data<=16'd2475;
      88672:data<=16'd390;
      88673:data<=-16'd182;
      88674:data<=-16'd717;
      88675:data<=-16'd864;
      88676:data<=-16'd306;
      88677:data<=-16'd459;
      88678:data<=-16'd629;
      88679:data<=-16'd1287;
      88680:data<=-16'd1996;
      88681:data<=-16'd1427;
      88682:data<=-16'd1262;
      88683:data<=-16'd1823;
      88684:data<=-16'd1726;
      88685:data<=-16'd1354;
      88686:data<=-16'd1130;
      88687:data<=-16'd854;
      88688:data<=-16'd491;
      88689:data<=-16'd557;
      88690:data<=-16'd989;
      88691:data<=-16'd126;
      88692:data<=16'd1577;
      88693:data<=16'd2035;
      88694:data<=16'd1859;
      88695:data<=16'd1718;
      88696:data<=16'd1307;
      88697:data<=16'd1997;
      88698:data<=16'd3654;
      88699:data<=16'd3852;
      88700:data<=16'd3201;
      88701:data<=16'd3698;
      88702:data<=16'd3694;
      88703:data<=16'd3124;
      88704:data<=16'd4687;
      88705:data<=16'd5742;
      88706:data<=16'd4616;
      88707:data<=16'd5069;
      88708:data<=16'd5068;
      88709:data<=16'd3889;
      88710:data<=16'd6046;
      88711:data<=16'd4986;
      88712:data<=-16'd2554;
      88713:data<=-16'd5275;
      88714:data<=-16'd3450;
      88715:data<=-16'd4118;
      88716:data<=-16'd3153;
      88717:data<=-16'd629;
      88718:data<=-16'd567;
      88719:data<=-16'd526;
      88720:data<=-16'd379;
      88721:data<=-16'd983;
      88722:data<=-16'd114;
      88723:data<=16'd1525;
      88724:data<=16'd2015;
      88725:data<=16'd1720;
      88726:data<=16'd1601;
      88727:data<=16'd1538;
      88728:data<=16'd1645;
      88729:data<=16'd2993;
      88730:data<=16'd3786;
      88731:data<=16'd2983;
      88732:data<=16'd3539;
      88733:data<=16'd4229;
      88734:data<=16'd3174;
      88735:data<=16'd3888;
      88736:data<=16'd6094;
      88737:data<=16'd6460;
      88738:data<=16'd6014;
      88739:data<=16'd5609;
      88740:data<=16'd4608;
      88741:data<=16'd5060;
      88742:data<=16'd7453;
      88743:data<=16'd7988;
      88744:data<=16'd6802;
      88745:data<=16'd6893;
      88746:data<=16'd6531;
      88747:data<=16'd6551;
      88748:data<=16'd8652;
      88749:data<=16'd8404;
      88750:data<=16'd7409;
      88751:data<=16'd8088;
      88752:data<=16'd6310;
      88753:data<=16'd8125;
      88754:data<=16'd16548;
      88755:data<=16'd19787;
      88756:data<=16'd17732;
      88757:data<=16'd17462;
      88758:data<=16'd16471;
      88759:data<=16'd15277;
      88760:data<=16'd16240;
      88761:data<=16'd16977;
      88762:data<=16'd16698;
      88763:data<=16'd15879;
      88764:data<=16'd15139;
      88765:data<=16'd14672;
      88766:data<=16'd14131;
      88767:data<=16'd14411;
      88768:data<=16'd14492;
      88769:data<=16'd13452;
      88770:data<=16'd12698;
      88771:data<=16'd12255;
      88772:data<=16'd12316;
      88773:data<=16'd12631;
      88774:data<=16'd11955;
      88775:data<=16'd11223;
      88776:data<=16'd10837;
      88777:data<=16'd10633;
      88778:data<=16'd10775;
      88779:data<=16'd10646;
      88780:data<=16'd10939;
      88781:data<=16'd10722;
      88782:data<=16'd9188;
      88783:data<=16'd9003;
      88784:data<=16'd9060;
      88785:data<=16'd7803;
      88786:data<=16'd7168;
      88787:data<=16'd6398;
      88788:data<=16'd5504;
      88789:data<=16'd5216;
      88790:data<=16'd4572;
      88791:data<=16'd4202;
      88792:data<=16'd2582;
      88793:data<=16'd743;
      88794:data<=16'd1842;
      88795:data<=-16'd400;
      88796:data<=-16'd7347;
      88797:data<=-16'd10549;
      88798:data<=-16'd10771;
      88799:data<=-16'd11605;
      88800:data<=-16'd11577;
      88801:data<=-16'd11186;
      88802:data<=-16'd10657;
      88803:data<=-16'd10375;
      88804:data<=-16'd11339;
      88805:data<=-16'd12188;
      88806:data<=-16'd12525;
      88807:data<=-16'd12387;
      88808:data<=-16'd11759;
      88809:data<=-16'd11391;
      88810:data<=-16'd11336;
      88811:data<=-16'd12322;
      88812:data<=-16'd12933;
      88813:data<=-16'd11920;
      88814:data<=-16'd11926;
      88815:data<=-16'd11731;
      88816:data<=-16'd10749;
      88817:data<=-16'd12002;
      88818:data<=-16'd12613;
      88819:data<=-16'd11888;
      88820:data<=-16'd12242;
      88821:data<=-16'd11098;
      88822:data<=-16'd10293;
      88823:data<=-16'd11891;
      88824:data<=-16'd12208;
      88825:data<=-16'd11906;
      88826:data<=-16'd11911;
      88827:data<=-16'd11069;
      88828:data<=-16'd10598;
      88829:data<=-16'd10608;
      88830:data<=-16'd11623;
      88831:data<=-16'd12252;
      88832:data<=-16'd10819;
      88833:data<=-16'd10671;
      88834:data<=-16'd10308;
      88835:data<=-16'd9592;
      88836:data<=-16'd12669;
      88837:data<=-16'd10922;
      88838:data<=-16'd2106;
      88839:data<=16'd1007;
      88840:data<=-16'd438;
      88841:data<=-16'd694;
      88842:data<=-16'd2217;
      88843:data<=-16'd2581;
      88844:data<=-16'd1626;
      88845:data<=-16'd2134;
      88846:data<=-16'd1992;
      88847:data<=-16'd1874;
      88848:data<=-16'd2963;
      88849:data<=-16'd3797;
      88850:data<=-16'd4070;
      88851:data<=-16'd3460;
      88852:data<=-16'd3046;
      88853:data<=-16'd3133;
      88854:data<=-16'd3366;
      88855:data<=-16'd5060;
      88856:data<=-16'd5497;
      88857:data<=-16'd4117;
      88858:data<=-16'd4498;
      88859:data<=-16'd4361;
      88860:data<=-16'd3806;
      88861:data<=-16'd5438;
      88862:data<=-16'd5636;
      88863:data<=-16'd4698;
      88864:data<=-16'd5053;
      88865:data<=-16'd4696;
      88866:data<=-16'd4628;
      88867:data<=-16'd5739;
      88868:data<=-16'd6172;
      88869:data<=-16'd5824;
      88870:data<=-16'd5456;
      88871:data<=-16'd5715;
      88872:data<=-16'd5665;
      88873:data<=-16'd5894;
      88874:data<=-16'd7444;
      88875:data<=-16'd6584;
      88876:data<=-16'd5031;
      88877:data<=-16'd5671;
      88878:data<=-16'd4018;
      88879:data<=-16'd5488;
      88880:data<=-16'd13900;
      88881:data<=-16'd17094;
      88882:data<=-16'd14669;
      88883:data<=-16'd14728;
      88884:data<=-16'd14483;
      88885:data<=-16'd13676;
      88886:data<=-16'd13737;
      88887:data<=-16'd12395;
      88888:data<=-16'd11412;
      88889:data<=-16'd11242;
      88890:data<=-16'd10528;
      88891:data<=-16'd9779;
      88892:data<=-16'd8105;
      88893:data<=-16'd6414;
      88894:data<=-16'd6026;
      88895:data<=-16'd5758;
      88896:data<=-16'd5630;
      88897:data<=-16'd5359;
      88898:data<=-16'd4300;
      88899:data<=-16'd3013;
      88900:data<=-16'd1783;
      88901:data<=-16'd1172;
      88902:data<=-16'd1227;
      88903:data<=-16'd1527;
      88904:data<=-16'd1034;
      88905:data<=16'd1304;
      88906:data<=16'd2813;
      88907:data<=16'd2661;
      88908:data<=16'd3107;
      88909:data<=16'd2678;
      88910:data<=16'd2361;
      88911:data<=16'd4346;
      88912:data<=16'd5324;
      88913:data<=16'd5101;
      88914:data<=16'd5309;
      88915:data<=16'd4830;
      88916:data<=16'd4898;
      88917:data<=16'd5736;
      88918:data<=16'd6692;
      88919:data<=16'd7586;
      88920:data<=16'd6708;
      88921:data<=16'd7877;
      88922:data<=16'd13603;
      88923:data<=16'd17653;
      88924:data<=16'd18457;
      88925:data<=16'd18181;
      88926:data<=16'd16947;
      88927:data<=16'd16866;
      88928:data<=16'd16982;
      88929:data<=16'd16462;
      88930:data<=16'd17555;
      88931:data<=16'd17585;
      88932:data<=16'd16195;
      88933:data<=16'd16390;
      88934:data<=16'd15932;
      88935:data<=16'd15291;
      88936:data<=16'd16675;
      88937:data<=16'd17124;
      88938:data<=16'd16299;
      88939:data<=16'd16114;
      88940:data<=16'd15706;
      88941:data<=16'd14944;
      88942:data<=16'd14919;
      88943:data<=16'd15587;
      88944:data<=16'd15462;
      88945:data<=16'd14424;
      88946:data<=16'd13860;
      88947:data<=16'd13562;
      88948:data<=16'd13911;
      88949:data<=16'd14671;
      88950:data<=16'd13803;
      88951:data<=16'd12866;
      88952:data<=16'd12739;
      88953:data<=16'd11913;
      88954:data<=16'd12192;
      88955:data<=16'd13254;
      88956:data<=16'd12854;
      88957:data<=16'd12000;
      88958:data<=16'd11232;
      88959:data<=16'd11171;
      88960:data<=16'd11318;
      88961:data<=16'd10806;
      88962:data<=16'd12058;
      88963:data<=16'd10931;
      88964:data<=16'd3489;
      88965:data<=-16'd1196;
      88966:data<=16'd2;
      88967:data<=16'd879;
      88968:data<=16'd1183;
      88969:data<=16'd977;
      88970:data<=16'd82;
      88971:data<=16'd469;
      88972:data<=16'd928;
      88973:data<=16'd1707;
      88974:data<=16'd2801;
      88975:data<=16'd2002;
      88976:data<=16'd1471;
      88977:data<=16'd1959;
      88978:data<=16'd1861;
      88979:data<=16'd2608;
      88980:data<=16'd3472;
      88981:data<=16'd3196;
      88982:data<=16'd2958;
      88983:data<=16'd2799;
      88984:data<=16'd2861;
      88985:data<=16'd2886;
      88986:data<=16'd2393;
      88987:data<=16'd2164;
      88988:data<=16'd1569;
      88989:data<=16'd690;
      88990:data<=16'd878;
      88991:data<=16'd1318;
      88992:data<=16'd605;
      88993:data<=-16'd1168;
      88994:data<=-16'd1982;
      88995:data<=-16'd1457;
      88996:data<=-16'd1491;
      88997:data<=-16'd1350;
      88998:data<=-16'd1918;
      88999:data<=-16'd4153;
      89000:data<=-16'd4191;
      89001:data<=-16'd3345;
      89002:data<=-16'd3683;
      89003:data<=-16'd2645;
      89004:data<=-16'd3777;
      89005:data<=-16'd5345;
      89006:data<=16'd202;
      89007:data<=16'd5577;
      89008:data<=16'd4874;
      89009:data<=16'd4617;
      89010:data<=16'd4678;
      89011:data<=16'd2732;
      89012:data<=16'd1996;
      89013:data<=16'd2032;
      89014:data<=16'd1027;
      89015:data<=16'd754;
      89016:data<=16'd1762;
      89017:data<=16'd1122;
      89018:data<=-16'd1142;
      89019:data<=-16'd1554;
      89020:data<=-16'd1465;
      89021:data<=-16'd2256;
      89022:data<=-16'd1865;
      89023:data<=-16'd2478;
      89024:data<=-16'd4282;
      89025:data<=-16'd4055;
      89026:data<=-16'd4059;
      89027:data<=-16'd5062;
      89028:data<=-16'd4780;
      89029:data<=-16'd4546;
      89030:data<=-16'd5077;
      89031:data<=-16'd5601;
      89032:data<=-16'd5817;
      89033:data<=-16'd5676;
      89034:data<=-16'd5724;
      89035:data<=-16'd5550;
      89036:data<=-16'd6322;
      89037:data<=-16'd8055;
      89038:data<=-16'd7216;
      89039:data<=-16'd6167;
      89040:data<=-16'd7268;
      89041:data<=-16'd6996;
      89042:data<=-16'd7127;
      89043:data<=-16'd8534;
      89044:data<=-16'd8255;
      89045:data<=-16'd8651;
      89046:data<=-16'd8551;
      89047:data<=-16'd7715;
      89048:data<=-16'd13265;
      89049:data<=-16'd20205;
      89050:data<=-16'd20011;
      89051:data<=-16'd18507;
      89052:data<=-16'd18483;
      89053:data<=-16'd17171;
      89054:data<=-16'd17308;
      89055:data<=-16'd18516;
      89056:data<=-16'd17849;
      89057:data<=-16'd16835;
      89058:data<=-16'd16269;
      89059:data<=-16'd15629;
      89060:data<=-16'd15729;
      89061:data<=-16'd16368;
      89062:data<=-16'd16311;
      89063:data<=-16'd15443;
      89064:data<=-16'd14600;
      89065:data<=-16'd13775;
      89066:data<=-16'd13288;
      89067:data<=-16'd14211;
      89068:data<=-16'd14642;
      89069:data<=-16'd13217;
      89070:data<=-16'd12610;
      89071:data<=-16'd12483;
      89072:data<=-16'd11086;
      89073:data<=-16'd11168;
      89074:data<=-16'd12828;
      89075:data<=-16'd12627;
      89076:data<=-16'd11342;
      89077:data<=-16'd10913;
      89078:data<=-16'd10379;
      89079:data<=-16'd9758;
      89080:data<=-16'd10337;
      89081:data<=-16'd10859;
      89082:data<=-16'd9750;
      89083:data<=-16'd8668;
      89084:data<=-16'd8510;
      89085:data<=-16'd8149;
      89086:data<=-16'd7294;
      89087:data<=-16'd5871;
      89088:data<=-16'd5598;
      89089:data<=-16'd5721;
      89090:data<=-16'd602;
      89091:data<=16'd6056;
      89092:data<=16'd6883;
      89093:data<=16'd6749;
      89094:data<=16'd8003;
      89095:data<=16'd7081;
      89096:data<=16'd6655;
      89097:data<=16'd7171;
      89098:data<=16'd7460;
      89099:data<=16'd9156;
      89100:data<=16'd9726;
      89101:data<=16'd9074;
      89102:data<=16'd9307;
      89103:data<=16'd8478;
      89104:data<=16'd8167;
      89105:data<=16'd9544;
      89106:data<=16'd9884;
      89107:data<=16'd9840;
      89108:data<=16'd9735;
      89109:data<=16'd9021;
      89110:data<=16'd8786;
      89111:data<=16'd9136;
      89112:data<=16'd10396;
      89113:data<=16'd11066;
      89114:data<=16'd10079;
      89115:data<=16'd9790;
      89116:data<=16'd9558;
      89117:data<=16'd9342;
      89118:data<=16'd10937;
      89119:data<=16'd11679;
      89120:data<=16'd10880;
      89121:data<=16'd10383;
      89122:data<=16'd9899;
      89123:data<=16'd10003;
      89124:data<=16'd10884;
      89125:data<=16'd11878;
      89126:data<=16'd11445;
      89127:data<=16'd9727;
      89128:data<=16'd10263;
      89129:data<=16'd10554;
      89130:data<=16'd9492;
      89131:data<=16'd10877;
      89132:data<=16'd7834;
      89133:data<=16'd584;
      89134:data<=-16'd42;
      89135:data<=16'd836;
      89136:data<=-16'd106;
      89137:data<=16'd1833;
      89138:data<=16'd1394;
      89139:data<=16'd190;
      89140:data<=16'd2243;
      89141:data<=16'd2102;
      89142:data<=16'd1885;
      89143:data<=16'd3001;
      89144:data<=16'd2265;
      89145:data<=16'd2813;
      89146:data<=16'd3504;
      89147:data<=16'd2719;
      89148:data<=16'd3576;
      89149:data<=16'd4672;
      89150:data<=16'd5221;
      89151:data<=16'd5445;
      89152:data<=16'd4911;
      89153:data<=16'd5101;
      89154:data<=16'd4854;
      89155:data<=16'd5194;
      89156:data<=16'd6684;
      89157:data<=16'd5488;
      89158:data<=16'd4728;
      89159:data<=16'd5870;
      89160:data<=16'd4842;
      89161:data<=16'd4454;
      89162:data<=16'd5477;
      89163:data<=16'd5732;
      89164:data<=16'd6575;
      89165:data<=16'd6517;
      89166:data<=16'd5471;
      89167:data<=16'd5456;
      89168:data<=16'd6496;
      89169:data<=16'd7705;
      89170:data<=16'd6466;
      89171:data<=16'd5727;
      89172:data<=16'd6699;
      89173:data<=16'd4913;
      89174:data<=16'd8369;
      89175:data<=16'd17385;
      89176:data<=16'd17697;
      89177:data<=16'd14716;
      89178:data<=16'd15347;
      89179:data<=16'd13706;
      89180:data<=16'd13547;
      89181:data<=16'd14784;
      89182:data<=16'd13364;
      89183:data<=16'd13362;
      89184:data<=16'd13048;
      89185:data<=16'd12091;
      89186:data<=16'd12633;
      89187:data<=16'd10912;
      89188:data<=16'd9840;
      89189:data<=16'd10671;
      89190:data<=16'd9873;
      89191:data<=16'd10207;
      89192:data<=16'd9536;
      89193:data<=16'd6549;
      89194:data<=16'd5780;
      89195:data<=16'd4444;
      89196:data<=16'd2787;
      89197:data<=16'd3938;
      89198:data<=16'd3626;
      89199:data<=16'd1243;
      89200:data<=-16'd613;
      89201:data<=-16'd1052;
      89202:data<=16'd30;
      89203:data<=-16'd171;
      89204:data<=-16'd1298;
      89205:data<=-16'd2234;
      89206:data<=-16'd3900;
      89207:data<=-16'd3850;
      89208:data<=-16'd3148;
      89209:data<=-16'd3617;
      89210:data<=-16'd3436;
      89211:data<=-16'd4438;
      89212:data<=-16'd6111;
      89213:data<=-16'd6822;
      89214:data<=-16'd7168;
      89215:data<=-16'd5438;
      89216:data<=-16'd7641;
      89217:data<=-16'd15723;
      89218:data<=-16'd18069;
      89219:data<=-16'd16384;
      89220:data<=-16'd17117;
      89221:data<=-16'd15902;
      89222:data<=-16'd15341;
      89223:data<=-16'd16759;
      89224:data<=-16'd16116;
      89225:data<=-16'd16472;
      89226:data<=-16'd16889;
      89227:data<=-16'd15528;
      89228:data<=-16'd15778;
      89229:data<=-16'd15784;
      89230:data<=-16'd15655;
      89231:data<=-16'd16824;
      89232:data<=-16'd15646;
      89233:data<=-16'd14586;
      89234:data<=-16'd16128;
      89235:data<=-16'd16083;
      89236:data<=-16'd15286;
      89237:data<=-16'd15941;
      89238:data<=-16'd15975;
      89239:data<=-16'd15553;
      89240:data<=-16'd15245;
      89241:data<=-16'd13796;
      89242:data<=-16'd13107;
      89243:data<=-16'd14862;
      89244:data<=-16'd15188;
      89245:data<=-16'd13082;
      89246:data<=-16'd12684;
      89247:data<=-16'd13245;
      89248:data<=-16'd12910;
      89249:data<=-16'd13230;
      89250:data<=-16'd13236;
      89251:data<=-16'd12524;
      89252:data<=-16'd11969;
      89253:data<=-16'd11150;
      89254:data<=-16'd11304;
      89255:data<=-16'd11671;
      89256:data<=-16'd11711;
      89257:data<=-16'd12442;
      89258:data<=-16'd8860;
      89259:data<=-16'd1525;
      89260:data<=16'd1096;
      89261:data<=16'd332;
      89262:data<=-16'd400;
      89263:data<=-16'd2275;
      89264:data<=-16'd2510;
      89265:data<=-16'd1043;
      89266:data<=-16'd660;
      89267:data<=-16'd925;
      89268:data<=-16'd2200;
      89269:data<=-16'd3177;
      89270:data<=-16'd2299;
      89271:data<=-16'd1723;
      89272:data<=-16'd1572;
      89273:data<=-16'd1548;
      89274:data<=-16'd2387;
      89275:data<=-16'd2664;
      89276:data<=-16'd2801;
      89277:data<=-16'd3610;
      89278:data<=-16'd3378;
      89279:data<=-16'd2532;
      89280:data<=-16'd2984;
      89281:data<=-16'd4290;
      89282:data<=-16'd4300;
      89283:data<=-16'd2872;
      89284:data<=-16'd2488;
      89285:data<=-16'd3513;
      89286:data<=-16'd4132;
      89287:data<=-16'd3242;
      89288:data<=-16'd1566;
      89289:data<=-16'd1574;
      89290:data<=-16'd2105;
      89291:data<=-16'd970;
      89292:data<=-16'd144;
      89293:data<=16'd1036;
      89294:data<=16'd2461;
      89295:data<=16'd1553;
      89296:data<=16'd2144;
      89297:data<=16'd3703;
      89298:data<=16'd2476;
      89299:data<=16'd3588;
      89300:data<=16'd3595;
      89301:data<=-16'd3186;
      89302:data<=-16'd6232;
      89303:data<=-16'd3979;
      89304:data<=-16'd4349;
      89305:data<=-16'd3345;
      89306:data<=-16'd581;
      89307:data<=-16'd429;
      89308:data<=-16'd97;
      89309:data<=-16'd20;
      89310:data<=-16'd978;
      89311:data<=16'd220;
      89312:data<=16'd1832;
      89313:data<=16'd2146;
      89314:data<=16'd2863;
      89315:data<=16'd3782;
      89316:data<=16'd3924;
      89317:data<=16'd3557;
      89318:data<=16'd4103;
      89319:data<=16'd4830;
      89320:data<=16'd4077;
      89321:data<=16'd4458;
      89322:data<=16'd5952;
      89323:data<=16'd5474;
      89324:data<=16'd5533;
      89325:data<=16'd7022;
      89326:data<=16'd6965;
      89327:data<=16'd6925;
      89328:data<=16'd7755;
      89329:data<=16'd7451;
      89330:data<=16'd7746;
      89331:data<=16'd9415;
      89332:data<=16'd9379;
      89333:data<=16'd8072;
      89334:data<=16'd7808;
      89335:data<=16'd7280;
      89336:data<=16'd7028;
      89337:data<=16'd8904;
      89338:data<=16'd10084;
      89339:data<=16'd9711;
      89340:data<=16'd9298;
      89341:data<=16'd8241;
      89342:data<=16'd10878;
      89343:data<=16'd18298;
      89344:data<=16'd21144;
      89345:data<=16'd19105;
      89346:data<=16'd19052;
      89347:data<=16'd18572;
      89348:data<=16'd16865;
      89349:data<=16'd17757;
      89350:data<=16'd18766;
      89351:data<=16'd17655;
      89352:data<=16'd16728;
      89353:data<=16'd16284;
      89354:data<=16'd15808;
      89355:data<=16'd16266;
      89356:data<=16'd16989;
      89357:data<=16'd16410;
      89358:data<=16'd15279;
      89359:data<=16'd14882;
      89360:data<=16'd14792;
      89361:data<=16'd14292;
      89362:data<=16'd13547;
      89363:data<=16'd13320;
      89364:data<=16'd13496;
      89365:data<=16'd13534;
      89366:data<=16'd13480;
      89367:data<=16'd12533;
      89368:data<=16'd11735;
      89369:data<=16'd12560;
      89370:data<=16'd12070;
      89371:data<=16'd10813;
      89372:data<=16'd11160;
      89373:data<=16'd9794;
      89374:data<=16'd8913;
      89375:data<=16'd11297;
      89376:data<=16'd11327;
      89377:data<=16'd10317;
      89378:data<=16'd10883;
      89379:data<=16'd9360;
      89380:data<=16'd8757;
      89381:data<=16'd9347;
      89382:data<=16'd7982;
      89383:data<=16'd8722;
      89384:data<=16'd7272;
      89385:data<=-16'd466;
      89386:data<=-16'd4501;
      89387:data<=-16'd3936;
      89388:data<=-16'd4112;
      89389:data<=-16'd2682;
      89390:data<=-16'd2083;
      89391:data<=-16'd3542;
      89392:data<=-16'd2931;
      89393:data<=-16'd3137;
      89394:data<=-16'd5163;
      89395:data<=-16'd5583;
      89396:data<=-16'd6108;
      89397:data<=-16'd6256;
      89398:data<=-16'd4687;
      89399:data<=-16'd5503;
      89400:data<=-16'd8079;
      89401:data<=-16'd8602;
      89402:data<=-16'd8737;
      89403:data<=-16'd8705;
      89404:data<=-16'd7048;
      89405:data<=-16'd6645;
      89406:data<=-16'd8363;
      89407:data<=-16'd9174;
      89408:data<=-16'd8895;
      89409:data<=-16'd9423;
      89410:data<=-16'd10125;
      89411:data<=-16'd9260;
      89412:data<=-16'd8658;
      89413:data<=-16'd9881;
      89414:data<=-16'd9820;
      89415:data<=-16'd8821;
      89416:data<=-16'd9367;
      89417:data<=-16'd9110;
      89418:data<=-16'd9042;
      89419:data<=-16'd11580;
      89420:data<=-16'd14731;
      89421:data<=-16'd17964;
      89422:data<=-16'd18484;
      89423:data<=-16'd16054;
      89424:data<=-16'd17092;
      89425:data<=-16'd18263;
      89426:data<=-16'd16718;
      89427:data<=-16'd17653;
      89428:data<=-16'd14477;
      89429:data<=-16'd5315;
      89430:data<=-16'd1501;
      89431:data<=-16'd1139;
      89432:data<=16'd1063;
      89433:data<=16'd1826;
      89434:data<=16'd1600;
      89435:data<=16'd1721;
      89436:data<=16'd2238;
      89437:data<=16'd2725;
      89438:data<=16'd2320;
      89439:data<=16'd2760;
      89440:data<=16'd2218;
      89441:data<=16'd811;
      89442:data<=16'd1838;
      89443:data<=16'd1477;
      89444:data<=16'd2819;
      89445:data<=16'd10151;
      89446:data<=16'd13218;
      89447:data<=16'd10830;
      89448:data<=16'd9849;
      89449:data<=16'd9007;
      89450:data<=16'd9062;
      89451:data<=16'd8939;
      89452:data<=16'd7498;
      89453:data<=16'd8032;
      89454:data<=16'd7454;
      89455:data<=16'd6664;
      89456:data<=16'd6790;
      89457:data<=-16'd453;
      89458:data<=-16'd11154;
      89459:data<=-16'd17127;
      89460:data<=-16'd20177;
      89461:data<=-16'd19676;
      89462:data<=-16'd18342;
      89463:data<=-16'd19036;
      89464:data<=-16'd17920;
      89465:data<=-16'd16657;
      89466:data<=-16'd16120;
      89467:data<=-16'd14851;
      89468:data<=-16'd14885;
      89469:data<=-16'd14226;
      89470:data<=-16'd13203;
      89471:data<=-16'd14061;
      89472:data<=-16'd14205;
      89473:data<=-16'd13292;
      89474:data<=-16'd12172;
      89475:data<=-16'd15465;
      89476:data<=-16'd24864;
      89477:data<=-16'd28665;
      89478:data<=-16'd26069;
      89479:data<=-16'd25840;
      89480:data<=-16'd25205;
      89481:data<=-16'd24380;
      89482:data<=-16'd24118;
      89483:data<=-16'd21024;
      89484:data<=-16'd20274;
      89485:data<=-16'd21840;
      89486:data<=-16'd21152;
      89487:data<=-16'd20698;
      89488:data<=-16'd19411;
      89489:data<=-16'd17346;
      89490:data<=-16'd17479;
      89491:data<=-16'd17494;
      89492:data<=-16'd16231;
      89493:data<=-16'd14164;
      89494:data<=-16'd13071;
      89495:data<=-16'd13564;
      89496:data<=-16'd11544;
      89497:data<=-16'd9834;
      89498:data<=-16'd11741;
      89499:data<=-16'd12528;
      89500:data<=-16'd11909;
      89501:data<=-16'd11097;
      89502:data<=-16'd9705;
      89503:data<=-16'd8739;
      89504:data<=-16'd7682;
      89505:data<=-16'd8381;
      89506:data<=-16'd9031;
      89507:data<=-16'd6625;
      89508:data<=-16'd5571;
      89509:data<=-16'd4352;
      89510:data<=-16'd3362;
      89511:data<=-16'd6476;
      89512:data<=-16'd4449;
      89513:data<=16'd1397;
      89514:data<=16'd2015;
      89515:data<=16'd3231;
      89516:data<=16'd4182;
      89517:data<=16'd3148;
      89518:data<=16'd3935;
      89519:data<=16'd2734;
      89520:data<=16'd8069;
      89521:data<=16'd21416;
      89522:data<=16'd23928;
      89523:data<=16'd20563;
      89524:data<=16'd21191;
      89525:data<=16'd18480;
      89526:data<=16'd16666;
      89527:data<=16'd17741;
      89528:data<=16'd16763;
      89529:data<=16'd17202;
      89530:data<=16'd17048;
      89531:data<=16'd15393;
      89532:data<=16'd15817;
      89533:data<=16'd15380;
      89534:data<=16'd14868;
      89535:data<=16'd15356;
      89536:data<=16'd14604;
      89537:data<=16'd13549;
      89538:data<=16'd10944;
      89539:data<=16'd8933;
      89540:data<=16'd10026;
      89541:data<=16'd9420;
      89542:data<=16'd8375;
      89543:data<=16'd8886;
      89544:data<=16'd7982;
      89545:data<=16'd8220;
      89546:data<=16'd9397;
      89547:data<=16'd8493;
      89548:data<=16'd7787;
      89549:data<=16'd7407;
      89550:data<=16'd6269;
      89551:data<=16'd5192;
      89552:data<=16'd4472;
      89553:data<=16'd4360;
      89554:data<=16'd4309;
      89555:data<=16'd4874;
      89556:data<=16'd5900;
      89557:data<=16'd5906;
      89558:data<=16'd5779;
      89559:data<=16'd4784;
      89560:data<=16'd3924;
      89561:data<=16'd5092;
      89562:data<=16'd4626;
      89563:data<=16'd4293;
      89564:data<=16'd2344;
      89565:data<=-16'd10859;
      89566:data<=-16'd24242;
      89567:data<=-16'd24682;
      89568:data<=-16'd22542;
      89569:data<=-16'd22259;
      89570:data<=-16'd20315;
      89571:data<=-16'd20186;
      89572:data<=-16'd20359;
      89573:data<=-16'd18475;
      89574:data<=-16'd17007;
      89575:data<=-16'd16084;
      89576:data<=-16'd15479;
      89577:data<=-16'd15247;
      89578:data<=-16'd15374;
      89579:data<=-16'd15286;
      89580:data<=-16'd13594;
      89581:data<=-16'd12551;
      89582:data<=-16'd12602;
      89583:data<=-16'd11083;
      89584:data<=-16'd9888;
      89585:data<=-16'd9812;
      89586:data<=-16'd8772;
      89587:data<=-16'd7724;
      89588:data<=-16'd7330;
      89589:data<=-16'd7010;
      89590:data<=-16'd7272;
      89591:data<=-16'd7894;
      89592:data<=-16'd7201;
      89593:data<=-16'd5554;
      89594:data<=-16'd5964;
      89595:data<=-16'd7060;
      89596:data<=-16'd5844;
      89597:data<=-16'd4511;
      89598:data<=-16'd3987;
      89599:data<=-16'd3903;
      89600:data<=-16'd4573;
      89601:data<=-16'd3788;
      89602:data<=-16'd2757;
      89603:data<=-16'd2828;
      89604:data<=-16'd2863;
      89605:data<=-16'd4573;
      89606:data<=-16'd3899;
      89607:data<=-16'd790;
      89608:data<=-16'd3119;
      89609:data<=-16'd429;
      89610:data<=16'd12580;
      89611:data<=16'd17593;
      89612:data<=16'd15603;
      89613:data<=16'd17279;
      89614:data<=16'd16334;
      89615:data<=16'd14885;
      89616:data<=16'd15746;
      89617:data<=16'd13153;
      89618:data<=16'd14041;
      89619:data<=16'd20192;
      89620:data<=16'd21422;
      89621:data<=16'd19553;
      89622:data<=16'd19050;
      89623:data<=16'd18387;
      89624:data<=16'd17973;
      89625:data<=16'd17114;
      89626:data<=16'd15803;
      89627:data<=16'd15133;
      89628:data<=16'd14522;
      89629:data<=16'd14592;
      89630:data<=16'd13687;
      89631:data<=16'd11122;
      89632:data<=16'd10922;
      89633:data<=16'd11950;
      89634:data<=16'd11599;
      89635:data<=16'd11906;
      89636:data<=16'd11668;
      89637:data<=16'd9691;
      89638:data<=16'd8854;
      89639:data<=16'd9451;
      89640:data<=16'd9861;
      89641:data<=16'd9482;
      89642:data<=16'd8378;
      89643:data<=16'd8102;
      89644:data<=16'd9016;
      89645:data<=16'd8710;
      89646:data<=16'd7394;
      89647:data<=16'd7864;
      89648:data<=16'd8181;
      89649:data<=16'd6711;
      89650:data<=16'd6925;
      89651:data<=16'd7400;
      89652:data<=16'd7009;
      89653:data<=16'd7850;
      89654:data<=16'd1715;
      89655:data<=-16'd10853;
      89656:data<=-16'd13808;
      89657:data<=-16'd9888;
      89658:data<=-16'd9459;
      89659:data<=-16'd8470;
      89660:data<=-16'd7083;
      89661:data<=-16'd7245;
      89662:data<=-16'd6822;
      89663:data<=-16'd7451;
      89664:data<=-16'd7068;
      89665:data<=-16'd5752;
      89666:data<=-16'd6367;
      89667:data<=-16'd4868;
      89668:data<=-16'd3636;
      89669:data<=-16'd4772;
      89670:data<=-16'd2513;
      89671:data<=-16'd2221;
      89672:data<=-16'd6692;
      89673:data<=-16'd7717;
      89674:data<=-16'd7060;
      89675:data<=-16'd7562;
      89676:data<=-16'd6704;
      89677:data<=-16'd6310;
      89678:data<=-16'd6217;
      89679:data<=-16'd5532;
      89680:data<=-16'd5090;
      89681:data<=-16'd4190;
      89682:data<=-16'd4770;
      89683:data<=-16'd5418;
      89684:data<=-16'd2649;
      89685:data<=-16'd902;
      89686:data<=-16'd1230;
      89687:data<=16'd138;
      89688:data<=16'd509;
      89689:data<=-16'd466;
      89690:data<=16'd281;
      89691:data<=16'd237;
      89692:data<=-16'd326;
      89693:data<=16'd1199;
      89694:data<=16'd1325;
      89695:data<=16'd581;
      89696:data<=16'd1695;
      89697:data<=16'd1287;
      89698:data<=16'd4485;
      89699:data<=16'd15782;
      89700:data<=16'd21996;
      89701:data<=16'd19890;
      89702:data<=16'd19644;
      89703:data<=16'd19340;
      89704:data<=16'd17447;
      89705:data<=16'd17509;
      89706:data<=16'd16913;
      89707:data<=16'd16516;
      89708:data<=16'd17067;
      89709:data<=16'd16340;
      89710:data<=16'd17250;
      89711:data<=16'd17951;
      89712:data<=16'd15922;
      89713:data<=16'd15693;
      89714:data<=16'd15524;
      89715:data<=16'd13305;
      89716:data<=16'd12925;
      89717:data<=16'd12966;
      89718:data<=16'd11819;
      89719:data<=16'd11323;
      89720:data<=16'd10786;
      89721:data<=16'd10586;
      89722:data<=16'd10898;
      89723:data<=16'd10457;
      89724:data<=16'd12149;
      89725:data<=16'd17029;
      89726:data<=16'd20162;
      89727:data<=16'd20113;
      89728:data<=16'd19229;
      89729:data<=16'd17943;
      89730:data<=16'd17440;
      89731:data<=16'd17274;
      89732:data<=16'd15496;
      89733:data<=16'd14939;
      89734:data<=16'd15041;
      89735:data<=16'd13324;
      89736:data<=16'd14395;
      89737:data<=16'd15800;
      89738:data<=16'd13256;
      89739:data<=16'd12734;
      89740:data<=16'd12468;
      89741:data<=16'd11103;
      89742:data<=16'd13285;
      89743:data<=16'd8226;
      89744:data<=-16'd4863;
      89745:data<=-16'd8581;
      89746:data<=-16'd6398;
      89747:data<=-16'd7485;
      89748:data<=-16'd7163;
      89749:data<=-16'd6385;
      89750:data<=-16'd6068;
      89751:data<=-16'd3943;
      89752:data<=-16'd3463;
      89753:data<=-16'd4413;
      89754:data<=-16'd4475;
      89755:data<=-16'd4746;
      89756:data<=-16'd4628;
      89757:data<=-16'd4014;
      89758:data<=-16'd4017;
      89759:data<=-16'd4032;
      89760:data<=-16'd3239;
      89761:data<=-16'd2826;
      89762:data<=-16'd3811;
      89763:data<=-16'd3127;
      89764:data<=-16'd481;
      89765:data<=-16'd158;
      89766:data<=-16'd829;
      89767:data<=-16'd497;
      89768:data<=-16'd1384;
      89769:data<=-16'd1971;
      89770:data<=-16'd719;
      89771:data<=-16'd716;
      89772:data<=-16'd2199;
      89773:data<=-16'd1844;
      89774:data<=-16'd914;
      89775:data<=-16'd1920;
      89776:data<=-16'd984;
      89777:data<=16'd808;
      89778:data<=-16'd2949;
      89779:data<=-16'd7307;
      89780:data<=-16'd7482;
      89781:data<=-16'd7551;
      89782:data<=-16'd7573;
      89783:data<=-16'd7362;
      89784:data<=-16'd6965;
      89785:data<=-16'd5836;
      89786:data<=-16'd7715;
      89787:data<=-16'd5970;
      89788:data<=16'd5380;
      89789:data<=16'd13235;
      89790:data<=16'd13242;
      89791:data<=16'd13262;
      89792:data<=16'd12906;
      89793:data<=16'd12413;
      89794:data<=16'd12516;
      89795:data<=16'd11097;
      89796:data<=16'd10081;
      89797:data<=16'd9873;
      89798:data<=16'd9950;
      89799:data<=16'd10202;
      89800:data<=16'd8439;
      89801:data<=16'd6937;
      89802:data<=16'd7673;
      89803:data<=16'd8158;
      89804:data<=16'd7783;
      89805:data<=16'd6579;
      89806:data<=16'd5782;
      89807:data<=16'd6064;
      89808:data<=16'd5292;
      89809:data<=16'd4704;
      89810:data<=16'd5134;
      89811:data<=16'd5065;
      89812:data<=16'd5150;
      89813:data<=16'd4602;
      89814:data<=16'd3271;
      89815:data<=16'd3011;
      89816:data<=16'd4243;
      89817:data<=16'd6185;
      89818:data<=16'd5548;
      89819:data<=16'd3664;
      89820:data<=16'd4746;
      89821:data<=16'd4802;
      89822:data<=16'd3271;
      89823:data<=16'd2772;
      89824:data<=16'd1055;
      89825:data<=16'd1706;
      89826:data<=16'd3054;
      89827:data<=-16'd39;
      89828:data<=16'd238;
      89829:data<=16'd1562;
      89830:data<=-16'd82;
      89831:data<=16'd5680;
      89832:data<=16'd7843;
      89833:data<=-16'd4252;
      89834:data<=-16'd10710;
      89835:data<=-16'd7978;
      89836:data<=-16'd7991;
      89837:data<=-16'd7529;
      89838:data<=-16'd7121;
      89839:data<=-16'd8745;
      89840:data<=-16'd7750;
      89841:data<=-16'd6470;
      89842:data<=-16'd6237;
      89843:data<=-16'd5024;
      89844:data<=-16'd4510;
      89845:data<=-16'd4391;
      89846:data<=-16'd4285;
      89847:data<=-16'd4505;
      89848:data<=-16'd3990;
      89849:data<=-16'd3680;
      89850:data<=-16'd3724;
      89851:data<=-16'd4159;
      89852:data<=-16'd5306;
      89853:data<=-16'd4689;
      89854:data<=-16'd3635;
      89855:data<=-16'd4642;
      89856:data<=-16'd4896;
      89857:data<=-16'd4297;
      89858:data<=-16'd4701;
      89859:data<=-16'd4378;
      89860:data<=-16'd3545;
      89861:data<=-16'd4338;
      89862:data<=-16'd5245;
      89863:data<=-16'd4241;
      89864:data<=-16'd3485;
      89865:data<=-16'd3936;
      89866:data<=-16'd3641;
      89867:data<=-16'd3706;
      89868:data<=-16'd4150;
      89869:data<=-16'd4256;
      89870:data<=-16'd6369;
      89871:data<=-16'd7181;
      89872:data<=-16'd5513;
      89873:data<=-16'd6308;
      89874:data<=-16'd6375;
      89875:data<=-16'd6038;
      89876:data<=-16'd6740;
      89877:data<=16'd1921;
      89878:data<=16'd13233;
      89879:data<=16'd13115;
      89880:data<=16'd11244;
      89881:data<=16'd11919;
      89882:data<=16'd10044;
      89883:data<=16'd9417;
      89884:data<=16'd6222;
      89885:data<=-16'd1037;
      89886:data<=-16'd3451;
      89887:data<=-16'd2598;
      89888:data<=-16'd2699;
      89889:data<=-16'd2652;
      89890:data<=-16'd2813;
      89891:data<=-16'd2611;
      89892:data<=-16'd3221;
      89893:data<=-16'd4393;
      89894:data<=-16'd3536;
      89895:data<=-16'd3680;
      89896:data<=-16'd5203;
      89897:data<=-16'd5153;
      89898:data<=-16'd5565;
      89899:data<=-16'd6686;
      89900:data<=-16'd6731;
      89901:data<=-16'd6240;
      89902:data<=-16'd5843;
      89903:data<=-16'd6115;
      89904:data<=-16'd6223;
      89905:data<=-16'd5691;
      89906:data<=-16'd5642;
      89907:data<=-16'd5412;
      89908:data<=-16'd4884;
      89909:data<=-16'd5315;
      89910:data<=-16'd6507;
      89911:data<=-16'd7115;
      89912:data<=-16'd7233;
      89913:data<=-16'd8296;
      89914:data<=-16'd7982;
      89915:data<=-16'd5956;
      89916:data<=-16'd6482;
      89917:data<=-16'd6972;
      89918:data<=-16'd6543;
      89919:data<=-16'd7608;
      89920:data<=-16'd5512;
      89921:data<=-16'd7262;
      89922:data<=-16'd19591;
      89923:data<=-16'd26156;
      89924:data<=-16'd23595;
      89925:data<=-16'd23376;
      89926:data<=-16'd22483;
      89927:data<=-16'd20553;
      89928:data<=-16'd20480;
      89929:data<=-16'd18958;
      89930:data<=-16'd18472;
      89931:data<=-16'd18456;
      89932:data<=-16'd16654;
      89933:data<=-16'd16701;
      89934:data<=-16'd15978;
      89935:data<=-16'd15048;
      89936:data<=-16'd17702;
      89937:data<=-16'd15793;
      89938:data<=-16'd8434;
      89939:data<=-16'd5777;
      89940:data<=-16'd6552;
      89941:data<=-16'd5330;
      89942:data<=-16'd4451;
      89943:data<=-16'd5385;
      89944:data<=-16'd5865;
      89945:data<=-16'd5327;
      89946:data<=-16'd4584;
      89947:data<=-16'd4150;
      89948:data<=-16'd4958;
      89949:data<=-16'd6023;
      89950:data<=-16'd6369;
      89951:data<=-16'd6830;
      89952:data<=-16'd6120;
      89953:data<=-16'd5204;
      89954:data<=-16'd5480;
      89955:data<=-16'd4303;
      89956:data<=-16'd4021;
      89957:data<=-16'd5113;
      89958:data<=-16'd3876;
      89959:data<=-16'd4185;
      89960:data<=-16'd4467;
      89961:data<=-16'd2188;
      89962:data<=-16'd4099;
      89963:data<=-16'd5115;
      89964:data<=-16'd3462;
      89965:data<=-16'd6399;
      89966:data<=-16'd1177;
      89967:data<=16'd12624;
      89968:data<=16'd14719;
      89969:data<=16'd11094;
      89970:data<=16'd12198;
      89971:data<=16'd11665;
      89972:data<=16'd10871;
      89973:data<=16'd11089;
      89974:data<=16'd10099;
      89975:data<=16'd9835;
      89976:data<=16'd8449;
      89977:data<=16'd6937;
      89978:data<=16'd7297;
      89979:data<=16'd6314;
      89980:data<=16'd5877;
      89981:data<=16'd6566;
      89982:data<=16'd5137;
      89983:data<=16'd4288;
      89984:data<=16'd4899;
      89985:data<=16'd5078;
      89986:data<=16'd5520;
      89987:data<=16'd4995;
      89988:data<=16'd4073;
      89989:data<=16'd4358;
      89990:data<=16'd1695;
      89991:data<=-16'd4205;
      89992:data<=-16'd6651;
      89993:data<=-16'd5482;
      89994:data<=-16'd5277;
      89995:data<=-16'd5597;
      89996:data<=-16'd5750;
      89997:data<=-16'd5994;
      89998:data<=-16'd4558;
      89999:data<=-16'd2917;
      90000:data<=-16'd2887;
      90001:data<=-16'd3594;
      90002:data<=-16'd5247;
      90003:data<=-16'd5517;
      90004:data<=-16'd4053;
      90005:data<=-16'd4238;
      90006:data<=-16'd3883;
      90007:data<=-16'd3610;
      90008:data<=-16'd4921;
      90009:data<=-16'd2977;
      90010:data<=-16'd4875;
      90011:data<=-16'd15769;
      90012:data<=-16'd21086;
      90013:data<=-16'd18618;
      90014:data<=-16'd18069;
      90015:data<=-16'd17750;
      90016:data<=-16'd17575;
      90017:data<=-16'd18407;
      90018:data<=-16'd16713;
      90019:data<=-16'd15346;
      90020:data<=-16'd15403;
      90021:data<=-16'd14314;
      90022:data<=-16'd13624;
      90023:data<=-16'd12743;
      90024:data<=-16'd11354;
      90025:data<=-16'd11294;
      90026:data<=-16'd10461;
      90027:data<=-16'd8992;
      90028:data<=-16'd9639;
      90029:data<=-16'd10351;
      90030:data<=-16'd9388;
      90031:data<=-16'd8683;
      90032:data<=-16'd8319;
      90033:data<=-16'd7341;
      90034:data<=-16'd6928;
      90035:data<=-16'd7078;
      90036:data<=-16'd6846;
      90037:data<=-16'd6710;
      90038:data<=-16'd5962;
      90039:data<=-16'd5083;
      90040:data<=-16'd5145;
      90041:data<=-16'd4484;
      90042:data<=-16'd4792;
      90043:data<=-16'd4872;
      90044:data<=16'd649;
      90045:data<=16'd5018;
      90046:data<=16'd4044;
      90047:data<=16'd5238;
      90048:data<=16'd6137;
      90049:data<=16'd4617;
      90050:data<=16'd5077;
      90051:data<=16'd4558;
      90052:data<=16'd5271;
      90053:data<=16'd7250;
      90054:data<=16'd3915;
      90055:data<=16'd6596;
      90056:data<=16'd18726;
      90057:data<=16'd22870;
      90058:data<=16'd20154;
      90059:data<=16'd19408;
      90060:data<=16'd18337;
      90061:data<=16'd18456;
      90062:data<=16'd18653;
      90063:data<=16'd17054;
      90064:data<=16'd17217;
      90065:data<=16'd16879;
      90066:data<=16'd15893;
      90067:data<=16'd16468;
      90068:data<=16'd14963;
      90069:data<=16'd13540;
      90070:data<=16'd14894;
      90071:data<=16'd14747;
      90072:data<=16'd13204;
      90073:data<=16'd12637;
      90074:data<=16'd12709;
      90075:data<=16'd12636;
      90076:data<=16'd11665;
      90077:data<=16'd11336;
      90078:data<=16'd11765;
      90079:data<=16'd10968;
      90080:data<=16'd10281;
      90081:data<=16'd10877;
      90082:data<=16'd11693;
      90083:data<=16'd11943;
      90084:data<=16'd11635;
      90085:data<=16'd11247;
      90086:data<=16'd10223;
      90087:data<=16'd9368;
      90088:data<=16'd9529;
      90089:data<=16'd8912;
      90090:data<=16'd8495;
      90091:data<=16'd8769;
      90092:data<=16'd8028;
      90093:data<=16'd7677;
      90094:data<=16'd7780;
      90095:data<=16'd9054;
      90096:data<=16'd10345;
      90097:data<=16'd5207;
      90098:data<=-16'd174;
      90099:data<=-16'd734;
      90100:data<=-16'd8319;
      90101:data<=-16'd18378;
      90102:data<=-16'd18099;
      90103:data<=-16'd15386;
      90104:data<=-16'd14933;
      90105:data<=-16'd13649;
      90106:data<=-16'd13585;
      90107:data<=-16'd12900;
      90108:data<=-16'd11057;
      90109:data<=-16'd10154;
      90110:data<=-16'd9154;
      90111:data<=-16'd9297;
      90112:data<=-16'd9696;
      90113:data<=-16'd8889;
      90114:data<=-16'd8643;
      90115:data<=-16'd7614;
      90116:data<=-16'd6772;
      90117:data<=-16'd7131;
      90118:data<=-16'd5560;
      90119:data<=-16'd4701;
      90120:data<=-16'd5557;
      90121:data<=-16'd4135;
      90122:data<=-16'd2496;
      90123:data<=-16'd2382;
      90124:data<=-16'd2229;
      90125:data<=-16'd2209;
      90126:data<=-16'd1980;
      90127:data<=-16'd1709;
      90128:data<=-16'd1430;
      90129:data<=-16'd588;
      90130:data<=-16'd117;
      90131:data<=-16'd287;
      90132:data<=-16'd852;
      90133:data<=-16'd675;
      90134:data<=16'd766;
      90135:data<=16'd1791;
      90136:data<=16'd2631;
      90137:data<=16'd2626;
      90138:data<=16'd1765;
      90139:data<=16'd2093;
      90140:data<=16'd1322;
      90141:data<=16'd1563;
      90142:data<=16'd3266;
      90143:data<=16'd461;
      90144:data<=16'd4328;
      90145:data<=16'd17728;
      90146:data<=16'd20433;
      90147:data<=16'd17239;
      90148:data<=16'd19108;
      90149:data<=16'd17394;
      90150:data<=16'd18859;
      90151:data<=16'd25737;
      90152:data<=16'd24980;
      90153:data<=16'd22563;
      90154:data<=16'd23334;
      90155:data<=16'd22008;
      90156:data<=16'd21346;
      90157:data<=16'd20541;
      90158:data<=16'd18958;
      90159:data<=16'd18859;
      90160:data<=16'd17478;
      90161:data<=16'd17144;
      90162:data<=16'd18589;
      90163:data<=16'd17643;
      90164:data<=16'd16644;
      90165:data<=16'd16404;
      90166:data<=16'd15559;
      90167:data<=16'd15432;
      90168:data<=16'd15154;
      90169:data<=16'd14260;
      90170:data<=16'd12986;
      90171:data<=16'd12193;
      90172:data<=16'd12657;
      90173:data<=16'd11770;
      90174:data<=16'd10636;
      90175:data<=16'd11259;
      90176:data<=16'd11297;
      90177:data<=16'd10862;
      90178:data<=16'd10229;
      90179:data<=16'd9747;
      90180:data<=16'd9817;
      90181:data<=16'd8537;
      90182:data<=16'd8249;
      90183:data<=16'd8313;
      90184:data<=16'd6899;
      90185:data<=16'd8202;
      90186:data<=16'd7492;
      90187:data<=16'd5333;
      90188:data<=16'd8748;
      90189:data<=16'd3808;
      90190:data<=-16'd9423;
      90191:data<=-16'd11191;
      90192:data<=-16'd8536;
      90193:data<=-16'd9823;
      90194:data<=-16'd8774;
      90195:data<=-16'd8492;
      90196:data<=-16'd8567;
      90197:data<=-16'd7802;
      90198:data<=-16'd9027;
      90199:data<=-16'd8166;
      90200:data<=-16'd7750;
      90201:data<=-16'd8410;
      90202:data<=-16'd5241;
      90203:data<=-16'd6871;
      90204:data<=-16'd13650;
      90205:data<=-16'd14675;
      90206:data<=-16'd12966;
      90207:data<=-16'd12660;
      90208:data<=-16'd12471;
      90209:data<=-16'd12812;
      90210:data<=-16'd12225;
      90211:data<=-16'd11191;
      90212:data<=-16'd10665;
      90213:data<=-16'd10202;
      90214:data<=-16'd10155;
      90215:data<=-16'd8883;
      90216:data<=-16'd7746;
      90217:data<=-16'd8366;
      90218:data<=-16'd7827;
      90219:data<=-16'd6996;
      90220:data<=-16'd6946;
      90221:data<=-16'd6425;
      90222:data<=-16'd6757;
      90223:data<=-16'd6989;
      90224:data<=-16'd5896;
      90225:data<=-16'd5288;
      90226:data<=-16'd5485;
      90227:data<=-16'd4793;
      90228:data<=-16'd2904;
      90229:data<=-16'd2940;
      90230:data<=-16'd3704;
      90231:data<=-16'd2820;
      90232:data<=-16'd4570;
      90233:data<=-16'd2328;
      90234:data<=16'd9535;
      90235:data<=16'd15247;
      90236:data<=16'd12483;
      90237:data<=16'd12751;
      90238:data<=16'd12542;
      90239:data<=16'd11268;
      90240:data<=16'd11564;
      90241:data<=16'd10399;
      90242:data<=16'd10889;
      90243:data<=16'd11573;
      90244:data<=16'd9944;
      90245:data<=16'd10525;
      90246:data<=16'd10149;
      90247:data<=16'd8335;
      90248:data<=16'd8995;
      90249:data<=16'd8316;
      90250:data<=16'd7715;
      90251:data<=16'd8291;
      90252:data<=16'd6020;
      90253:data<=16'd5504;
      90254:data<=16'd6930;
      90255:data<=16'd5583;
      90256:data<=16'd7262;
      90257:data<=16'd13035;
      90258:data<=16'd14848;
      90259:data<=16'd13141;
      90260:data<=16'd13098;
      90261:data<=16'd13285;
      90262:data<=16'd12046;
      90263:data<=16'd11402;
      90264:data<=16'd10182;
      90265:data<=16'd8387;
      90266:data<=16'd8658;
      90267:data<=16'd9060;
      90268:data<=16'd9597;
      90269:data<=16'd10464;
      90270:data<=16'd8900;
      90271:data<=16'd8552;
      90272:data<=16'd8933;
      90273:data<=16'd7080;
      90274:data<=16'd7947;
      90275:data<=16'd7397;
      90276:data<=16'd4652;
      90277:data<=16'd7269;
      90278:data<=16'd2921;
      90279:data<=-16'd10554;
      90280:data<=-16'd13985;
      90281:data<=-16'd11453;
      90282:data<=-16'd12088;
      90283:data<=-16'd10831;
      90284:data<=-16'd10759;
      90285:data<=-16'd11814;
      90286:data<=-16'd9976;
      90287:data<=-16'd9588;
      90288:data<=-16'd10103;
      90289:data<=-16'd9802;
      90290:data<=-16'd10608;
      90291:data<=-16'd10210;
      90292:data<=-16'd8978;
      90293:data<=-16'd9398;
      90294:data<=-16'd10188;
      90295:data<=-16'd10320;
      90296:data<=-16'd9788;
      90297:data<=-16'd9799;
      90298:data<=-16'd10281;
      90299:data<=-16'd9236;
      90300:data<=-16'd8343;
      90301:data<=-16'd8857;
      90302:data<=-16'd9172;
      90303:data<=-16'd9721;
      90304:data<=-16'd10013;
      90305:data<=-16'd9074;
      90306:data<=-16'd9098;
      90307:data<=-16'd9800;
      90308:data<=-16'd8969;
      90309:data<=-16'd10078;
      90310:data<=-16'd15059;
      90311:data<=-16'd17525;
      90312:data<=-16'd16145;
      90313:data<=-16'd16019;
      90314:data<=-16'd15803;
      90315:data<=-16'd14475;
      90316:data<=-16'd14424;
      90317:data<=-16'd13963;
      90318:data<=-16'd13342;
      90319:data<=-16'd13133;
      90320:data<=-16'd12542;
      90321:data<=-16'd14580;
      90322:data<=-16'd13367;
      90323:data<=-16'd2708;
      90324:data<=16'd5031;
      90325:data<=16'd3971;
      90326:data<=16'd2839;
      90327:data<=16'd2704;
      90328:data<=16'd2608;
      90329:data<=16'd3287;
      90330:data<=16'd2497;
      90331:data<=16'd2467;
      90332:data<=16'd3262;
      90333:data<=16'd1560;
      90334:data<=16'd526;
      90335:data<=16'd675;
      90336:data<=-16'd851;
      90337:data<=-16'd1454;
      90338:data<=-16'd558;
      90339:data<=-16'd384;
      90340:data<=-16'd435;
      90341:data<=-16'd499;
      90342:data<=-16'd487;
      90343:data<=-16'd629;
      90344:data<=-16'd1712;
      90345:data<=-16'd1965;
      90346:data<=-16'd1240;
      90347:data<=-16'd1973;
      90348:data<=-16'd2999;
      90349:data<=-16'd2710;
      90350:data<=-16'd2684;
      90351:data<=-16'd3251;
      90352:data<=-16'd3419;
      90353:data<=-16'd3022;
      90354:data<=-16'd2109;
      90355:data<=-16'd1968;
      90356:data<=-16'd2754;
      90357:data<=-16'd2322;
      90358:data<=-16'd1670;
      90359:data<=-16'd1906;
      90360:data<=-16'd1989;
      90361:data<=-16'd3932;
      90362:data<=-16'd4096;
      90363:data<=16'd2347;
      90364:data<=16'd5338;
      90365:data<=16'd3078;
      90366:data<=16'd5535;
      90367:data<=16'd2525;
      90368:data<=-16'd10519;
      90369:data<=-16'd15130;
      90370:data<=-16'd12075;
      90371:data<=-16'd12689;
      90372:data<=-16'd12516;
      90373:data<=-16'd11828;
      90374:data<=-16'd13135;
      90375:data<=-16'd12377;
      90376:data<=-16'd11582;
      90377:data<=-16'd11655;
      90378:data<=-16'd10539;
      90379:data<=-16'd10258;
      90380:data<=-16'd9700;
      90381:data<=-16'd7962;
      90382:data<=-16'd7670;
      90383:data<=-16'd8270;
      90384:data<=-16'd8182;
      90385:data<=-16'd7421;
      90386:data<=-16'd7439;
      90387:data<=-16'd8812;
      90388:data<=-16'd9125;
      90389:data<=-16'd8558;
      90390:data<=-16'd8416;
      90391:data<=-16'd7712;
      90392:data<=-16'd7062;
      90393:data<=-16'd6554;
      90394:data<=-16'd5908;
      90395:data<=-16'd6202;
      90396:data<=-16'd6044;
      90397:data<=-16'd4608;
      90398:data<=-16'd3858;
      90399:data<=-16'd4913;
      90400:data<=-16'd6269;
      90401:data<=-16'd5676;
      90402:data<=-16'd5124;
      90403:data<=-16'd5876;
      90404:data<=-16'd5473;
      90405:data<=-16'd5031;
      90406:data<=-16'd4761;
      90407:data<=-16'd4170;
      90408:data<=-16'd4827;
      90409:data<=-16'd3751;
      90410:data<=-16'd3380;
      90411:data<=-16'd4922;
      90412:data<=16'd2695;
      90413:data<=16'd13083;
      90414:data<=16'd12750;
      90415:data<=16'd10288;
      90416:data<=16'd7950;
      90417:data<=16'd2267;
      90418:data<=16'd1254;
      90419:data<=16'd2215;
      90420:data<=16'd957;
      90421:data<=16'd2347;
      90422:data<=16'd3010;
      90423:data<=16'd1695;
      90424:data<=16'd2226;
      90425:data<=16'd2431;
      90426:data<=16'd1554;
      90427:data<=16'd528;
      90428:data<=-16'd20;
      90429:data<=16'd379;
      90430:data<=-16'd185;
      90431:data<=-16'd214;
      90432:data<=16'd661;
      90433:data<=-16'd123;
      90434:data<=-16'd135;
      90435:data<=16'd623;
      90436:data<=16'd194;
      90437:data<=16'd723;
      90438:data<=16'd1089;
      90439:data<=16'd18;
      90440:data<=-16'd758;
      90441:data<=-16'd1472;
      90442:data<=-16'd1856;
      90443:data<=-16'd1475;
      90444:data<=-16'd1068;
      90445:data<=-16'd1010;
      90446:data<=-16'd1538;
      90447:data<=-16'd1729;
      90448:data<=-16'd989;
      90449:data<=16'd105;
      90450:data<=16'd194;
      90451:data<=-16'd508;
      90452:data<=16'd722;
      90453:data<=16'd331;
      90454:data<=-16'd2566;
      90455:data<=-16'd863;
      90456:data<=-16'd2861;
      90457:data<=-16'd14390;
      90458:data<=-16'd19287;
      90459:data<=-16'd16352;
      90460:data<=-16'd15784;
      90461:data<=-16'd14965;
      90462:data<=-16'd14446;
      90463:data<=-16'd14025;
      90464:data<=-16'd11536;
      90465:data<=-16'd11805;
      90466:data<=-16'd11914;
      90467:data<=-16'd10921;
      90468:data<=-16'd12972;
      90469:data<=-16'd9846;
      90470:data<=-16'd2252;
      90471:data<=-16'd1121;
      90472:data<=-16'd2264;
      90473:data<=-16'd1190;
      90474:data<=-16'd1381;
      90475:data<=-16'd1592;
      90476:data<=-16'd431;
      90477:data<=16'd375;
      90478:data<=16'd447;
      90479:data<=16'd277;
      90480:data<=-16'd678;
      90481:data<=-16'd1619;
      90482:data<=-16'd696;
      90483:data<=-16'd140;
      90484:data<=-16'd628;
      90485:data<=16'd44;
      90486:data<=16'd27;
      90487:data<=16'd71;
      90488:data<=16'd1078;
      90489:data<=16'd321;
      90490:data<=16'd666;
      90491:data<=16'd2074;
      90492:data<=16'd1488;
      90493:data<=16'd1856;
      90494:data<=16'd1862;
      90495:data<=16'd1256;
      90496:data<=16'd2417;
      90497:data<=16'd1569;
      90498:data<=16'd1915;
      90499:data<=16'd3583;
      90500:data<=16'd758;
      90501:data<=16'd5374;
      90502:data<=16'd18389;
      90503:data<=16'd21359;
      90504:data<=16'd18399;
      90505:data<=16'd19174;
      90506:data<=16'd18991;
      90507:data<=16'd18974;
      90508:data<=16'd19229;
      90509:data<=16'd17264;
      90510:data<=16'd16819;
      90511:data<=16'd17071;
      90512:data<=16'd16031;
      90513:data<=16'd15452;
      90514:data<=16'd14703;
      90515:data<=16'd14192;
      90516:data<=16'd14305;
      90517:data<=16'd13929;
      90518:data<=16'd13708;
      90519:data<=16'd13170;
      90520:data<=16'd12942;
      90521:data<=16'd13826;
      90522:data<=16'd11176;
      90523:data<=16'd4886;
      90524:data<=16'd2126;
      90525:data<=16'd3113;
      90526:data<=16'd3180;
      90527:data<=16'd2816;
      90528:data<=16'd2978;
      90529:data<=16'd3048;
      90530:data<=16'd3419;
      90531:data<=16'd2836;
      90532:data<=16'd2237;
      90533:data<=16'd4322;
      90534:data<=16'd5347;
      90535:data<=16'd3607;
      90536:data<=16'd3383;
      90537:data<=16'd4020;
      90538:data<=16'd3920;
      90539:data<=16'd3764;
      90540:data<=16'd3078;
      90541:data<=16'd3562;
      90542:data<=16'd3688;
      90543:data<=16'd2291;
      90544:data<=16'd3996;
      90545:data<=16'd2487;
      90546:data<=-16'd7454;
      90547:data<=-16'd12739;
      90548:data<=-16'd10784;
      90549:data<=-16'd10903;
      90550:data<=-16'd11176;
      90551:data<=-16'd10583;
      90552:data<=-16'd10807;
      90553:data<=-16'd9109;
      90554:data<=-16'd8273;
      90555:data<=-16'd9360;
      90556:data<=-16'd8692;
      90557:data<=-16'd8281;
      90558:data<=-16'd8025;
      90559:data<=-16'd5547;
      90560:data<=-16'd3958;
      90561:data<=-16'd4181;
      90562:data<=-16'd4296;
      90563:data<=-16'd4121;
      90564:data<=-16'd3360;
      90565:data<=-16'd2681;
      90566:data<=-16'd2429;
      90567:data<=-16'd1979;
      90568:data<=-16'd1804;
      90569:data<=-16'd1195;
      90570:data<=-16'd717;
      90571:data<=-16'd1859;
      90572:data<=-16'd1249;
      90573:data<=16'd1172;
      90574:data<=16'd883;
      90575:data<=16'd2255;
      90576:data<=16'd8243;
      90577:data<=16'd10046;
      90578:data<=16'd7703;
      90579:data<=16'd8962;
      90580:data<=16'd9743;
      90581:data<=16'd7642;
      90582:data<=16'd7588;
      90583:data<=16'd7304;
      90584:data<=16'd6466;
      90585:data<=16'd7548;
      90586:data<=16'd7462;
      90587:data<=16'd8654;
      90588:data<=16'd10255;
      90589:data<=16'd6962;
      90590:data<=16'd10328;
      90591:data<=16'd22532;
      90592:data<=16'd25611;
      90593:data<=16'd22024;
      90594:data<=16'd22341;
      90595:data<=16'd21570;
      90596:data<=16'd20116;
      90597:data<=16'd19852;
      90598:data<=16'd18057;
      90599:data<=16'd18682;
      90600:data<=16'd20260;
      90601:data<=16'd18407;
      90602:data<=16'd17719;
      90603:data<=16'd17976;
      90604:data<=16'd15872;
      90605:data<=16'd14736;
      90606:data<=16'd14900;
      90607:data<=16'd14220;
      90608:data<=16'd13870;
      90609:data<=16'd13239;
      90610:data<=16'd11198;
      90611:data<=16'd10114;
      90612:data<=16'd11077;
      90613:data<=16'd11887;
      90614:data<=16'd11673;
      90615:data<=16'd11041;
      90616:data<=16'd10138;
      90617:data<=16'd9497;
      90618:data<=16'd9097;
      90619:data<=16'd8678;
      90620:data<=16'd7908;
      90621:data<=16'd6184;
      90622:data<=16'd5658;
      90623:data<=16'd6536;
      90624:data<=16'd5498;
      90625:data<=16'd4625;
      90626:data<=16'd6523;
      90627:data<=16'd7885;
      90628:data<=16'd5398;
      90629:data<=-16'd506;
      90630:data<=-16'd3862;
      90631:data<=-16'd3045;
      90632:data<=-16'd4244;
      90633:data<=-16'd4767;
      90634:data<=-16'd4187;
      90635:data<=-16'd11950;
      90636:data<=-16'd20926;
      90637:data<=-16'd20770;
      90638:data<=-16'd18836;
      90639:data<=-16'd18171;
      90640:data<=-16'd16622;
      90641:data<=-16'd16242;
      90642:data<=-16'd15587;
      90643:data<=-16'd15076;
      90644:data<=-16'd15676;
      90645:data<=-16'd14499;
      90646:data<=-16'd13355;
      90647:data<=-16'd13770;
      90648:data<=-16'd13355;
      90649:data<=-16'd12519;
      90650:data<=-16'd12135;
      90651:data<=-16'd11975;
      90652:data<=-16'd11127;
      90653:data<=-16'd9042;
      90654:data<=-16'd8052;
      90655:data<=-16'd8270;
      90656:data<=-16'd7688;
      90657:data<=-16'd6987;
      90658:data<=-16'd6546;
      90659:data<=-16'd6440;
      90660:data<=-16'd7330;
      90661:data<=-16'd7814;
      90662:data<=-16'd6898;
      90663:data<=-16'd6229;
      90664:data<=-16'd6536;
      90665:data<=-16'd5780;
      90666:data<=-16'd4062;
      90667:data<=-16'd3557;
      90668:data<=-16'd3096;
      90669:data<=-16'd2485;
      90670:data<=-16'd3001;
      90671:data<=-16'd2887;
      90672:data<=-16'd2679;
      90673:data<=-16'd3052;
      90674:data<=-16'd2713;
      90675:data<=-16'd2535;
      90676:data<=-16'd1115;
      90677:data<=-16'd867;
      90678:data<=-16'd3836;
      90679:data<=16'd1785;
      90680:data<=16'd14528;
      90681:data<=16'd18897;
      90682:data<=16'd20522;
      90683:data<=16'd24732;
      90684:data<=16'd23857;
      90685:data<=16'd22453;
      90686:data<=16'd22830;
      90687:data<=16'd20122;
      90688:data<=16'd18716;
      90689:data<=16'd19017;
      90690:data<=16'd17290;
      90691:data<=16'd16064;
      90692:data<=16'd16293;
      90693:data<=16'd17058;
      90694:data<=16'd17290;
      90695:data<=16'd15951;
      90696:data<=16'd14759;
      90697:data<=16'd14054;
      90698:data<=16'd13397;
      90699:data<=16'd12778;
      90700:data<=16'd11271;
      90701:data<=16'd10060;
      90702:data<=16'd9392;
      90703:data<=16'd8768;
      90704:data<=16'd9115;
      90705:data<=16'd8734;
      90706:data<=16'd7758;
      90707:data<=16'd8003;
      90708:data<=16'd7884;
      90709:data<=16'd7204;
      90710:data<=16'd6261;
      90711:data<=16'd5447;
      90712:data<=16'd5815;
      90713:data<=16'd4901;
      90714:data<=16'd3453;
      90715:data<=16'd3623;
      90716:data<=16'd3397;
      90717:data<=16'd3770;
      90718:data<=16'd3277;
      90719:data<=16'd570;
      90720:data<=16'd259;
      90721:data<=-16'd792;
      90722:data<=-16'd2082;
      90723:data<=16'd1011;
      90724:data<=-16'd4100;
      90725:data<=-16'd17259;
      90726:data<=-16'd20157;
      90727:data<=-16'd17236;
      90728:data<=-16'd18190;
      90729:data<=-16'd18007;
      90730:data<=-16'd16583;
      90731:data<=-16'd16486;
      90732:data<=-16'd17408;
      90733:data<=-16'd17807;
      90734:data<=-16'd16442;
      90735:data<=-16'd18889;
      90736:data<=-16'd24236;
      90737:data<=-16'd24077;
      90738:data<=-16'd21899;
      90739:data<=-16'd22137;
      90740:data<=-16'd21284;
      90741:data<=-16'd19801;
      90742:data<=-16'd19309;
      90743:data<=-16'd18820;
      90744:data<=-16'd18017;
      90745:data<=-16'd17532;
      90746:data<=-16'd18251;
      90747:data<=-16'd18390;
      90748:data<=-16'd17191;
      90749:data<=-16'd17130;
      90750:data<=-16'd16960;
      90751:data<=-16'd15223;
      90752:data<=-16'd14712;
      90753:data<=-16'd15212;
      90754:data<=-16'd13828;
      90755:data<=-16'd12126;
      90756:data<=-16'd12320;
      90757:data<=-16'd12043;
      90758:data<=-16'd11492;
      90759:data<=-16'd12859;
      90760:data<=-16'd12724;
      90761:data<=-16'd11074;
      90762:data<=-16'd11624;
      90763:data<=-16'd11861;
      90764:data<=-16'd10822;
      90765:data<=-16'd9644;
      90766:data<=-16'd8530;
      90767:data<=-16'd9909;
      90768:data<=-16'd7001;
      90769:data<=16'd4652;
      90770:data<=16'd11297;
      90771:data<=16'd9081;
      90772:data<=16'd7673;
      90773:data<=16'd7700;
      90774:data<=16'd7844;
      90775:data<=16'd7444;
      90776:data<=16'd5724;
      90777:data<=16'd6213;
      90778:data<=16'd7127;
      90779:data<=16'd6633;
      90780:data<=16'd7359;
      90781:data<=16'd6977;
      90782:data<=16'd6088;
      90783:data<=16'd6498;
      90784:data<=16'd5021;
      90785:data<=16'd3980;
      90786:data<=16'd3968;
      90787:data<=16'd2288;
      90788:data<=16'd4349;
      90789:data<=16'd9824;
      90790:data<=16'd11156;
      90791:data<=16'd9796;
      90792:data<=16'd9412;
      90793:data<=16'd9388;
      90794:data<=16'd9444;
      90795:data<=16'd9062;
      90796:data<=16'd8599;
      90797:data<=16'd8752;
      90798:data<=16'd7477;
      90799:data<=16'd5074;
      90800:data<=16'd5491;
      90801:data<=16'd6672;
      90802:data<=16'd4734;
      90803:data<=16'd4191;
      90804:data<=16'd5441;
      90805:data<=16'd3946;
      90806:data<=16'd3868;
      90807:data<=16'd4792;
      90808:data<=16'd2667;
      90809:data<=16'd2999;
      90810:data<=16'd3541;
      90811:data<=16'd1189;
      90812:data<=16'd2076;
      90813:data<=-16'd2284;
      90814:data<=-16'd15039;
      90815:data<=-16'd18964;
      90816:data<=-16'd15302;
      90817:data<=-16'd15208;
      90818:data<=-16'd15106;
      90819:data<=-16'd14258;
      90820:data<=-16'd14001;
      90821:data<=-16'd12801;
      90822:data<=-16'd12549;
      90823:data<=-16'd11794;
      90824:data<=-16'd10877;
      90825:data<=-16'd12630;
      90826:data<=-16'd13069;
      90827:data<=-16'd11732;
      90828:data<=-16'd11693;
      90829:data<=-16'd11098;
      90830:data<=-16'd10240;
      90831:data<=-16'd10231;
      90832:data<=-16'd9765;
      90833:data<=-16'd8971;
      90834:data<=-16'd8114;
      90835:data<=-16'd7941;
      90836:data<=-16'd7823;
      90837:data<=-16'd6757;
      90838:data<=-16'd8058;
      90839:data<=-16'd9758;
      90840:data<=-16'd7952;
      90841:data<=-16'd9966;
      90842:data<=-16'd16531;
      90843:data<=-16'd17221;
      90844:data<=-16'd14622;
      90845:data<=-16'd15412;
      90846:data<=-16'd14731;
      90847:data<=-16'd12104;
      90848:data<=-16'd11940;
      90849:data<=-16'd11765;
      90850:data<=-16'd10734;
      90851:data<=-16'd11072;
      90852:data<=-16'd11499;
      90853:data<=-16'd11859;
      90854:data<=-16'd11638;
      90855:data<=-16'd10079;
      90856:data<=-16'd10598;
      90857:data<=-16'd9069;
      90858:data<=16'd1298;
      90859:data<=16'd10725;
      90860:data<=16'd10707;
      90861:data<=16'd8930;
      90862:data<=16'd9671;
      90863:data<=16'd9941;
      90864:data<=16'd8526;
      90865:data<=16'd5906;
      90866:data<=16'd5210;
      90867:data<=16'd6435;
      90868:data<=16'd5909;
      90869:data<=16'd5171;
      90870:data<=16'd5404;
      90871:data<=16'd5318;
      90872:data<=16'd6276;
      90873:data<=16'd6636;
      90874:data<=16'd5080;
      90875:data<=16'd4857;
      90876:data<=16'd5251;
      90877:data<=16'd4428;
      90878:data<=16'd3610;
      90879:data<=16'd2625;
      90880:data<=16'd1979;
      90881:data<=16'd1989;
      90882:data<=16'd1747;
      90883:data<=16'd2469;
      90884:data<=16'd3062;
      90885:data<=16'd2250;
      90886:data<=16'd3049;
      90887:data<=16'd4109;
      90888:data<=16'd3072;
      90889:data<=16'd3333;
      90890:data<=16'd4024;
      90891:data<=16'd2664;
      90892:data<=16'd1771;
      90893:data<=16'd808;
      90894:data<=16'd1475;
      90895:data<=16'd7426;
      90896:data<=16'd10925;
      90897:data<=16'd9229;
      90898:data<=16'd9849;
      90899:data<=16'd9227;
      90900:data<=16'd7207;
      90901:data<=16'd10019;
      90902:data<=16'd6237;
      90903:data<=-16'd6830;
      90904:data<=-16'd12214;
      90905:data<=-16'd10687;
      90906:data<=-16'd10753;
      90907:data<=-16'd9724;
      90908:data<=-16'd8933;
      90909:data<=-16'd8998;
      90910:data<=-16'd7661;
      90911:data<=-16'd7565;
      90912:data<=-16'd7924;
      90913:data<=-16'd7306;
      90914:data<=-16'd7101;
      90915:data<=-16'd6460;
      90916:data<=-16'd6296;
      90917:data<=-16'd6520;
      90918:data<=-16'd5426;
      90919:data<=-16'd4720;
      90920:data<=-16'd4090;
      90921:data<=-16'd3162;
      90922:data<=-16'd3407;
      90923:data<=-16'd2924;
      90924:data<=-16'd1741;
      90925:data<=-16'd1726;
      90926:data<=-16'd1764;
      90927:data<=-16'd1357;
      90928:data<=-16'd802;
      90929:data<=-16'd470;
      90930:data<=-16'd490;
      90931:data<=16'd92;
      90932:data<=16'd969;
      90933:data<=16'd1539;
      90934:data<=16'd1228;
      90935:data<=16'd829;
      90936:data<=16'd2264;
      90937:data<=16'd2676;
      90938:data<=16'd1453;
      90939:data<=16'd1932;
      90940:data<=16'd1892;
      90941:data<=16'd1451;
      90942:data<=16'd2147;
      90943:data<=16'd1503;
      90944:data<=16'd2517;
      90945:data<=16'd4440;
      90946:data<=16'd3970;
      90947:data<=16'd8384;
      90948:data<=16'd15209;
      90949:data<=16'd14636;
      90950:data<=16'd12145;
      90951:data<=16'd12340;
      90952:data<=16'd11802;
      90953:data<=16'd10969;
      90954:data<=16'd10693;
      90955:data<=16'd10577;
      90956:data<=16'd10345;
      90957:data<=16'd10495;
      90958:data<=16'd11558;
      90959:data<=16'd11282;
      90960:data<=16'd10546;
      90961:data<=16'd10968;
      90962:data<=16'd10372;
      90963:data<=16'd10111;
      90964:data<=16'd10226;
      90965:data<=16'd8343;
      90966:data<=16'd7450;
      90967:data<=16'd8061;
      90968:data<=16'd7808;
      90969:data<=16'd7674;
      90970:data<=16'd7909;
      90971:data<=16'd8540;
      90972:data<=16'd9098;
      90973:data<=16'd8257;
      90974:data<=16'd7567;
      90975:data<=16'd7796;
      90976:data<=16'd7699;
      90977:data<=16'd7142;
      90978:data<=16'd6901;
      90979:data<=16'd6784;
      90980:data<=16'd5468;
      90981:data<=16'd4881;
      90982:data<=16'd5548;
      90983:data<=16'd4611;
      90984:data<=16'd5072;
      90985:data<=16'd6795;
      90986:data<=16'd6141;
      90987:data<=16'd7056;
      90988:data<=16'd7119;
      90989:data<=16'd4763;
      90990:data<=16'd6918;
      90991:data<=16'd4306;
      90992:data<=-16'd7991;
      90993:data<=-16'd13659;
      90994:data<=-16'd11723;
      90995:data<=-16'd11564;
      90996:data<=-16'd11624;
      90997:data<=-16'd10683;
      90998:data<=-16'd8978;
      90999:data<=-16'd8185;
      91000:data<=-16'd7779;
      91001:data<=-16'd2358;
      91002:data<=16'd2290;
      91003:data<=16'd547;
      91004:data<=-16'd146;
      91005:data<=16'd986;
      91006:data<=16'd511;
      91007:data<=16'd716;
      91008:data<=16'd1099;
      91009:data<=16'd711;
      91010:data<=16'd1162;
      91011:data<=16'd2781;
      91012:data<=16'd3908;
      91013:data<=16'd3392;
      91014:data<=16'd3629;
      91015:data<=16'd4501;
      91016:data<=16'd3492;
      91017:data<=16'd2648;
      91018:data<=16'd2710;
      91019:data<=16'd2347;
      91020:data<=16'd2073;
      91021:data<=16'd1829;
      91022:data<=16'd2062;
      91023:data<=16'd2177;
      91024:data<=16'd2608;
      91025:data<=16'd4983;
      91026:data<=16'd5203;
      91027:data<=16'd3914;
      91028:data<=16'd5178;
      91029:data<=16'd4572;
      91030:data<=16'd3648;
      91031:data<=16'd4705;
      91032:data<=16'd2661;
      91033:data<=16'd2737;
      91034:data<=16'd4405;
      91035:data<=16'd1071;
      91036:data<=16'd6072;
      91037:data<=16'd19746;
      91038:data<=16'd22735;
      91039:data<=16'd19358;
      91040:data<=16'd19892;
      91041:data<=16'd19203;
      91042:data<=16'd17285;
      91043:data<=16'd16654;
      91044:data<=16'd15948;
      91045:data<=16'd15220;
      91046:data<=16'd13867;
      91047:data<=16'd13029;
      91048:data<=16'd13762;
      91049:data<=16'd13811;
      91050:data<=16'd12872;
      91051:data<=16'd12175;
      91052:data<=16'd12577;
      91053:data<=16'd12468;
      91054:data<=16'd8050;
      91055:data<=16'd2319;
      91056:data<=16'd760;
      91057:data<=16'd1171;
      91058:data<=16'd622;
      91059:data<=16'd199;
      91060:data<=16'd343;
      91061:data<=-16'd33;
      91062:data<=-16'd811;
      91063:data<=16'd94;
      91064:data<=16'd1932;
      91065:data<=16'd1762;
      91066:data<=16'd795;
      91067:data<=16'd928;
      91068:data<=16'd1133;
      91069:data<=16'd617;
      91070:data<=-16'd364;
      91071:data<=-16'd901;
      91072:data<=-16'd807;
      91073:data<=-16'd858;
      91074:data<=-16'd1300;
      91075:data<=-16'd1864;
      91076:data<=-16'd1083;
      91077:data<=16'd206;
      91078:data<=16'd32;
      91079:data<=16'd881;
      91080:data<=-16'd977;
      91081:data<=-16'd11104;
      91082:data<=-16'd18842;
      91083:data<=-16'd17566;
      91084:data<=-16'd16349;
      91085:data<=-16'd17194;
      91086:data<=-16'd16894;
      91087:data<=-16'd15961;
      91088:data<=-16'd14521;
      91089:data<=-16'd14389;
      91090:data<=-16'd14051;
      91091:data<=-16'd11482;
      91092:data<=-16'd10843;
      91093:data<=-16'd11238;
      91094:data<=-16'd10369;
      91095:data<=-16'd10589;
      91096:data<=-16'd10063;
      91097:data<=-16'd8862;
      91098:data<=-16'd9059;
      91099:data<=-16'd8519;
      91100:data<=-16'd8146;
      91101:data<=-16'd8087;
      91102:data<=-16'd6936;
      91103:data<=-16'd6513;
      91104:data<=-16'd5093;
      91105:data<=-16'd3800;
      91106:data<=-16'd5228;
      91107:data<=-16'd2191;
      91108:data<=16'd4123;
      91109:data<=16'd3933;
      91110:data<=16'd2088;
      91111:data<=16'd4162;
      91112:data<=16'd4502;
      91113:data<=16'd3377;
      91114:data<=16'd4200;
      91115:data<=16'd3864;
      91116:data<=16'd3187;
      91117:data<=16'd5106;
      91118:data<=16'd5700;
      91119:data<=16'd4852;
      91120:data<=16'd5266;
      91121:data<=16'd4247;
      91122:data<=16'd4082;
      91123:data<=16'd4831;
      91124:data<=16'd1936;
      91125:data<=16'd5752;
      91126:data<=16'd18167;
      91127:data<=16'd21634;
      91128:data<=16'd18037;
      91129:data<=16'd18157;
      91130:data<=16'd18137;
      91131:data<=16'd17514;
      91132:data<=16'd17012;
      91133:data<=16'd15018;
      91134:data<=16'd14622;
      91135:data<=16'd14304;
      91136:data<=16'd13167;
      91137:data<=16'd13527;
      91138:data<=16'd12575;
      91139:data<=16'd11018;
      91140:data<=16'd10780;
      91141:data<=16'd9871;
      91142:data<=16'd9265;
      91143:data<=16'd8316;
      91144:data<=16'd6199;
      91145:data<=16'd5300;
      91146:data<=16'd4534;
      91147:data<=16'd3516;
      91148:data<=16'd3606;
      91149:data<=16'd3738;
      91150:data<=16'd3356;
      91151:data<=16'd2153;
      91152:data<=16'd1621;
      91153:data<=16'd2767;
      91154:data<=16'd2620;
      91155:data<=16'd1894;
      91156:data<=16'd1404;
      91157:data<=-16'd1413;
      91158:data<=-16'd3071;
      91159:data<=-16'd1744;
      91160:data<=-16'd3876;
      91161:data<=-16'd9922;
      91162:data<=-16'd12313;
      91163:data<=-16'd10490;
      91164:data<=-16'd10772;
      91165:data<=-16'd11559;
      91166:data<=-16'd9969;
      91167:data<=-16'd10753;
      91168:data<=-16'd11035;
      91169:data<=-16'd9456;
      91170:data<=-16'd16944;
      91171:data<=-16'd28268;
      91172:data<=-16'd29561;
      91173:data<=-16'd26821;
      91174:data<=-16'd26536;
      91175:data<=-16'd25642;
      91176:data<=-16'd24697;
      91177:data<=-16'd24005;
      91178:data<=-16'd22664;
      91179:data<=-16'd21440;
      91180:data<=-16'd20657;
      91181:data<=-16'd20854;
      91182:data<=-16'd21102;
      91183:data<=-16'd20562;
      91184:data<=-16'd20218;
      91185:data<=-16'd19840;
      91186:data<=-16'd19394;
      91187:data<=-16'd18951;
      91188:data<=-16'd17888;
      91189:data<=-16'd16826;
      91190:data<=-16'd15954;
      91191:data<=-16'd15083;
      91192:data<=-16'd14210;
      91193:data<=-16'd13048;
      91194:data<=-16'd12220;
      91195:data<=-16'd11724;
      91196:data<=-16'd11934;
      91197:data<=-16'd13324;
      91198:data<=-16'd13220;
      91199:data<=-16'd11486;
      91200:data<=-16'd11124;
      91201:data<=-16'd11318;
      91202:data<=-16'd10276;
      91203:data<=-16'd8610;
      91204:data<=-16'd7641;
      91205:data<=-16'd7700;
      91206:data<=-16'd7682;
      91207:data<=-16'd7075;
      91208:data<=-16'd5909;
      91209:data<=-16'd5785;
      91210:data<=-16'd7259;
      91211:data<=-16'd6728;
      91212:data<=-16'd6405;
      91213:data<=-16'd6616;
      91214:data<=16'd3360;
      91215:data<=16'd17728;
      91216:data<=16'd20865;
      91217:data<=16'd19531;
      91218:data<=16'd20354;
      91219:data<=16'd18539;
      91220:data<=16'd17713;
      91221:data<=16'd18606;
      91222:data<=16'd16907;
      91223:data<=16'd15255;
      91224:data<=16'd14283;
      91225:data<=16'd13362;
      91226:data<=16'd13841;
      91227:data<=16'd13565;
      91228:data<=16'd12342;
      91229:data<=16'd11806;
      91230:data<=16'd11286;
      91231:data<=16'd11051;
      91232:data<=16'd10796;
      91233:data<=16'd9938;
      91234:data<=16'd9429;
      91235:data<=16'd8983;
      91236:data<=16'd7946;
      91237:data<=16'd6567;
      91238:data<=16'd5651;
      91239:data<=16'd5667;
      91240:data<=16'd5785;
      91241:data<=16'd5903;
      91242:data<=16'd5749;
      91243:data<=16'd4931;
      91244:data<=16'd4846;
      91245:data<=16'd4843;
      91246:data<=16'd3921;
      91247:data<=16'd3333;
      91248:data<=16'd2723;
      91249:data<=16'd1982;
      91250:data<=16'd1096;
      91251:data<=-16'd208;
      91252:data<=16'd111;
      91253:data<=16'd440;
      91254:data<=-16'd227;
      91255:data<=16'd902;
      91256:data<=16'd62;
      91257:data<=-16'd1422;
      91258:data<=16'd1562;
      91259:data<=-16'd2611;
      91260:data<=-16'd15359;
      91261:data<=-16'd18722;
      91262:data<=-16'd15596;
      91263:data<=-16'd17705;
      91264:data<=-16'd18659;
      91265:data<=-16'd16340;
      91266:data<=-16'd17764;
      91267:data<=-16'd22024;
      91268:data<=-16'd23890;
      91269:data<=-16'd22527;
      91270:data<=-16'd21294;
      91271:data<=-16'd20970;
      91272:data<=-16'd19273;
      91273:data<=-16'd17631;
      91274:data<=-16'd17280;
      91275:data<=-16'd16633;
      91276:data<=-16'd16266;
      91277:data<=-16'd16706;
      91278:data<=-16'd16422;
      91279:data<=-16'd14916;
      91280:data<=-16'd13581;
      91281:data<=-16'd13242;
      91282:data<=-16'd12574;
      91283:data<=-16'd11303;
      91284:data<=-16'd10285;
      91285:data<=-16'd9351;
      91286:data<=-16'd9207;
      91287:data<=-16'd9439;
      91288:data<=-16'd8827;
      91289:data<=-16'd8824;
      91290:data<=-16'd9480;
      91291:data<=-16'd9356;
      91292:data<=-16'd8837;
      91293:data<=-16'd8094;
      91294:data<=-16'd6987;
      91295:data<=-16'd5802;
      91296:data<=-16'd5285;
      91297:data<=-16'd5084;
      91298:data<=-16'd4017;
      91299:data<=-16'd3849;
      91300:data<=-16'd3544;
      91301:data<=-16'd2079;
      91302:data<=-16'd4322;
      91303:data<=-16'd3576;
      91304:data<=16'd7201;
      91305:data<=16'd14038;
      91306:data<=16'd12827;
      91307:data<=16'd13423;
      91308:data<=16'd13317;
      91309:data<=16'd12236;
      91310:data<=16'd13339;
      91311:data<=16'd12542;
      91312:data<=16'd11764;
      91313:data<=16'd12490;
      91314:data<=16'd11517;
      91315:data<=16'd10787;
      91316:data<=16'd10539;
      91317:data<=16'd9747;
      91318:data<=16'd9201;
      91319:data<=16'd9370;
      91320:data<=16'd12649;
      91321:data<=16'd15656;
      91322:data<=16'd14381;
      91323:data<=16'd13720;
      91324:data<=16'd14304;
      91325:data<=16'd13438;
      91326:data<=16'd12719;
      91327:data<=16'd12211;
      91328:data<=16'd11565;
      91329:data<=16'd10213;
      91330:data<=16'd8784;
      91331:data<=16'd9374;
      91332:data<=16'd9303;
      91333:data<=16'd8378;
      91334:data<=16'd8517;
      91335:data<=16'd7215;
      91336:data<=16'd6273;
      91337:data<=16'd7183;
      91338:data<=16'd6921;
      91339:data<=16'd5888;
      91340:data<=16'd5087;
      91341:data<=16'd5782;
      91342:data<=16'd6912;
      91343:data<=16'd5938;
      91344:data<=16'd6038;
      91345:data<=16'd5262;
      91346:data<=16'd3557;
      91347:data<=16'd6560;
      91348:data<=16'd2596;
      91349:data<=-16'd10765;
      91350:data<=-16'd14381;
      91351:data<=-16'd11104;
      91352:data<=-16'd11424;
      91353:data<=-16'd10947;
      91354:data<=-16'd10608;
      91355:data<=-16'd9962;
      91356:data<=-16'd7254;
      91357:data<=-16'd7312;
      91358:data<=-16'd7988;
      91359:data<=-16'd7491;
      91360:data<=-16'd7811;
      91361:data<=-16'd6916;
      91362:data<=-16'd6128;
      91363:data<=-16'd6070;
      91364:data<=-16'd5360;
      91365:data<=-16'd5529;
      91366:data<=-16'd5171;
      91367:data<=-16'd4217;
      91368:data<=-16'd3764;
      91369:data<=-16'd2272;
      91370:data<=-16'd1739;
      91371:data<=-16'd2109;
      91372:data<=-16'd1989;
      91373:data<=-16'd4168;
      91374:data<=-16'd6808;
      91375:data<=-16'd7321;
      91376:data<=-16'd7365;
      91377:data<=-16'd7142;
      91378:data<=-16'd6708;
      91379:data<=-16'd5497;
      91380:data<=-16'd4046;
      91381:data<=-16'd4270;
      91382:data<=-16'd3794;
      91383:data<=-16'd2138;
      91384:data<=-16'd1391;
      91385:data<=-16'd934;
      91386:data<=-16'd1108;
      91387:data<=-16'd1031;
      91388:data<=-16'd306;
      91389:data<=-16'd297;
      91390:data<=16'd346;
      91391:data<=-16'd341;
      91392:data<=16'd21;
      91393:data<=16'd8959;
      91394:data<=16'd17852;
      91395:data<=16'd18316;
      91396:data<=16'd18120;
      91397:data<=16'd18830;
      91398:data<=16'd17873;
      91399:data<=16'd17587;
      91400:data<=16'd17000;
      91401:data<=16'd16322;
      91402:data<=16'd16204;
      91403:data<=16'd14879;
      91404:data<=16'd14275;
      91405:data<=16'd14910;
      91406:data<=16'd14404;
      91407:data<=16'd13294;
      91408:data<=16'd13277;
      91409:data<=16'd14457;
      91410:data<=16'd14628;
      91411:data<=16'd13449;
      91412:data<=16'd13019;
      91413:data<=16'd12483;
      91414:data<=16'd12047;
      91415:data<=16'd12551;
      91416:data<=16'd11605;
      91417:data<=16'd10217;
      91418:data<=16'd10128;
      91419:data<=16'd9677;
      91420:data<=16'd9251;
      91421:data<=16'd9279;
      91422:data<=16'd9236;
      91423:data<=16'd9550;
      91424:data<=16'd8998;
      91425:data<=16'd7909;
      91426:data<=16'd9746;
      91427:data<=16'd13970;
      91428:data<=16'd14904;
      91429:data<=16'd12181;
      91430:data<=16'd11445;
      91431:data<=16'd11480;
      91432:data<=16'd10329;
      91433:data<=16'd11126;
      91434:data<=16'd9947;
      91435:data<=16'd8122;
      91436:data<=16'd11849;
      91437:data<=16'd8777;
      91438:data<=-16'd3908;
      91439:data<=-16'd8296;
      91440:data<=-16'd6347;
      91441:data<=-16'd7539;
      91442:data<=-16'd7286;
      91443:data<=-16'd6934;
      91444:data<=-16'd8419;
      91445:data<=-16'd7912;
      91446:data<=-16'd7280;
      91447:data<=-16'd7048;
      91448:data<=-16'd5500;
      91449:data<=-16'd4420;
      91450:data<=-16'd4299;
      91451:data<=-16'd4228;
      91452:data<=-16'd3739;
      91453:data<=-16'd3771;
      91454:data<=-16'd4730;
      91455:data<=-16'd4417;
      91456:data<=-16'd3853;
      91457:data<=-16'd4273;
      91458:data<=-16'd3900;
      91459:data<=-16'd4115;
      91460:data<=-16'd4943;
      91461:data<=-16'd4143;
      91462:data<=-16'd2811;
      91463:data<=-16'd1782;
      91464:data<=-16'd1767;
      91465:data<=-16'd2253;
      91466:data<=-16'd1327;
      91467:data<=-16'd1506;
      91468:data<=-16'd2666;
      91469:data<=-16'd1874;
      91470:data<=-16'd1583;
      91471:data<=-16'd1838;
      91472:data<=-16'd1204;
      91473:data<=-16'd1434;
      91474:data<=-16'd1008;
      91475:data<=16'd149;
      91476:data<=16'd0;
      91477:data<=16'd105;
      91478:data<=16'd296;
      91479:data<=-16'd1289;
      91480:data<=-16'd5604;
      91481:data<=-16'd8619;
      91482:data<=-16'd1497;
      91483:data<=16'd9687;
      91484:data<=16'd11358;
      91485:data<=16'd8933;
      91486:data<=16'd9850;
      91487:data<=16'd10052;
      91488:data<=16'd9956;
      91489:data<=16'd11127;
      91490:data<=16'd10921;
      91491:data<=16'd9705;
      91492:data<=16'd8971;
      91493:data<=16'd8927;
      91494:data<=16'd9195;
      91495:data<=16'd8934;
      91496:data<=16'd8081;
      91497:data<=16'd7040;
      91498:data<=16'd6872;
      91499:data<=16'd7195;
      91500:data<=16'd6361;
      91501:data<=16'd6035;
      91502:data<=16'd7057;
      91503:data<=16'd7315;
      91504:data<=16'd7192;
      91505:data<=16'd7468;
      91506:data<=16'd7051;
      91507:data<=16'd5891;
      91508:data<=16'd5309;
      91509:data<=16'd5492;
      91510:data<=16'd4937;
      91511:data<=16'd4451;
      91512:data<=16'd4825;
      91513:data<=16'd3953;
      91514:data<=16'd3471;
      91515:data<=16'd4596;
      91516:data<=16'd4252;
      91517:data<=16'd3750;
      91518:data<=16'd4478;
      91519:data<=16'd4243;
      91520:data<=16'd3500;
      91521:data<=16'd3137;
      91522:data<=16'd3136;
      91523:data<=16'd2309;
      91524:data<=16'd1293;
      91525:data<=16'd3163;
      91526:data<=16'd262;
      91527:data<=-16'd11392;
      91528:data<=-16'd16751;
      91529:data<=-16'd13215;
      91530:data<=-16'd12533;
      91531:data<=-16'd13132;
      91532:data<=-16'd10486;
      91533:data<=-16'd6617;
      91534:data<=-16'd4507;
      91535:data<=-16'd5724;
      91536:data<=-16'd6288;
      91537:data<=-16'd5043;
      91538:data<=-16'd4874;
      91539:data<=-16'd4851;
      91540:data<=-16'd5485;
      91541:data<=-16'd5632;
      91542:data<=-16'd3550;
      91543:data<=-16'd3081;
      91544:data<=-16'd3447;
      91545:data<=-16'd2895;
      91546:data<=-16'd3212;
      91547:data<=-16'd2413;
      91548:data<=-16'd1897;
      91549:data<=-16'd3386;
      91550:data<=-16'd3497;
      91551:data<=-16'd3096;
      91552:data<=-16'd2983;
      91553:data<=-16'd2366;
      91554:data<=-16'd2587;
      91555:data<=-16'd2732;
      91556:data<=-16'd2942;
      91557:data<=-16'd3048;
      91558:data<=-16'd2044;
      91559:data<=-16'd2164;
      91560:data<=-16'd2320;
      91561:data<=-16'd1980;
      91562:data<=-16'd2513;
      91563:data<=-16'd2041;
      91564:data<=-16'd2921;
      91565:data<=-16'd4044;
      91566:data<=-16'd2100;
      91567:data<=-16'd2977;
      91568:data<=-16'd4540;
      91569:data<=-16'd3926;
      91570:data<=-16'd5973;
      91571:data<=-16'd1057;
      91572:data<=16'd11245;
      91573:data<=16'd13778;
      91574:data<=16'd10742;
      91575:data<=16'd11489;
      91576:data<=16'd10994;
      91577:data<=16'd10075;
      91578:data<=16'd10539;
      91579:data<=16'd9639;
      91580:data<=16'd8254;
      91581:data<=16'd7151;
      91582:data<=16'd5700;
      91583:data<=16'd4602;
      91584:data<=16'd5071;
      91585:data<=16'd4009;
      91586:data<=-16'd960;
      91587:data<=-16'd3112;
      91588:data<=-16'd1663;
      91589:data<=-16'd2425;
      91590:data<=-16'd2707;
      91591:data<=-16'd2607;
      91592:data<=-16'd3999;
      91593:data<=-16'd3018;
      91594:data<=-16'd2655;
      91595:data<=-16'd4670;
      91596:data<=-16'd4896;
      91597:data<=-16'd4781;
      91598:data<=-16'd4722;
      91599:data<=-16'd4355;
      91600:data<=-16'd5216;
      91601:data<=-16'd4770;
      91602:data<=-16'd3927;
      91603:data<=-16'd4875;
      91604:data<=-16'd5112;
      91605:data<=-16'd4587;
      91606:data<=-16'd4267;
      91607:data<=-16'd5016;
      91608:data<=-16'd6811;
      91609:data<=-16'd6757;
      91610:data<=-16'd6061;
      91611:data<=-16'd5962;
      91612:data<=-16'd5749;
      91613:data<=-16'd6746;
      91614:data<=-16'd5796;
      91615:data<=-16'd5918;
      91616:data<=-16'd15003;
      91617:data<=-16'd23090;
      91618:data<=-16'd21910;
      91619:data<=-16'd19975;
      91620:data<=-16'd19917;
      91621:data<=-16'd19957;
      91622:data<=-16'd20905;
      91623:data<=-16'd20720;
      91624:data<=-16'd19735;
      91625:data<=-16'd18841;
      91626:data<=-16'd17497;
      91627:data<=-16'd17162;
      91628:data<=-16'd17076;
      91629:data<=-16'd16152;
      91630:data<=-16'd15127;
      91631:data<=-16'd14146;
      91632:data<=-16'd13690;
      91633:data<=-16'd13127;
      91634:data<=-16'd12777;
      91635:data<=-16'd13342;
      91636:data<=-16'd12859;
      91637:data<=-16'd12454;
      91638:data<=-16'd11925;
      91639:data<=-16'd7829;
      91640:data<=-16'd4179;
      91641:data<=-16'd4199;
      91642:data<=-16'd4284;
      91643:data<=-16'd3748;
      91644:data<=-16'd3240;
      91645:data<=-16'd2689;
      91646:data<=-16'd2576;
      91647:data<=-16'd2737;
      91648:data<=-16'd3635;
      91649:data<=-16'd3795;
      91650:data<=-16'd2922;
      91651:data<=-16'd3430;
      91652:data<=-16'd3392;
      91653:data<=-16'd2319;
      91654:data<=-16'd2279;
      91655:data<=-16'd2121;
      91656:data<=-16'd2033;
      91657:data<=-16'd983;
      91658:data<=-16'd227;
      91659:data<=-16'd2804;
      91660:data<=16'd1130;
      91661:data<=16'd12502;
      91662:data<=16'd15282;
      91663:data<=16'd12254;
      91664:data<=16'd13062;
      91665:data<=16'd12775;
      91666:data<=16'd11693;
      91667:data<=16'd12213;
      91668:data<=16'd11844;
      91669:data<=16'd11762;
      91670:data<=16'd11179;
      91671:data<=16'd10041;
      91672:data<=16'd10615;
      91673:data<=16'd10257;
      91674:data<=16'd8481;
      91675:data<=16'd7147;
      91676:data<=16'd6432;
      91677:data<=16'd7188;
      91678:data<=16'd7301;
      91679:data<=16'd6062;
      91680:data<=16'd5832;
      91681:data<=16'd5488;
      91682:data<=16'd5565;
      91683:data<=16'd6601;
      91684:data<=16'd5796;
      91685:data<=16'd4570;
      91686:data<=16'd4501;
      91687:data<=16'd4173;
      91688:data<=16'd3248;
      91689:data<=16'd1733;
      91690:data<=16'd1791;
      91691:data<=16'd2385;
      91692:data<=-16'd934;
      91693:data<=-16'd4420;
      91694:data<=-16'd4634;
      91695:data<=-16'd4485;
      91696:data<=-16'd3704;
      91697:data<=-16'd3046;
      91698:data<=-16'd4058;
      91699:data<=-16'd4205;
      91700:data<=-16'd3576;
      91701:data<=-16'd4112;
      91702:data<=-16'd5535;
      91703:data<=-16'd5169;
      91704:data<=-16'd3808;
      91705:data<=-16'd10122;
      91706:data<=-16'd20968;
      91707:data<=-16'd22618;
      91708:data<=-16'd19141;
      91709:data<=-16'd18854;
      91710:data<=-16'd18351;
      91711:data<=-16'd17405;
      91712:data<=-16'd16718;
      91713:data<=-16'd16107;
      91714:data<=-16'd17431;
      91715:data<=-16'd17270;
      91716:data<=-16'd15371;
      91717:data<=-16'd15382;
      91718:data<=-16'd14882;
      91719:data<=-16'd13450;
      91720:data<=-16'd12813;
      91721:data<=-16'd11982;
      91722:data<=-16'd11435;
      91723:data<=-16'd10934;
      91724:data<=-16'd10066;
      91725:data<=-16'd9168;
      91726:data<=-16'd8238;
      91727:data<=-16'd9003;
      91728:data<=-16'd9999;
      91729:data<=-16'd9013;
      91730:data<=-16'd8311;
      91731:data<=-16'd8087;
      91732:data<=-16'd7905;
      91733:data<=-16'd7882;
      91734:data<=-16'd6746;
      91735:data<=-16'd6087;
      91736:data<=-16'd5636;
      91737:data<=-16'd4328;
      91738:data<=-16'd4259;
      91739:data<=-16'd3654;
      91740:data<=-16'd2911;
      91741:data<=-16'd4575;
      91742:data<=-16'd4407;
      91743:data<=-16'd2925;
      91744:data<=-16'd3826;
      91745:data<=-16'd2159;
      91746:data<=16'd3527;
      91747:data<=16'd5359;
      91748:data<=16'd2437;
      91749:data<=16'd6640;
      91750:data<=16'd18891;
      91751:data<=16'd23388;
      91752:data<=16'd20248;
      91753:data<=16'd20064;
      91754:data<=16'd19203;
      91755:data<=16'd17205;
      91756:data<=16'd17506;
      91757:data<=16'd16554;
      91758:data<=16'd16137;
      91759:data<=16'd16904;
      91760:data<=16'd15790;
      91761:data<=16'd15405;
      91762:data<=16'd15057;
      91763:data<=16'd13817;
      91764:data<=16'd14139;
      91765:data<=16'd13776;
      91766:data<=16'd12580;
      91767:data<=16'd12349;
      91768:data<=16'd11797;
      91769:data<=16'd11276;
      91770:data<=16'd10771;
      91771:data<=16'd10413;
      91772:data<=16'd11013;
      91773:data<=16'd10874;
      91774:data<=16'd9820;
      91775:data<=16'd8790;
      91776:data<=16'd8652;
      91777:data<=16'd9662;
      91778:data<=16'd9186;
      91779:data<=16'd8263;
      91780:data<=16'd8913;
      91781:data<=16'd9092;
      91782:data<=16'd9480;
      91783:data<=16'd9656;
      91784:data<=16'd8460;
      91785:data<=16'd8457;
      91786:data<=16'd8205;
      91787:data<=16'd7194;
      91788:data<=16'd7489;
      91789:data<=16'd7194;
      91790:data<=16'd7125;
      91791:data<=16'd6769;
      91792:data<=16'd5573;
      91793:data<=16'd7506;
      91794:data<=16'd3943;
      91795:data<=-16'd8519;
      91796:data<=-16'd11999;
      91797:data<=-16'd7398;
      91798:data<=-16'd10172;
      91799:data<=-16'd15088;
      91800:data<=-16'd15350;
      91801:data<=-16'd14493;
      91802:data<=-16'd13503;
      91803:data<=-16'd13095;
      91804:data<=-16'd13092;
      91805:data<=-16'd12242;
      91806:data<=-16'd11194;
      91807:data<=-16'd9679;
      91808:data<=-16'd8624;
      91809:data<=-16'd8402;
      91810:data<=-16'd7304;
      91811:data<=-16'd6663;
      91812:data<=-16'd6866;
      91813:data<=-16'd6466;
      91814:data<=-16'd6150;
      91815:data<=-16'd5285;
      91816:data<=-16'd4237;
      91817:data<=-16'd4986;
      91818:data<=-16'd5368;
      91819:data<=-16'd4108;
      91820:data<=-16'd3049;
      91821:data<=-16'd1898;
      91822:data<=-16'd1022;
      91823:data<=-16'd1710;
      91824:data<=-16'd2096;
      91825:data<=-16'd1413;
      91826:data<=-16'd1407;
      91827:data<=-16'd1222;
      91828:data<=-16'd224;
      91829:data<=-16'd227;
      91830:data<=-16'd293;
      91831:data<=16'd523;
      91832:data<=16'd522;
      91833:data<=16'd604;
      91834:data<=16'd1704;
      91835:data<=16'd2790;
      91836:data<=16'd3095;
      91837:data<=16'd1551;
      91838:data<=16'd3419;
      91839:data<=16'd13526;
      91840:data<=16'd21056;
      91841:data<=16'd19070;
      91842:data<=16'd17094;
      91843:data<=16'd18210;
      91844:data<=16'd17616;
      91845:data<=16'd16581;
      91846:data<=16'd16927;
      91847:data<=16'd17202;
      91848:data<=16'd17079;
      91849:data<=16'd16933;
      91850:data<=16'd16375;
      91851:data<=16'd16865;
      91852:data<=16'd19828;
      91853:data<=16'd21494;
      91854:data<=16'd20269;
      91855:data<=16'd19603;
      91856:data<=16'd18591;
      91857:data<=16'd16677;
      91858:data<=16'd16531;
      91859:data<=16'd16873;
      91860:data<=16'd16909;
      91861:data<=16'd16960;
      91862:data<=16'd15867;
      91863:data<=16'd14822;
      91864:data<=16'd14240;
      91865:data<=16'd13720;
      91866:data<=16'd13609;
      91867:data<=16'd12736;
      91868:data<=16'd11815;
      91869:data<=16'd11330;
      91870:data<=16'd10463;
      91871:data<=16'd10075;
      91872:data<=16'd9435;
      91873:data<=16'd9644;
      91874:data<=16'd10883;
      91875:data<=16'd9409;
      91876:data<=16'd8505;
      91877:data<=16'd9471;
      91878:data<=16'd8363;
      91879:data<=16'd8440;
      91880:data<=16'd8243;
      91881:data<=16'd6451;
      91882:data<=16'd7843;
      91883:data<=16'd2855;
      91884:data<=-16'd9906;
      91885:data<=-16'd13474;
      91886:data<=-16'd10151;
      91887:data<=-16'd9618;
      91888:data<=-16'd9189;
      91889:data<=-16'd9471;
      91890:data<=-16'd9855;
      91891:data<=-16'd8348;
      91892:data<=-16'd8184;
      91893:data<=-16'd8599;
      91894:data<=-16'd8392;
      91895:data<=-16'd8542;
      91896:data<=-16'd8319;
      91897:data<=-16'd8658;
      91898:data<=-16'd8962;
      91899:data<=-16'd7779;
      91900:data<=-16'd6560;
      91901:data<=-16'd6002;
      91902:data<=-16'd5917;
      91903:data<=-16'd5591;
      91904:data<=-16'd6522;
      91905:data<=-16'd10674;
      91906:data<=-16'd13018;
      91907:data<=-16'd11659;
      91908:data<=-16'd11408;
      91909:data<=-16'd11966;
      91910:data<=-16'd11790;
      91911:data<=-16'd11025;
      91912:data<=-16'd9350;
      91913:data<=-16'd8481;
      91914:data<=-16'd7997;
      91915:data<=-16'd7447;
      91916:data<=-16'd7626;
      91917:data<=-16'd6487;
      91918:data<=-16'd5844;
      91919:data<=-16'd6996;
      91920:data<=-16'd6469;
      91921:data<=-16'd5823;
      91922:data<=-16'd6131;
      91923:data<=-16'd6055;
      91924:data<=-16'd6311;
      91925:data<=-16'd4939;
      91926:data<=-16'd3829;
      91927:data<=-16'd2723;
      91928:data<=16'd5835;
      91929:data<=16'd14380;
      91930:data<=16'd13524;
      91931:data<=16'd11621;
      91932:data<=16'd11955;
      91933:data<=16'd11276;
      91934:data<=16'd10771;
      91935:data<=16'd9991;
      91936:data<=16'd10032;
      91937:data<=16'd10376;
      91938:data<=16'd8921;
      91939:data<=16'd9310;
      91940:data<=16'd10760;
      91941:data<=16'd10293;
      91942:data<=16'd9953;
      91943:data<=16'd9119;
      91944:data<=16'd8034;
      91945:data<=16'd7530;
      91946:data<=16'd6229;
      91947:data<=16'd6231;
      91948:data<=16'd6587;
      91949:data<=16'd5403;
      91950:data<=16'd5536;
      91951:data<=16'd5758;
      91952:data<=16'd5192;
      91953:data<=16'd5859;
      91954:data<=16'd6422;
      91955:data<=16'd6384;
      91956:data<=16'd5456;
      91957:data<=16'd5260;
      91958:data<=16'd8848;
      91959:data<=16'd11473;
      91960:data<=16'd10314;
      91961:data<=16'd9257;
      91962:data<=16'd8792;
      91963:data<=16'd8549;
      91964:data<=16'd8340;
      91965:data<=16'd8023;
      91966:data<=16'd8226;
      91967:data<=16'd7662;
      91968:data<=16'd7621;
      91969:data<=16'd7357;
      91970:data<=16'd5576;
      91971:data<=16'd6493;
      91972:data<=16'd3535;
      91973:data<=-16'd7060;
      91974:data<=-16'd10963;
      91975:data<=-16'd8434;
      91976:data<=-16'd9133;
      91977:data<=-16'd9432;
      91978:data<=-16'd8851;
      91979:data<=-16'd8570;
      91980:data<=-16'd7759;
      91981:data<=-16'd8830;
      91982:data<=-16'd8984;
      91983:data<=-16'd8050;
      91984:data<=-16'd8352;
      91985:data<=-16'd7574;
      91986:data<=-16'd8116;
      91987:data<=-16'd8796;
      91988:data<=-16'd6907;
      91989:data<=-16'd7518;
      91990:data<=-16'd7994;
      91991:data<=-16'd6307;
      91992:data<=-16'd7410;
      91993:data<=-16'd8346;
      91994:data<=-16'd8307;
      91995:data<=-16'd8975;
      91996:data<=-16'd8053;
      91997:data<=-16'd7814;
      91998:data<=-16'd7755;
      91999:data<=-16'd6831;
      92000:data<=-16'd7724;
      92001:data<=-16'd7583;
      92002:data<=-16'd7118;
      92003:data<=-16'd7867;
      92004:data<=-16'd6689;
      92005:data<=-16'd7175;
      92006:data<=-16'd8947;
      92007:data<=-16'd8370;
      92008:data<=-16'd8757;
      92009:data<=-16'd8423;
      92010:data<=-16'd7959;
      92011:data<=-16'd11320;
      92012:data<=-16'd13787;
      92013:data<=-16'd13735;
      92014:data<=-16'd12222;
      92015:data<=-16'd11552;
      92016:data<=-16'd14451;
      92017:data<=-16'd9668;
      92018:data<=16'd2211;
      92019:data<=16'd3732;
      92020:data<=16'd141;
      92021:data<=16'd957;
      92022:data<=16'd1060;
      92023:data<=16'd1345;
      92024:data<=16'd1569;
      92025:data<=16'd273;
      92026:data<=16'd895;
      92027:data<=16'd1212;
      92028:data<=16'd843;
      92029:data<=16'd1030;
      92030:data<=16'd149;
      92031:data<=16'd776;
      92032:data<=16'd1105;
      92033:data<=-16'd1225;
      92034:data<=-16'd1779;
      92035:data<=-16'd1541;
      92036:data<=-16'd2094;
      92037:data<=-16'd2003;
      92038:data<=-16'd2531;
      92039:data<=-16'd2453;
      92040:data<=-16'd1903;
      92041:data<=-16'd2311;
      92042:data<=-16'd1974;
      92043:data<=-16'd1826;
      92044:data<=-16'd1762;
      92045:data<=-16'd1632;
      92046:data<=-16'd3368;
      92047:data<=-16'd3824;
      92048:data<=-16'd3049;
      92049:data<=-16'd3967;
      92050:data<=-16'd3871;
      92051:data<=-16'd3428;
      92052:data<=-16'd4034;
      92053:data<=-16'd3632;
      92054:data<=-16'd3271;
      92055:data<=-16'd3127;
      92056:data<=-16'd2751;
      92057:data<=-16'd2898;
      92058:data<=-16'd3612;
      92059:data<=-16'd4834;
      92060:data<=-16'd3835;
      92061:data<=-16'd4811;
      92062:data<=-16'd14314;
      92063:data<=-16'd20760;
      92064:data<=-16'd16387;
      92065:data<=-16'd11579;
      92066:data<=-16'd10173;
      92067:data<=-16'd9756;
      92068:data<=-16'd9591;
      92069:data<=-16'd8423;
      92070:data<=-16'd7988;
      92071:data<=-16'd7738;
      92072:data<=-16'd7420;
      92073:data<=-16'd9144;
      92074:data<=-16'd9306;
      92075:data<=-16'd7973;
      92076:data<=-16'd8481;
      92077:data<=-16'd8232;
      92078:data<=-16'd7503;
      92079:data<=-16'd7322;
      92080:data<=-16'd6147;
      92081:data<=-16'd5739;
      92082:data<=-16'd6058;
      92083:data<=-16'd5708;
      92084:data<=-16'd5286;
      92085:data<=-16'd5239;
      92086:data<=-16'd6372;
      92087:data<=-16'd7025;
      92088:data<=-16'd6222;
      92089:data<=-16'd5780;
      92090:data<=-16'd5013;
      92091:data<=-16'd4708;
      92092:data<=-16'd5460;
      92093:data<=-16'd4683;
      92094:data<=-16'd3401;
      92095:data<=-16'd2887;
      92096:data<=-16'd2845;
      92097:data<=-16'd3297;
      92098:data<=-16'd3149;
      92099:data<=-16'd4011;
      92100:data<=-16'd4773;
      92101:data<=-16'd3401;
      92102:data<=-16'd3877;
      92103:data<=-16'd3536;
      92104:data<=-16'd1588;
      92105:data<=-16'd3676;
      92106:data<=-16'd120;
      92107:data<=16'd11212;
      92108:data<=16'd14111;
      92109:data<=16'd11412;
      92110:data<=16'd12254;
      92111:data<=16'd11220;
      92112:data<=16'd9216;
      92113:data<=16'd9397;
      92114:data<=16'd8489;
      92115:data<=16'd7918;
      92116:data<=16'd8672;
      92117:data<=16'd6793;
      92118:data<=16'd2525;
      92119:data<=16'd675;
      92120:data<=16'd1663;
      92121:data<=16'd1509;
      92122:data<=16'd481;
      92123:data<=16'd699;
      92124:data<=16'd843;
      92125:data<=16'd50;
      92126:data<=-16'd1115;
      92127:data<=-16'd1447;
      92128:data<=-16'd511;
      92129:data<=-16'd202;
      92130:data<=-16'd522;
      92131:data<=-16'd317;
      92132:data<=-16'd123;
      92133:data<=-16'd77;
      92134:data<=-16'd243;
      92135:data<=-16'd250;
      92136:data<=16'd176;
      92137:data<=16'd299;
      92138:data<=-16'd29;
      92139:data<=-16'd1600;
      92140:data<=-16'd2840;
      92141:data<=-16'd1553;
      92142:data<=-16'd1290;
      92143:data<=-16'd2170;
      92144:data<=-16'd1421;
      92145:data<=-16'd1441;
      92146:data<=-16'd1048;
      92147:data<=-16'd133;
      92148:data<=-16'd1650;
      92149:data<=-16'd819;
      92150:data<=-16'd626;
      92151:data<=-16'd9250;
      92152:data<=-16'd16988;
      92153:data<=-16'd16512;
      92154:data<=-16'd15424;
      92155:data<=-16'd15299;
      92156:data<=-16'd13753;
      92157:data<=-16'd12745;
      92158:data<=-16'd12615;
      92159:data<=-16'd12507;
      92160:data<=-16'd12007;
      92161:data<=-16'd10889;
      92162:data<=-16'd10340;
      92163:data<=-16'd10734;
      92164:data<=-16'd10414;
      92165:data<=-16'd9506;
      92166:data<=-16'd9800;
      92167:data<=-16'd9521;
      92168:data<=-16'd8017;
      92169:data<=-16'd8106;
      92170:data<=-16'd6267;
      92171:data<=-16'd566;
      92172:data<=16'd1636;
      92173:data<=16'd200;
      92174:data<=16'd529;
      92175:data<=16'd1181;
      92176:data<=16'd1245;
      92177:data<=16'd1412;
      92178:data<=16'd757;
      92179:data<=16'd127;
      92180:data<=-16'd120;
      92181:data<=-16'd35;
      92182:data<=16'd502;
      92183:data<=16'd735;
      92184:data<=16'd1086;
      92185:data<=16'd951;
      92186:data<=16'd698;
      92187:data<=16'd1715;
      92188:data<=16'd1348;
      92189:data<=16'd779;
      92190:data<=16'd2150;
      92191:data<=16'd1753;
      92192:data<=16'd2278;
      92193:data<=16'd3915;
      92194:data<=16'd1401;
      92195:data<=16'd4722;
      92196:data<=16'd15957;
      92197:data<=16'd18710;
      92198:data<=16'd15571;
      92199:data<=16'd16433;
      92200:data<=16'd16301;
      92201:data<=16'd15406;
      92202:data<=16'd15913;
      92203:data<=16'd14882;
      92204:data<=16'd14957;
      92205:data<=16'd16228;
      92206:data<=16'd15769;
      92207:data<=16'd15355;
      92208:data<=16'd15188;
      92209:data<=16'd14759;
      92210:data<=16'd14571;
      92211:data<=16'd13988;
      92212:data<=16'd13706;
      92213:data<=16'd13127;
      92214:data<=16'd11684;
      92215:data<=16'd11326;
      92216:data<=16'd11339;
      92217:data<=16'd10831;
      92218:data<=16'd11262;
      92219:data<=16'd11808;
      92220:data<=16'd10930;
      92221:data<=16'd10238;
      92222:data<=16'd11135;
      92223:data<=16'd10008;
      92224:data<=16'd5580;
      92225:data<=16'd3425;
      92226:data<=16'd3688;
      92227:data<=16'd2881;
      92228:data<=16'd2654;
      92229:data<=16'd2725;
      92230:data<=16'd2554;
      92231:data<=16'd3547;
      92232:data<=16'd4206;
      92233:data<=16'd4505;
      92234:data<=16'd4329;
      92235:data<=16'd3820;
      92236:data<=16'd4689;
      92237:data<=16'd3495;
      92238:data<=16'd2379;
      92239:data<=16'd4326;
      92240:data<=-16'd1107;
      92241:data<=-16'd11109;
      92242:data<=-16'd12326;
      92243:data<=-16'd10278;
      92244:data<=-16'd9976;
      92245:data<=-16'd8249;
      92246:data<=-16'd7647;
      92247:data<=-16'd7565;
      92248:data<=-16'd6783;
      92249:data<=-16'd7063;
      92250:data<=-16'd7013;
      92251:data<=-16'd6705;
      92252:data<=-16'd6209;
      92253:data<=-16'd5471;
      92254:data<=-16'd5741;
      92255:data<=-16'd5212;
      92256:data<=-16'd4534;
      92257:data<=-16'd4548;
      92258:data<=-16'd2934;
      92259:data<=-16'd1786;
      92260:data<=-16'd1839;
      92261:data<=-16'd1431;
      92262:data<=-16'd1478;
      92263:data<=-16'd875;
      92264:data<=-16'd321;
      92265:data<=-16'd1092;
      92266:data<=-16'd1028;
      92267:data<=-16'd711;
      92268:data<=-16'd473;
      92269:data<=-16'd234;
      92270:data<=-16'd698;
      92271:data<=16'd500;
      92272:data<=16'd1999;
      92273:data<=16'd2126;
      92274:data<=16'd2619;
      92275:data<=16'd2009;
      92276:data<=16'd2711;
      92277:data<=16'd6525;
      92278:data<=16'd8508;
      92279:data<=16'd8636;
      92280:data<=16'd8258;
      92281:data<=16'd8437;
      92282:data<=16'd9427;
      92283:data<=16'd7183;
      92284:data<=16'd9632;
      92285:data<=16'd20688;
      92286:data<=16'd24521;
      92287:data<=16'd21607;
      92288:data<=16'd22089;
      92289:data<=16'd21143;
      92290:data<=16'd19581;
      92291:data<=16'd20298;
      92292:data<=16'd19420;
      92293:data<=16'd18334;
      92294:data<=16'd17752;
      92295:data<=16'd16910;
      92296:data<=16'd16333;
      92297:data<=16'd15418;
      92298:data<=16'd16078;
      92299:data<=16'd16456;
      92300:data<=16'd14578;
      92301:data<=16'd14257;
      92302:data<=16'd14160;
      92303:data<=16'd13036;
      92304:data<=16'd12713;
      92305:data<=16'd11649;
      92306:data<=16'd11121;
      92307:data<=16'd11091;
      92308:data<=16'd9659;
      92309:data<=16'd9145;
      92310:data<=16'd9115;
      92311:data<=16'd9502;
      92312:data<=16'd10464;
      92313:data<=16'd9174;
      92314:data<=16'd8542;
      92315:data<=16'd8815;
      92316:data<=16'd6872;
      92317:data<=16'd6134;
      92318:data<=16'd6084;
      92319:data<=16'd5468;
      92320:data<=16'd6053;
      92321:data<=16'd5325;
      92322:data<=16'd4743;
      92323:data<=16'd4528;
      92324:data<=16'd3080;
      92325:data<=16'd4915;
      92326:data<=16'd5147;
      92327:data<=16'd2379;
      92328:data<=16'd4733;
      92329:data<=16'd529;
      92330:data<=-16'd14131;
      92331:data<=-16'd19864;
      92332:data<=-16'd17747;
      92333:data<=-16'd18237;
      92334:data<=-16'd17895;
      92335:data<=-16'd17327;
      92336:data<=-16'd17623;
      92337:data<=-16'd16199;
      92338:data<=-16'd14727;
      92339:data<=-16'd13932;
      92340:data<=-16'd13717;
      92341:data<=-16'd13711;
      92342:data<=-16'd12742;
      92343:data<=-16'd12298;
      92344:data<=-16'd12348;
      92345:data<=-16'd12005;
      92346:data<=-16'd11960;
      92347:data<=-16'd11356;
      92348:data<=-16'd10531;
      92349:data<=-16'd10217;
      92350:data<=-16'd9403;
      92351:data<=-16'd8378;
      92352:data<=-16'd7456;
      92353:data<=-16'd6912;
      92354:data<=-16'd7060;
      92355:data<=-16'd6899;
      92356:data<=-16'd6789;
      92357:data<=-16'd6966;
      92358:data<=-16'd6590;
      92359:data<=-16'd6352;
      92360:data<=-16'd6373;
      92361:data<=-16'd6015;
      92362:data<=-16'd5506;
      92363:data<=-16'd5404;
      92364:data<=-16'd5362;
      92365:data<=-16'd4018;
      92366:data<=-16'd3025;
      92367:data<=-16'd3550;
      92368:data<=-16'd3005;
      92369:data<=-16'd2728;
      92370:data<=-16'd3090;
      92371:data<=-16'd1968;
      92372:data<=-16'd2942;
      92373:data<=-16'd2071;
      92374:data<=16'd7072;
      92375:data<=16'd13388;
      92376:data<=16'd11632;
      92377:data<=16'd11843;
      92378:data<=16'd13385;
      92379:data<=16'd12072;
      92380:data<=16'd11925;
      92381:data<=16'd12254;
      92382:data<=16'd11054;
      92383:data<=16'd12422;
      92384:data<=16'd15898;
      92385:data<=16'd16089;
      92386:data<=16'd14668;
      92387:data<=16'd15114;
      92388:data<=16'd14334;
      92389:data<=16'd12602;
      92390:data<=16'd13062;
      92391:data<=16'd13330;
      92392:data<=16'd12889;
      92393:data<=16'd12692;
      92394:data<=16'd11464;
      92395:data<=16'd10972;
      92396:data<=16'd10881;
      92397:data<=16'd9568;
      92398:data<=16'd9280;
      92399:data<=16'd9077;
      92400:data<=16'd8172;
      92401:data<=16'd8081;
      92402:data<=16'd7040;
      92403:data<=16'd5724;
      92404:data<=16'd5479;
      92405:data<=16'd4968;
      92406:data<=16'd4866;
      92407:data<=16'd4592;
      92408:data<=16'd4196;
      92409:data<=16'd4578;
      92410:data<=16'd3568;
      92411:data<=16'd2781;
      92412:data<=16'd2855;
      92413:data<=16'd1700;
      92414:data<=16'd2050;
      92415:data<=16'd1888;
      92416:data<=16'd331;
      92417:data<=16'd1190;
      92418:data<=-16'd3883;
      92419:data<=-16'd14828;
      92420:data<=-16'd17429;
      92421:data<=-16'd15644;
      92422:data<=-16'd16848;
      92423:data<=-16'd16424;
      92424:data<=-16'd15837;
      92425:data<=-16'd16043;
      92426:data<=-16'd14819;
      92427:data<=-16'd14862;
      92428:data<=-16'd15024;
      92429:data<=-16'd13658;
      92430:data<=-16'd13843;
      92431:data<=-16'd15273;
      92432:data<=-16'd15437;
      92433:data<=-16'd14678;
      92434:data<=-16'd14179;
      92435:data<=-16'd13570;
      92436:data<=-16'd14404;
      92437:data<=-16'd18172;
      92438:data<=-16'd19646;
      92439:data<=-16'd17711;
      92440:data<=-16'd17666;
      92441:data<=-16'd17584;
      92442:data<=-16'd16146;
      92443:data<=-16'd16277;
      92444:data<=-16'd16498;
      92445:data<=-16'd16688;
      92446:data<=-16'd16725;
      92447:data<=-16'd15335;
      92448:data<=-16'd14939;
      92449:data<=-16'd14672;
      92450:data<=-16'd13747;
      92451:data<=-16'd13914;
      92452:data<=-16'd13207;
      92453:data<=-16'd12595;
      92454:data<=-16'd12492;
      92455:data<=-16'd10704;
      92456:data<=-16'd10681;
      92457:data<=-16'd11653;
      92458:data<=-16'd10909;
      92459:data<=-16'd10798;
      92460:data<=-16'd9559;
      92461:data<=-16'd9156;
      92462:data<=-16'd10185;
      92463:data<=-16'd3280;
      92464:data<=16'd6149;
      92465:data<=16'd7095;
      92466:data<=16'd5911;
      92467:data<=16'd6404;
      92468:data<=16'd6256;
      92469:data<=16'd6534;
      92470:data<=16'd5485;
      92471:data<=16'd3964;
      92472:data<=16'd4425;
      92473:data<=16'd4232;
      92474:data<=16'd3345;
      92475:data<=16'd3648;
      92476:data<=16'd3985;
      92477:data<=16'd3660;
      92478:data<=16'd3471;
      92479:data<=16'd3491;
      92480:data<=16'd3051;
      92481:data<=16'd3130;
      92482:data<=16'd3704;
      92483:data<=16'd2772;
      92484:data<=16'd1607;
      92485:data<=16'd1271;
      92486:data<=16'd1071;
      92487:data<=16'd1237;
      92488:data<=16'd549;
      92489:data<=16'd1582;
      92490:data<=16'd6046;
      92491:data<=16'd7460;
      92492:data<=16'd6343;
      92493:data<=16'd7177;
      92494:data<=16'd7065;
      92495:data<=16'd6545;
      92496:data<=16'd6457;
      92497:data<=16'd4902;
      92498:data<=16'd4206;
      92499:data<=16'd3970;
      92500:data<=16'd3409;
      92501:data<=16'd3717;
      92502:data<=16'd3418;
      92503:data<=16'd3541;
      92504:data<=16'd2713;
      92505:data<=16'd1137;
      92506:data<=16'd3680;
      92507:data<=16'd1193;
      92508:data<=-16'd9659;
      92509:data<=-16'd13755;
      92510:data<=-16'd12777;
      92511:data<=-16'd14595;
      92512:data<=-16'd13922;
      92513:data<=-16'd12569;
      92514:data<=-16'd12963;
      92515:data<=-16'd12010;
      92516:data<=-16'd11455;
      92517:data<=-16'd11207;
      92518:data<=-16'd10751;
      92519:data<=-16'd10527;
      92520:data<=-16'd9280;
      92521:data<=-16'd8989;
      92522:data<=-16'd8896;
      92523:data<=-16'd8232;
      92524:data<=-16'd9734;
      92525:data<=-16'd10058;
      92526:data<=-16'd8599;
      92527:data<=-16'd8827;
      92528:data<=-16'd8457;
      92529:data<=-16'd7583;
      92530:data<=-16'd7298;
      92531:data<=-16'd6570;
      92532:data<=-16'd6408;
      92533:data<=-16'd5677;
      92534:data<=-16'd4965;
      92535:data<=-16'd5310;
      92536:data<=-16'd4896;
      92537:data<=-16'd5905;
      92538:data<=-16'd6968;
      92539:data<=-16'd5805;
      92540:data<=-16'd5897;
      92541:data<=-16'd5347;
      92542:data<=-16'd5674;
      92543:data<=-16'd10110;
      92544:data<=-16'd11264;
      92545:data<=-16'd9908;
      92546:data<=-16'd10331;
      92547:data<=-16'd9365;
      92548:data<=-16'd9154;
      92549:data<=-16'd8332;
      92550:data<=-16'd7247;
      92551:data<=-16'd10584;
      92552:data<=-16'd6338;
      92553:data<=16'd6028;
      92554:data<=16'd8957;
      92555:data<=16'd6898;
      92556:data<=16'd7915;
      92557:data<=16'd7423;
      92558:data<=16'd7253;
      92559:data<=16'd7497;
      92560:data<=16'd6878;
      92561:data<=16'd7724;
      92562:data<=16'd7453;
      92563:data<=16'd6120;
      92564:data<=16'd5368;
      92565:data<=16'd4176;
      92566:data<=16'd4555;
      92567:data<=16'd5304;
      92568:data<=16'd4714;
      92569:data<=16'd4878;
      92570:data<=16'd4493;
      92571:data<=16'd3967;
      92572:data<=16'd5072;
      92573:data<=16'd5371;
      92574:data<=16'd4837;
      92575:data<=16'd4590;
      92576:data<=16'd3554;
      92577:data<=16'd2255;
      92578:data<=16'd1898;
      92579:data<=16'd2361;
      92580:data<=16'd2588;
      92581:data<=16'd2801;
      92582:data<=16'd3354;
      92583:data<=16'd2907;
      92584:data<=16'd2584;
      92585:data<=16'd3157;
      92586:data<=16'd2958;
      92587:data<=16'd2766;
      92588:data<=16'd2529;
      92589:data<=16'd1827;
      92590:data<=16'd1530;
      92591:data<=16'd693;
      92592:data<=16'd861;
      92593:data<=16'd1283;
      92594:data<=-16'd332;
      92595:data<=16'd1845;
      92596:data<=16'd4323;
      92597:data<=-16'd2229;
      92598:data<=-16'd8078;
      92599:data<=-16'd6783;
      92600:data<=-16'd6347;
      92601:data<=-16'd6200;
      92602:data<=-16'd4686;
      92603:data<=-16'd5388;
      92604:data<=-16'd6737;
      92605:data<=-16'd7250;
      92606:data<=-16'd7250;
      92607:data<=-16'd6498;
      92608:data<=-16'd5761;
      92609:data<=-16'd4846;
      92610:data<=-16'd4469;
      92611:data<=-16'd4843;
      92612:data<=-16'd4196;
      92613:data<=-16'd3547;
      92614:data<=-16'd3570;
      92615:data<=-16'd3209;
      92616:data<=-16'd2892;
      92617:data<=-16'd2549;
      92618:data<=-16'd2522;
      92619:data<=-16'd2787;
      92620:data<=-16'd2067;
      92621:data<=-16'd1401;
      92622:data<=-16'd1154;
      92623:data<=-16'd575;
      92624:data<=-16'd561;
      92625:data<=-16'd596;
      92626:data<=-16'd92;
      92627:data<=16'd92;
      92628:data<=-16'd33;
      92629:data<=16'd384;
      92630:data<=16'd1985;
      92631:data<=16'd2651;
      92632:data<=16'd1938;
      92633:data<=16'd2705;
      92634:data<=16'd3008;
      92635:data<=16'd2393;
      92636:data<=16'd3294;
      92637:data<=16'd2998;
      92638:data<=16'd3292;
      92639:data<=16'd4657;
      92640:data<=16'd2341;
      92641:data<=16'd5615;
      92642:data<=16'd16809;
      92643:data<=16'd20183;
      92644:data<=16'd18207;
      92645:data<=16'd19699;
      92646:data<=16'd18842;
      92647:data<=16'd17264;
      92648:data<=16'd17487;
      92649:data<=16'd14076;
      92650:data<=16'd10229;
      92651:data<=16'd9777;
      92652:data<=16'd9547;
      92653:data<=16'd8583;
      92654:data<=16'd7577;
      92655:data<=16'd7621;
      92656:data<=16'd9179;
      92657:data<=16'd10117;
      92658:data<=16'd9714;
      92659:data<=16'd9197;
      92660:data<=16'd8966;
      92661:data<=16'd8496;
      92662:data<=16'd8061;
      92663:data<=16'd8222;
      92664:data<=16'd7899;
      92665:data<=16'd7260;
      92666:data<=16'd6842;
      92667:data<=16'd5483;
      92668:data<=16'd5166;
      92669:data<=16'd7191;
      92670:data<=16'd8172;
      92671:data<=16'd7571;
      92672:data<=16'd7477;
      92673:data<=16'd7718;
      92674:data<=16'd7262;
      92675:data<=16'd6387;
      92676:data<=16'd6225;
      92677:data<=16'd5977;
      92678:data<=16'd5412;
      92679:data<=16'd5582;
      92680:data<=16'd4960;
      92681:data<=16'd4493;
      92682:data<=16'd5418;
      92683:data<=16'd5310;
      92684:data<=16'd6172;
      92685:data<=16'd6026;
      92686:data<=-16'd1668;
      92687:data<=-16'd9238;
      92688:data<=-16'd9407;
      92689:data<=-16'd8733;
      92690:data<=-16'd9235;
      92691:data<=-16'd8715;
      92692:data<=-16'd8385;
      92693:data<=-16'd8153;
      92694:data<=-16'd8251;
      92695:data<=-16'd7968;
      92696:data<=-16'd6056;
      92697:data<=-16'd5062;
      92698:data<=-16'd5142;
      92699:data<=-16'd3956;
      92700:data<=-16'd3413;
      92701:data<=-16'd4501;
      92702:data<=-16'd2911;
      92703:data<=16'd1841;
      92704:data<=16'd3786;
      92705:data<=16'd2643;
      92706:data<=16'd2641;
      92707:data<=16'd2560;
      92708:data<=16'd2141;
      92709:data<=16'd3092;
      92710:data<=16'd3758;
      92711:data<=16'd4112;
      92712:data<=16'd4255;
      92713:data<=16'd3779;
      92714:data<=16'd3970;
      92715:data<=16'd3165;
      92716:data<=16'd2044;
      92717:data<=16'd2852;
      92718:data<=16'd2831;
      92719:data<=16'd2719;
      92720:data<=16'd3190;
      92721:data<=16'd1888;
      92722:data<=16'd2200;
      92723:data<=16'd3988;
      92724:data<=16'd4206;
      92725:data<=16'd4579;
      92726:data<=16'd4068;
      92727:data<=16'd4249;
      92728:data<=16'd5536;
      92729:data<=16'd3292;
      92730:data<=16'd5797;
      92731:data<=16'd15803;
      92732:data<=16'd19023;
      92733:data<=16'd16600;
      92734:data<=16'd16636;
      92735:data<=16'd16263;
      92736:data<=16'd16310;
      92737:data<=16'd16804;
      92738:data<=16'd15459;
      92739:data<=16'd14854;
      92740:data<=16'd14134;
      92741:data<=16'd12881;
      92742:data<=16'd12953;
      92743:data<=16'd12172;
      92744:data<=16'd10978;
      92745:data<=16'd10977;
      92746:data<=16'd10680;
      92747:data<=16'd10056;
      92748:data<=16'd9426;
      92749:data<=16'd8810;
      92750:data<=16'd8758;
      92751:data<=16'd9169;
      92752:data<=16'd9042;
      92753:data<=16'd7738;
      92754:data<=16'd7203;
      92755:data<=16'd5752;
      92756:data<=16'd811;
      92757:data<=-16'd1486;
      92758:data<=-16'd525;
      92759:data<=-16'd1706;
      92760:data<=-16'd1680;
      92761:data<=-16'd682;
      92762:data<=-16'd1480;
      92763:data<=-16'd238;
      92764:data<=16'd870;
      92765:data<=-16'd41;
      92766:data<=16'd112;
      92767:data<=-16'd387;
      92768:data<=-16'd879;
      92769:data<=-16'd514;
      92770:data<=-16'd1183;
      92771:data<=-16'd1111;
      92772:data<=-16'd2026;
      92773:data<=-16'd3113;
      92774:data<=-16'd1494;
      92775:data<=-16'd5724;
      92776:data<=-16'd14618;
      92777:data<=-16'd16216;
      92778:data<=-16'd14568;
      92779:data<=-16'd15121;
      92780:data<=-16'd14659;
      92781:data<=-16'd14264;
      92782:data<=-16'd14146;
      92783:data<=-16'd13488;
      92784:data<=-16'd13549;
      92785:data<=-16'd12960;
      92786:data<=-16'd12236;
      92787:data<=-16'd12463;
      92788:data<=-16'd11529;
      92789:data<=-16'd9893;
      92790:data<=-16'd9204;
      92791:data<=-16'd8799;
      92792:data<=-16'd8413;
      92793:data<=-16'd8214;
      92794:data<=-16'd7758;
      92795:data<=-16'd7445;
      92796:data<=-16'd7876;
      92797:data<=-16'd7999;
      92798:data<=-16'd7591;
      92799:data<=-16'd7362;
      92800:data<=-16'd6810;
      92801:data<=-16'd6579;
      92802:data<=-16'd6072;
      92803:data<=-16'd4349;
      92804:data<=-16'd4485;
      92805:data<=-16'd5143;
      92806:data<=-16'd3987;
      92807:data<=-16'd4300;
      92808:data<=-16'd3027;
      92809:data<=16'd1391;
      92810:data<=16'd2529;
      92811:data<=16'd2123;
      92812:data<=16'd2587;
      92813:data<=16'd1897;
      92814:data<=16'd2243;
      92815:data<=16'd2698;
      92816:data<=16'd3354;
      92817:data<=16'd4849;
      92818:data<=16'd2707;
      92819:data<=16'd4391;
      92820:data<=16'd14477;
      92821:data<=16'd18965;
      92822:data<=16'd16396;
      92823:data<=16'd15493;
      92824:data<=16'd15059;
      92825:data<=16'd14694;
      92826:data<=16'd14084;
      92827:data<=16'd12361;
      92828:data<=16'd11958;
      92829:data<=16'd11503;
      92830:data<=16'd10988;
      92831:data<=16'd11370;
      92832:data<=16'd10182;
      92833:data<=16'd9226;
      92834:data<=16'd9464;
      92835:data<=16'd8912;
      92836:data<=16'd8475;
      92837:data<=16'd7750;
      92838:data<=16'd6939;
      92839:data<=16'd6827;
      92840:data<=16'd6140;
      92841:data<=16'd5506;
      92842:data<=16'd4420;
      92843:data<=16'd3143;
      92844:data<=16'd3265;
      92845:data<=16'd2284;
      92846:data<=16'd1307;
      92847:data<=16'd1985;
      92848:data<=16'd1386;
      92849:data<=16'd1021;
      92850:data<=16'd1089;
      92851:data<=16'd402;
      92852:data<=16'd1061;
      92853:data<=16'd576;
      92854:data<=-16'd787;
      92855:data<=-16'd1216;
      92856:data<=-16'd3127;
      92857:data<=-16'd2734;
      92858:data<=-16'd1536;
      92859:data<=-16'd3627;
      92860:data<=-16'd2813;
      92861:data<=-16'd3877;
      92862:data<=-16'd9036;
      92863:data<=-16'd8126;
      92864:data<=-16'd11517;
      92865:data<=-16'd23353;
      92866:data<=-16'd25560;
      92867:data<=-16'd21816;
      92868:data<=-16'd22991;
      92869:data<=-16'd23728;
      92870:data<=-16'd22949;
      92871:data<=-16'd21849;
      92872:data<=-16'd20421;
      92873:data<=-16'd20592;
      92874:data<=-16'd20357;
      92875:data<=-16'd19456;
      92876:data<=-16'd18578;
      92877:data<=-16'd17241;
      92878:data<=-16'd17429;
      92879:data<=-16'd17153;
      92880:data<=-16'd15531;
      92881:data<=-16'd15945;
      92882:data<=-16'd16422;
      92883:data<=-16'd15687;
      92884:data<=-16'd15675;
      92885:data<=-16'd15520;
      92886:data<=-16'd14912;
      92887:data<=-16'd14025;
      92888:data<=-16'd13094;
      92889:data<=-16'd12762;
      92890:data<=-16'd12010;
      92891:data<=-16'd11085;
      92892:data<=-16'd10528;
      92893:data<=-16'd9941;
      92894:data<=-16'd9871;
      92895:data<=-16'd10052;
      92896:data<=-16'd10514;
      92897:data<=-16'd10489;
      92898:data<=-16'd9230;
      92899:data<=-16'd9139;
      92900:data<=-16'd9165;
      92901:data<=-16'd8190;
      92902:data<=-16'd8537;
      92903:data<=-16'd7840;
      92904:data<=-16'd6525;
      92905:data<=-16'd6849;
      92906:data<=-16'd5753;
      92907:data<=-16'd5970;
      92908:data<=-16'd5902;
      92909:data<=16'd1959;
      92910:data<=16'd8884;
      92911:data<=16'd8572;
      92912:data<=16'd8341;
      92913:data<=16'd7955;
      92914:data<=16'd7787;
      92915:data<=16'd11344;
      92916:data<=16'd13715;
      92917:data<=16'd13160;
      92918:data<=16'd12598;
      92919:data<=16'd12443;
      92920:data<=16'd12789;
      92921:data<=16'd11843;
      92922:data<=16'd9738;
      92923:data<=16'd9289;
      92924:data<=16'd9664;
      92925:data<=16'd9320;
      92926:data<=16'd8436;
      92927:data<=16'd7773;
      92928:data<=16'd7685;
      92929:data<=16'd7341;
      92930:data<=16'd7265;
      92931:data<=16'd7185;
      92932:data<=16'd6448;
      92933:data<=16'd6525;
      92934:data<=16'd6087;
      92935:data<=16'd4520;
      92936:data<=16'd3988;
      92937:data<=16'd3613;
      92938:data<=16'd3482;
      92939:data<=16'd3755;
      92940:data<=16'd2966;
      92941:data<=16'd2921;
      92942:data<=16'd3460;
      92943:data<=16'd3275;
      92944:data<=16'd3101;
      92945:data<=16'd2040;
      92946:data<=16'd2046;
      92947:data<=16'd3095;
      92948:data<=16'd1835;
      92949:data<=16'd1118;
      92950:data<=16'd423;
      92951:data<=-16'd745;
      92952:data<=16'd1823;
      92953:data<=-16'd917;
      92954:data<=-16'd11506;
      92955:data<=-16'd14909;
      92956:data<=-16'd12511;
      92957:data<=-16'd12790;
      92958:data<=-16'd12295;
      92959:data<=-16'd11335;
      92960:data<=-16'd10972;
      92961:data<=-16'd10329;
      92962:data<=-16'd11217;
      92963:data<=-16'd11285;
      92964:data<=-16'd10433;
      92965:data<=-16'd10624;
      92966:data<=-16'd9238;
      92967:data<=-16'd8590;
      92968:data<=-16'd11721;
      92969:data<=-16'd14475;
      92970:data<=-16'd14242;
      92971:data<=-16'd12496;
      92972:data<=-16'd11338;
      92973:data<=-16'd11332;
      92974:data<=-16'd11815;
      92975:data<=-16'd12525;
      92976:data<=-16'd12000;
      92977:data<=-16'd10851;
      92978:data<=-16'd10684;
      92979:data<=-16'd9703;
      92980:data<=-16'd8907;
      92981:data<=-16'd9317;
      92982:data<=-16'd8210;
      92983:data<=-16'd6984;
      92984:data<=-16'd6880;
      92985:data<=-16'd6002;
      92986:data<=-16'd5234;
      92987:data<=-16'd5354;
      92988:data<=-16'd5924;
      92989:data<=-16'd5968;
      92990:data<=-16'd5150;
      92991:data<=-16'd5483;
      92992:data<=-16'd5272;
      92993:data<=-16'd3767;
      92994:data<=-16'd3896;
      92995:data<=-16'd3102;
      92996:data<=-16'd2276;
      92997:data<=-16'd3203;
      92998:data<=16'd2716;
      92999:data<=16'd12496;
      93000:data<=16'd13954;
      93001:data<=16'd11424;
      93002:data<=16'd10957;
      93003:data<=16'd10328;
      93004:data<=16'd10060;
      93005:data<=16'd9718;
      93006:data<=16'd9130;
      93007:data<=16'd9776;
      93008:data<=16'd9650;
      93009:data<=16'd9147;
      93010:data<=16'd9592;
      93011:data<=16'd8925;
      93012:data<=16'd8534;
      93013:data<=16'd9653;
      93014:data<=16'd9380;
      93015:data<=16'd7835;
      93016:data<=16'd6408;
      93017:data<=16'd5084;
      93018:data<=16'd5600;
      93019:data<=16'd6572;
      93020:data<=16'd5520;
      93021:data<=16'd6972;
      93022:data<=16'd11439;
      93023:data<=16'd12132;
      93024:data<=16'd10812;
      93025:data<=16'd11502;
      93026:data<=16'd11159;
      93027:data<=16'd10276;
      93028:data<=16'd9882;
      93029:data<=16'd8137;
      93030:data<=16'd7344;
      93031:data<=16'd7608;
      93032:data<=16'd6960;
      93033:data<=16'd6670;
      93034:data<=16'd6172;
      93035:data<=16'd6018;
      93036:data<=16'd7001;
      93037:data<=16'd6865;
      93038:data<=16'd6546;
      93039:data<=16'd5702;
      93040:data<=16'd4440;
      93041:data<=16'd6091;
      93042:data<=16'd3532;
      93043:data<=-16'd6313;
      93044:data<=-16'd10904;
      93045:data<=-16'd9253;
      93046:data<=-16'd9342;
      93047:data<=-16'd9576;
      93048:data<=-16'd8795;
      93049:data<=-16'd8055;
      93050:data<=-16'd7036;
      93051:data<=-16'd6784;
      93052:data<=-16'd6684;
      93053:data<=-16'd6381;
      93054:data<=-16'd5488;
      93055:data<=-16'd3227;
      93056:data<=-16'd2858;
      93057:data<=-16'd4097;
      93058:data<=-16'd3316;
      93059:data<=-16'd2749;
      93060:data<=-16'd3265;
      93061:data<=-16'd2323;
      93062:data<=-16'd1418;
      93063:data<=-16'd2062;
      93064:data<=-16'd2147;
      93065:data<=-16'd1143;
      93066:data<=-16'd1172;
      93067:data<=-16'd1055;
      93068:data<=16'd1033;
      93069:data<=16'd2003;
      93070:data<=16'd1431;
      93071:data<=16'd1387;
      93072:data<=16'd1137;
      93073:data<=16'd1648;
      93074:data<=16'd890;
      93075:data<=-16'd3095;
      93076:data<=-16'd4313;
      93077:data<=-16'd3236;
      93078:data<=-16'd3814;
      93079:data<=-16'd3021;
      93080:data<=-16'd2408;
      93081:data<=-16'd2293;
      93082:data<=-16'd194;
      93083:data<=-16'd247;
      93084:data<=-16'd352;
      93085:data<=16'd749;
      93086:data<=-16'd1413;
      93087:data<=16'd2499;
      93088:data<=16'd13591;
      93089:data<=16'd16181;
      93090:data<=16'd13069;
      93091:data<=16'd13805;
      93092:data<=16'd14273;
      93093:data<=16'd13658;
      93094:data<=16'd14189;
      93095:data<=16'd14480;
      93096:data<=16'd14304;
      93097:data<=16'd13734;
      93098:data<=16'd13358;
      93099:data<=16'd13024;
      93100:data<=16'd12055;
      93101:data<=16'd11943;
      93102:data<=16'd11941;
      93103:data<=16'd10985;
      93104:data<=16'd10812;
      93105:data<=16'd10680;
      93106:data<=16'd9644;
      93107:data<=16'd9459;
      93108:data<=16'd10154;
      93109:data<=16'd10381;
      93110:data<=16'd10248;
      93111:data<=16'd9938;
      93112:data<=16'd8872;
      93113:data<=16'd8025;
      93114:data<=16'd8254;
      93115:data<=16'd8062;
      93116:data<=16'd7797;
      93117:data<=16'd7835;
      93118:data<=16'd6677;
      93119:data<=16'd6005;
      93120:data<=16'd6599;
      93121:data<=16'd7092;
      93122:data<=16'd7685;
      93123:data<=16'd6942;
      93124:data<=16'd6126;
      93125:data<=16'd6645;
      93126:data<=16'd5379;
      93127:data<=16'd6320;
      93128:data<=16'd10525;
      93129:data<=16'd10815;
      93130:data<=16'd10774;
      93131:data<=16'd9367;
      93132:data<=-16'd444;
      93133:data<=-16'd6616;
      93134:data<=-16'd3814;
      93135:data<=-16'd3319;
      93136:data<=-16'd4360;
      93137:data<=-16'd3917;
      93138:data<=-16'd4118;
      93139:data<=-16'd3418;
      93140:data<=-16'd3334;
      93141:data<=-16'd3859;
      93142:data<=-16'd3253;
      93143:data<=-16'd3592;
      93144:data<=-16'd3451;
      93145:data<=-16'd2964;
      93146:data<=-16'd3832;
      93147:data<=-16'd2830;
      93148:data<=-16'd1225;
      93149:data<=-16'd1339;
      93150:data<=-16'd867;
      93151:data<=-16'd446;
      93152:data<=-16'd886;
      93153:data<=-16'd1219;
      93154:data<=-16'd1248;
      93155:data<=-16'd1048;
      93156:data<=-16'd1287;
      93157:data<=-16'd834;
      93158:data<=-16'd397;
      93159:data<=-16'd1651;
      93160:data<=-16'd1033;
      93161:data<=16'd954;
      93162:data<=16'd1039;
      93163:data<=16'd1163;
      93164:data<=16'd1001;
      93165:data<=16'd399;
      93166:data<=16'd664;
      93167:data<=16'd356;
      93168:data<=16'd341;
      93169:data<=16'd100;
      93170:data<=-16'd523;
      93171:data<=16'd550;
      93172:data<=16'd42;
      93173:data<=16'd30;
      93174:data<=16'd2361;
      93175:data<=16'd1002;
      93176:data<=16'd3930;
      93177:data<=16'd14322;
      93178:data<=16'd17344;
      93179:data<=16'd15092;
      93180:data<=16'd14001;
      93181:data<=16'd9392;
      93182:data<=16'd6579;
      93183:data<=16'd7356;
      93184:data<=16'd6135;
      93185:data<=16'd5479;
      93186:data<=16'd5779;
      93187:data<=16'd6213;
      93188:data<=16'd7345;
      93189:data<=16'd6346;
      93190:data<=16'd5536;
      93191:data<=16'd6223;
      93192:data<=16'd5198;
      93193:data<=16'd4620;
      93194:data<=16'd5018;
      93195:data<=16'd4200;
      93196:data<=16'd3421;
      93197:data<=16'd3102;
      93198:data<=16'd2911;
      93199:data<=16'd2654;
      93200:data<=16'd2695;
      93201:data<=16'd3902;
      93202:data<=16'd4191;
      93203:data<=16'd3052;
      93204:data<=16'd2444;
      93205:data<=16'd2366;
      93206:data<=16'd2752;
      93207:data<=16'd2723;
      93208:data<=16'd1856;
      93209:data<=16'd1401;
      93210:data<=16'd949;
      93211:data<=16'd688;
      93212:data<=16'd318;
      93213:data<=-16'd246;
      93214:data<=16'd1213;
      93215:data<=16'd1915;
      93216:data<=16'd705;
      93217:data<=16'd1165;
      93218:data<=16'd801;
      93219:data<=16'd170;
      93220:data<=16'd171;
      93221:data<=-16'd6716;
      93222:data<=-16'd15289;
      93223:data<=-16'd15738;
      93224:data<=-16'd14689;
      93225:data<=-16'd15368;
      93226:data<=-16'd13790;
      93227:data<=-16'd12052;
      93228:data<=-16'd11543;
      93229:data<=-16'd11342;
      93230:data<=-16'd10645;
      93231:data<=-16'd9521;
      93232:data<=-16'd10025;
      93233:data<=-16'd9474;
      93234:data<=-16'd5624;
      93235:data<=-16'd3353;
      93236:data<=-16'd3838;
      93237:data<=-16'd3936;
      93238:data<=-16'd3747;
      93239:data<=-16'd3545;
      93240:data<=-16'd2325;
      93241:data<=-16'd930;
      93242:data<=-16'd923;
      93243:data<=-16'd1319;
      93244:data<=-16'd1090;
      93245:data<=-16'd1184;
      93246:data<=-16'd1284;
      93247:data<=-16'd1579;
      93248:data<=-16'd2250;
      93249:data<=-16'd1610;
      93250:data<=-16'd1422;
      93251:data<=-16'd2544;
      93252:data<=-16'd2261;
      93253:data<=-16'd1820;
      93254:data<=-16'd2073;
      93255:data<=-16'd1906;
      93256:data<=-16'd2073;
      93257:data<=-16'd2067;
      93258:data<=-16'd2379;
      93259:data<=-16'd2413;
      93260:data<=-16'd1207;
      93261:data<=-16'd2494;
      93262:data<=-16'd3483;
      93263:data<=-16'd2012;
      93264:data<=-16'd3410;
      93265:data<=-16'd227;
      93266:data<=16'd9894;
      93267:data<=16'd12222;
      93268:data<=16'd9085;
      93269:data<=16'd9395;
      93270:data<=16'd8833;
      93271:data<=16'd8043;
      93272:data<=16'd8158;
      93273:data<=16'd6928;
      93274:data<=16'd6714;
      93275:data<=16'd6131;
      93276:data<=16'd4617;
      93277:data<=16'd4805;
      93278:data<=16'd4683;
      93279:data<=16'd4202;
      93280:data<=16'd3818;
      93281:data<=16'd2165;
      93282:data<=16'd1586;
      93283:data<=16'd1964;
      93284:data<=16'd1356;
      93285:data<=16'd1008;
      93286:data<=16'd473;
      93287:data<=-16'd1885;
      93288:data<=-16'd5227;
      93289:data<=-16'd6601;
      93290:data<=-16'd5761;
      93291:data<=-16'd5750;
      93292:data<=-16'd5937;
      93293:data<=-16'd6167;
      93294:data<=-16'd7805;
      93295:data<=-16'd7743;
      93296:data<=-16'd6730;
      93297:data<=-16'd7350;
      93298:data<=-16'd7192;
      93299:data<=-16'd7062;
      93300:data<=-16'd7518;
      93301:data<=-16'd7147;
      93302:data<=-16'd7509;
      93303:data<=-16'd7118;
      93304:data<=-16'd6011;
      93305:data<=-16'd6467;
      93306:data<=-16'd6711;
      93307:data<=-16'd8178;
      93308:data<=-16'd8947;
      93309:data<=-16'd6149;
      93310:data<=-16'd10390;
      93311:data<=-16'd21156;
      93312:data<=-16'd23576;
      93313:data<=-16'd20685;
      93314:data<=-16'd20434;
      93315:data<=-16'd19837;
      93316:data<=-16'd19197;
      93317:data<=-16'd18891;
      93318:data<=-16'd17252;
      93319:data<=-16'd16866;
      93320:data<=-16'd17672;
      93321:data<=-16'd17177;
      93322:data<=-16'd16134;
      93323:data<=-16'd15749;
      93324:data<=-16'd15935;
      93325:data<=-16'd15753;
      93326:data<=-16'd14698;
      93327:data<=-16'd13493;
      93328:data<=-16'd12443;
      93329:data<=-16'd11731;
      93330:data<=-16'd11491;
      93331:data<=-16'd10962;
      93332:data<=-16'd10530;
      93333:data<=-16'd11320;
      93334:data<=-16'd11747;
      93335:data<=-16'd10754;
      93336:data<=-16'd10643;
      93337:data<=-16'd10774;
      93338:data<=-16'd9212;
      93339:data<=-16'd7785;
      93340:data<=-16'd5262;
      93341:data<=-16'd1149;
      93342:data<=-16'd558;
      93343:data<=-16'd1626;
      93344:data<=-16'd325;
      93345:data<=-16'd82;
      93346:data<=-16'd1137;
      93347:data<=-16'd1697;
      93348:data<=-16'd2130;
      93349:data<=-16'd1515;
      93350:data<=-16'd1434;
      93351:data<=-16'd1240;
      93352:data<=-16'd102;
      93353:data<=-16'd1868;
      93354:data<=16'd305;
      93355:data<=16'd10834;
      93356:data<=16'd16186;
      93357:data<=16'd14377;
      93358:data<=16'd14449;
      93359:data<=16'd13899;
      93360:data<=16'd11603;
      93361:data<=16'd10746;
      93362:data<=16'd10428;
      93363:data<=16'd10063;
      93364:data<=16'd8942;
      93365:data<=16'd7964;
      93366:data<=16'd8381;
      93367:data<=16'd8257;
      93368:data<=16'd8278;
      93369:data<=16'd8722;
      93370:data<=16'd8260;
      93371:data<=16'd8216;
      93372:data<=16'd7292;
      93373:data<=16'd5160;
      93374:data<=16'd4513;
      93375:data<=16'd4212;
      93376:data<=16'd3788;
      93377:data<=16'd3936;
      93378:data<=16'd3720;
      93379:data<=16'd3570;
      93380:data<=16'd3422;
      93381:data<=16'd3720;
      93382:data<=16'd4408;
      93383:data<=16'd3707;
      93384:data<=16'd3450;
      93385:data<=16'd3718;
      93386:data<=16'd2504;
      93387:data<=16'd1635;
      93388:data<=16'd1121;
      93389:data<=16'd1105;
      93390:data<=16'd1703;
      93391:data<=16'd849;
      93392:data<=16'd1162;
      93393:data<=16'd720;
      93394:data<=-16'd3206;
      93395:data<=-16'd3653;
      93396:data<=-16'd2899;
      93397:data<=-16'd3673;
      93398:data<=-16'd591;
      93399:data<=-16'd4290;
      93400:data<=-16'd17155;
      93401:data<=-16'd20983;
      93402:data<=-16'd17597;
      93403:data<=-16'd17500;
      93404:data<=-16'd17033;
      93405:data<=-16'd15803;
      93406:data<=-16'd15494;
      93407:data<=-16'd14795;
      93408:data<=-16'd14251;
      93409:data<=-16'd13268;
      93410:data<=-16'd12072;
      93411:data<=-16'd11433;
      93412:data<=-16'd11555;
      93413:data<=-16'd12918;
      93414:data<=-16'd12965;
      93415:data<=-16'd11442;
      93416:data<=-16'd10705;
      93417:data<=-16'd9661;
      93418:data<=-16'd8593;
      93419:data<=-16'd8175;
      93420:data<=-16'd7348;
      93421:data<=-16'd6930;
      93422:data<=-16'd6552;
      93423:data<=-16'd5698;
      93424:data<=-16'd5253;
      93425:data<=-16'd5336;
      93426:data<=-16'd6454;
      93427:data<=-16'd6831;
      93428:data<=-16'd5482;
      93429:data<=-16'd5110;
      93430:data<=-16'd4951;
      93431:data<=-16'd4108;
      93432:data<=-16'd3935;
      93433:data<=-16'd3425;
      93434:data<=-16'd2895;
      93435:data<=-16'd2488;
      93436:data<=-16'd1569;
      93437:data<=-16'd1316;
      93438:data<=-16'd1143;
      93439:data<=-16'd2099;
      93440:data<=-16'd3600;
      93441:data<=-16'd2235;
      93442:data<=-16'd2490;
      93443:data<=-16'd2370;
      93444:data<=16'd6363;
      93445:data<=16'd14225;
      93446:data<=16'd15141;
      93447:data<=16'd17588;
      93448:data<=16'd19358;
      93449:data<=16'd17238;
      93450:data<=16'd16392;
      93451:data<=16'd16674;
      93452:data<=16'd15926;
      93453:data<=16'd13954;
      93454:data<=16'd12339;
      93455:data<=16'd13091;
      93456:data<=16'd13359;
      93457:data<=16'd12505;
      93458:data<=16'd12445;
      93459:data<=16'd11734;
      93460:data<=16'd11256;
      93461:data<=16'd11438;
      93462:data<=16'd10593;
      93463:data<=16'd10005;
      93464:data<=16'd9855;
      93465:data<=16'd9771;
      93466:data<=16'd9956;
      93467:data<=16'd9439;
      93468:data<=16'd9089;
      93469:data<=16'd8862;
      93470:data<=16'd8504;
      93471:data<=16'd8689;
      93472:data<=16'd7515;
      93473:data<=16'd6595;
      93474:data<=16'd7630;
      93475:data<=16'd7523;
      93476:data<=16'd7183;
      93477:data<=16'd7218;
      93478:data<=16'd6690;
      93479:data<=16'd7711;
      93480:data<=16'd8338;
      93481:data<=16'd7846;
      93482:data<=16'd7853;
      93483:data<=16'd6893;
      93484:data<=16'd7094;
      93485:data<=16'd7269;
      93486:data<=16'd5949;
      93487:data<=16'd7655;
      93488:data<=16'd4466;
      93489:data<=-16'd6520;
      93490:data<=-16'd10176;
      93491:data<=-16'd7603;
      93492:data<=-16'd7295;
      93493:data<=-16'd6034;
      93494:data<=-16'd5324;
      93495:data<=-16'd5579;
      93496:data<=-16'd4478;
      93497:data<=-16'd4719;
      93498:data<=-16'd4761;
      93499:data<=-16'd4783;
      93500:data<=-16'd7047;
      93501:data<=-16'd8035;
      93502:data<=-16'd7893;
      93503:data<=-16'd7834;
      93504:data<=-16'd6601;
      93505:data<=-16'd5594;
      93506:data<=-16'd4548;
      93507:data<=-16'd3730;
      93508:data<=-16'd3704;
      93509:data<=-16'd2648;
      93510:data<=-16'd2405;
      93511:data<=-16'd3080;
      93512:data<=-16'd2378;
      93513:data<=-16'd2038;
      93514:data<=-16'd1897;
      93515:data<=-16'd1498;
      93516:data<=-16'd1829;
      93517:data<=-16'd1522;
      93518:data<=-16'd863;
      93519:data<=16'd188;
      93520:data<=16'd1463;
      93521:data<=16'd1077;
      93522:data<=16'd1468;
      93523:data<=16'd2877;
      93524:data<=16'd2823;
      93525:data<=16'd2839;
      93526:data<=16'd2596;
      93527:data<=16'd2546;
      93528:data<=16'd3019;
      93529:data<=16'd1451;
      93530:data<=16'd1630;
      93531:data<=16'd2786;
      93532:data<=16'd1589;
      93533:data<=16'd7944;
      93534:data<=16'd18991;
      93535:data<=16'd20212;
      93536:data<=16'd17649;
      93537:data<=16'd18119;
      93538:data<=16'd17101;
      93539:data<=16'd16333;
      93540:data<=16'd16201;
      93541:data<=16'd14783;
      93542:data<=16'd14405;
      93543:data<=16'd14088;
      93544:data<=16'd13123;
      93545:data<=16'd13559;
      93546:data<=16'd14504;
      93547:data<=16'd14416;
      93548:data<=16'd13335;
      93549:data<=16'd12665;
      93550:data<=16'd12481;
      93551:data<=16'd11047;
      93552:data<=16'd10422;
      93553:data<=16'd12410;
      93554:data<=16'd13955;
      93555:data<=16'd13550;
      93556:data<=16'd12490;
      93557:data<=16'd11850;
      93558:data<=16'd12340;
      93559:data<=16'd13458;
      93560:data<=16'd13391;
      93561:data<=16'd11937;
      93562:data<=16'd11668;
      93563:data<=16'd12044;
      93564:data<=16'd10504;
      93565:data<=16'd9552;
      93566:data<=16'd9727;
      93567:data<=16'd8434;
      93568:data<=16'd7765;
      93569:data<=16'd7871;
      93570:data<=16'd6845;
      93571:data<=16'd6602;
      93572:data<=16'd7700;
      93573:data<=16'd8762;
      93574:data<=16'd7777;
      93575:data<=16'd6288;
      93576:data<=16'd8070;
      93577:data<=16'd5090;
      93578:data<=-16'd5940;
      93579:data<=-16'd11126;
      93580:data<=-16'd9597;
      93581:data<=-16'd9726;
      93582:data<=-16'd9165;
      93583:data<=-16'd8851;
      93584:data<=-16'd9536;
      93585:data<=-16'd7532;
      93586:data<=-16'd6205;
      93587:data<=-16'd6573;
      93588:data<=-16'd6166;
      93589:data<=-16'd6114;
      93590:data<=-16'd5841;
      93591:data<=-16'd6003;
      93592:data<=-16'd6840;
      93593:data<=-16'd5973;
      93594:data<=-16'd5297;
      93595:data<=-16'd5535;
      93596:data<=-16'd5183;
      93597:data<=-16'd5228;
      93598:data<=-16'd4717;
      93599:data<=-16'd3550;
      93600:data<=-16'd3415;
      93601:data<=-16'd3381;
      93602:data<=-16'd2940;
      93603:data<=-16'd2637;
      93604:data<=-16'd2855;
      93605:data<=-16'd3422;
      93606:data<=-16'd4397;
      93607:data<=-16'd6696;
      93608:data<=-16'd7741;
      93609:data<=-16'd6831;
      93610:data<=-16'd7115;
      93611:data<=-16'd6216;
      93612:data<=-16'd3935;
      93613:data<=-16'd3806;
      93614:data<=-16'd3918;
      93615:data<=-16'd4038;
      93616:data<=-16'd3965;
      93617:data<=-16'd2943;
      93618:data<=-16'd4256;
      93619:data<=-16'd4341;
      93620:data<=-16'd2946;
      93621:data<=-16'd5231;
      93622:data<=-16'd1048;
      93623:data<=16'd10513;
      93624:data<=16'd13590;
      93625:data<=16'd11421;
      93626:data<=16'd12157;
      93627:data<=16'd11565;
      93628:data<=16'd10684;
      93629:data<=16'd10646;
      93630:data<=16'd9532;
      93631:data<=16'd9215;
      93632:data<=16'd9053;
      93633:data<=16'd8382;
      93634:data<=16'd8348;
      93635:data<=16'd7937;
      93636:data<=16'd7197;
      93637:data<=16'd6724;
      93638:data<=16'd6963;
      93639:data<=16'd7755;
      93640:data<=16'd7165;
      93641:data<=16'd6002;
      93642:data<=16'd5583;
      93643:data<=16'd4934;
      93644:data<=16'd4575;
      93645:data<=16'd4561;
      93646:data<=16'd4170;
      93647:data<=16'd3847;
      93648:data<=16'd3509;
      93649:data<=16'd2907;
      93650:data<=16'd2127;
      93651:data<=16'd2420;
      93652:data<=16'd3947;
      93653:data<=16'd3979;
      93654:data<=16'd3077;
      93655:data<=16'd2726;
      93656:data<=16'd1692;
      93657:data<=16'd1219;
      93658:data<=16'd1773;
      93659:data<=16'd2645;
      93660:data<=16'd4211;
      93661:data<=16'd4449;
      93662:data<=16'd4252;
      93663:data<=16'd4466;
      93664:data<=16'd3283;
      93665:data<=16'd4422;
      93666:data<=16'd3993;
      93667:data<=-16'd5133;
      93668:data<=-16'd12198;
      93669:data<=-16'd11662;
      93670:data<=-16'd11386;
      93671:data<=-16'd10966;
      93672:data<=-16'd10228;
      93673:data<=-16'd10918;
      93674:data<=-16'd10003;
      93675:data<=-16'd9257;
      93676:data<=-16'd9765;
      93677:data<=-16'd9565;
      93678:data<=-16'd9682;
      93679:data<=-16'd9433;
      93680:data<=-16'd9329;
      93681:data<=-16'd10081;
      93682:data<=-16'd9401;
      93683:data<=-16'd8721;
      93684:data<=-16'd8809;
      93685:data<=-16'd8320;
      93686:data<=-16'd8050;
      93687:data<=-16'd7456;
      93688:data<=-16'd7386;
      93689:data<=-16'd8008;
      93690:data<=-16'd7159;
      93691:data<=-16'd7457;
      93692:data<=-16'd9125;
      93693:data<=-16'd8813;
      93694:data<=-16'd8255;
      93695:data<=-16'd8596;
      93696:data<=-16'd8728;
      93697:data<=-16'd8281;
      93698:data<=-16'd7288;
      93699:data<=-16'd7016;
      93700:data<=-16'd6865;
      93701:data<=-16'd6692;
      93702:data<=-16'd6918;
      93703:data<=-16'd6111;
      93704:data<=-16'd6657;
      93705:data<=-16'd7956;
      93706:data<=-16'd7040;
      93707:data<=-16'd7300;
      93708:data<=-16'd6764;
      93709:data<=-16'd5422;
      93710:data<=-16'd7688;
      93711:data<=-16'd3221;
      93712:data<=16'd7307;
      93713:data<=16'd7652;
      93714:data<=16'd3924;
      93715:data<=16'd4827;
      93716:data<=16'd4234;
      93717:data<=16'd3021;
      93718:data<=16'd2443;
      93719:data<=16'd1189;
      93720:data<=16'd1428;
      93721:data<=16'd1275;
      93722:data<=16'd769;
      93723:data<=16'd1407;
      93724:data<=16'd928;
      93725:data<=16'd555;
      93726:data<=16'd708;
      93727:data<=-16'd141;
      93728:data<=-16'd209;
      93729:data<=16'd308;
      93730:data<=-16'd77;
      93731:data<=-16'd1277;
      93732:data<=-16'd2463;
      93733:data<=-16'd2209;
      93734:data<=-16'd1613;
      93735:data<=-16'd1717;
      93736:data<=-16'd1774;
      93737:data<=-16'd1905;
      93738:data<=-16'd1509;
      93739:data<=-16'd1134;
      93740:data<=-16'd1468;
      93741:data<=-16'd1371;
      93742:data<=-16'd1588;
      93743:data<=-16'd1700;
      93744:data<=-16'd1789;
      93745:data<=-16'd3788;
      93746:data<=-16'd4585;
      93747:data<=-16'd3862;
      93748:data<=-16'd4595;
      93749:data<=-16'd4323;
      93750:data<=-16'd3762;
      93751:data<=-16'd4081;
      93752:data<=-16'd3391;
      93753:data<=-16'd4231;
      93754:data<=-16'd4041;
      93755:data<=-16'd2224;
      93756:data<=-16'd8505;
      93757:data<=-16'd18163;
      93758:data<=-16'd19790;
      93759:data<=-16'd18403;
      93760:data<=-16'd18518;
      93761:data<=-16'd17741;
      93762:data<=-16'd16713;
      93763:data<=-16'd16213;
      93764:data<=-16'd16043;
      93765:data<=-16'd14710;
      93766:data<=-16'd11562;
      93767:data<=-16'd9367;
      93768:data<=-16'd8558;
      93769:data<=-16'd8090;
      93770:data<=-16'd8226;
      93771:data<=-16'd8608;
      93772:data<=-16'd9288;
      93773:data<=-16'd9226;
      93774:data<=-16'd7888;
      93775:data<=-16'd7382;
      93776:data<=-16'd7521;
      93777:data<=-16'd7134;
      93778:data<=-16'd6669;
      93779:data<=-16'd6240;
      93780:data<=-16'd5915;
      93781:data<=-16'd5382;
      93782:data<=-16'd5065;
      93783:data<=-16'd5159;
      93784:data<=-16'd5075;
      93785:data<=-16'd6405;
      93786:data<=-16'd7326;
      93787:data<=-16'd5700;
      93788:data<=-16'd5621;
      93789:data<=-16'd5849;
      93790:data<=-16'd4147;
      93791:data<=-16'd4496;
      93792:data<=-16'd4736;
      93793:data<=-16'd3289;
      93794:data<=-16'd3065;
      93795:data<=-16'd2393;
      93796:data<=-16'd2077;
      93797:data<=-16'd2309;
      93798:data<=-16'd2353;
      93799:data<=-16'd4918;
      93800:data<=-16'd1747;
      93801:data<=16'd9597;
      93802:data<=16'd14210;
      93803:data<=16'd12542;
      93804:data<=16'd12649;
      93805:data<=16'd11559;
      93806:data<=16'd10828;
      93807:data<=16'd11238;
      93808:data<=16'd10470;
      93809:data<=16'd10504;
      93810:data<=16'd9450;
      93811:data<=16'd7635;
      93812:data<=16'd7724;
      93813:data<=16'd7468;
      93814:data<=16'd7793;
      93815:data<=16'd8291;
      93816:data<=16'd7221;
      93817:data<=16'd7356;
      93818:data<=16'd6485;
      93819:data<=16'd3673;
      93820:data<=16'd2745;
      93821:data<=16'd2500;
      93822:data<=16'd2359;
      93823:data<=16'd1644;
      93824:data<=-16'd723;
      93825:data<=-16'd999;
      93826:data<=-16'd77;
      93827:data<=-16'd162;
      93828:data<=16'd470;
      93829:data<=16'd437;
      93830:data<=16'd196;
      93831:data<=16'd864;
      93832:data<=16'd886;
      93833:data<=16'd127;
      93834:data<=-16'd2378;
      93835:data<=-16'd3664;
      93836:data<=-16'd2156;
      93837:data<=-16'd3245;
      93838:data<=-16'd4197;
      93839:data<=-16'd3316;
      93840:data<=-16'd4531;
      93841:data<=-16'd3911;
      93842:data<=-16'd3601;
      93843:data<=-16'd4602;
      93844:data<=-16'd1318;
      93845:data<=-16'd5363;
      93846:data<=-16'd17399;
      93847:data<=-16'd19114;
      93848:data<=-16'd15641;
      93849:data<=-16'd15952;
      93850:data<=-16'd15082;
      93851:data<=-16'd15258;
      93852:data<=-16'd15916;
      93853:data<=-16'd14277;
      93854:data<=-16'd13681;
      93855:data<=-16'd12753;
      93856:data<=-16'd11574;
      93857:data<=-16'd11812;
      93858:data<=-16'd10968;
      93859:data<=-16'd9988;
      93860:data<=-16'd9905;
      93861:data<=-16'd9647;
      93862:data<=-16'd8854;
      93863:data<=-16'd7706;
      93864:data<=-16'd8431;
      93865:data<=-16'd9060;
      93866:data<=-16'd7327;
      93867:data<=-16'd6796;
      93868:data<=-16'd6816;
      93869:data<=-16'd5809;
      93870:data<=-16'd5348;
      93871:data<=-16'd5130;
      93872:data<=-16'd5045;
      93873:data<=-16'd2100;
      93874:data<=16'd3344;
      93875:data<=16'd4910;
      93876:data<=16'd4476;
      93877:data<=16'd3924;
      93878:data<=16'd2090;
      93879:data<=16'd3051;
      93880:data<=16'd4323;
      93881:data<=16'd3204;
      93882:data<=16'd3265;
      93883:data<=16'd3460;
      93884:data<=16'd4220;
      93885:data<=16'd5148;
      93886:data<=16'd4749;
      93887:data<=16'd5765;
      93888:data<=16'd4510;
      93889:data<=16'd5216;
      93890:data<=16'd15659;
      93891:data<=16'd21682;
      93892:data<=16'd19226;
      93893:data<=16'd19226;
      93894:data<=16'd18202;
      93895:data<=16'd16968;
      93896:data<=16'd18304;
      93897:data<=16'd16698;
      93898:data<=16'd15898;
      93899:data<=16'd16528;
      93900:data<=16'd15076;
      93901:data<=16'd15088;
      93902:data<=16'd15139;
      93903:data<=16'd15068;
      93904:data<=16'd16322;
      93905:data<=16'd15532;
      93906:data<=16'd14904;
      93907:data<=16'd14718;
      93908:data<=16'd13302;
      93909:data<=16'd13611;
      93910:data<=16'd13581;
      93911:data<=16'd12989;
      93912:data<=16'd13203;
      93913:data<=16'd11840;
      93914:data<=16'd11515;
      93915:data<=16'd11462;
      93916:data<=16'd10339;
      93917:data<=16'd11953;
      93918:data<=16'd12257;
      93919:data<=16'd10636;
      93920:data<=16'd11079;
      93921:data<=16'd10686;
      93922:data<=16'd10608;
      93923:data<=16'd10246;
      93924:data<=16'd8364;
      93925:data<=16'd9286;
      93926:data<=16'd6854;
      93927:data<=16'd497;
      93928:data<=-16'd564;
      93929:data<=-16'd121;
      93930:data<=16'd438;
      93931:data<=16'd1876;
      93932:data<=16'd646;
      93933:data<=16'd1950;
      93934:data<=-16'd106;
      93935:data<=-16'd11229;
      93936:data<=-16'd15470;
      93937:data<=-16'd12474;
      93938:data<=-16'd12640;
      93939:data<=-16'd11864;
      93940:data<=-16'd10859;
      93941:data<=-16'd10985;
      93942:data<=-16'd9383;
      93943:data<=-16'd8648;
      93944:data<=-16'd7641;
      93945:data<=-16'd6332;
      93946:data<=-16'd6724;
      93947:data<=-16'd5742;
      93948:data<=-16'd5083;
      93949:data<=-16'd5738;
      93950:data<=-16'd4987;
      93951:data<=-16'd4924;
      93952:data<=-16'd5178;
      93953:data<=-16'd4636;
      93954:data<=-16'd4564;
      93955:data<=-16'd3667;
      93956:data<=-16'd2889;
      93957:data<=-16'd2367;
      93958:data<=-16'd928;
      93959:data<=-16'd1048;
      93960:data<=-16'd1460;
      93961:data<=-16'd647;
      93962:data<=-16'd785;
      93963:data<=-16'd977;
      93964:data<=-16'd644;
      93965:data<=-16'd214;
      93966:data<=-16'd27;
      93967:data<=-16'd860;
      93968:data<=-16'd221;
      93969:data<=16'd1313;
      93970:data<=16'd1530;
      93971:data<=16'd2343;
      93972:data<=16'd2397;
      93973:data<=16'd1938;
      93974:data<=16'd2893;
      93975:data<=16'd2590;
      93976:data<=16'd2767;
      93977:data<=16'd2660;
      93978:data<=16'd1823;
      93979:data<=16'd11179;
      93980:data<=16'd24328;
      93981:data<=16'd25161;
      93982:data<=16'd22848;
      93983:data<=16'd24570;
      93984:data<=16'd23579;
      93985:data<=16'd22403;
      93986:data<=16'd22363;
      93987:data<=16'd20682;
      93988:data<=16'd19901;
      93989:data<=16'd19716;
      93990:data<=16'd18375;
      93991:data<=16'd17065;
      93992:data<=16'd16877;
      93993:data<=16'd17476;
      93994:data<=16'd16706;
      93995:data<=16'd15318;
      93996:data<=16'd15584;
      93997:data<=16'd16315;
      93998:data<=16'd16057;
      93999:data<=16'd14148;
      94000:data<=16'd12704;
      94001:data<=16'd13441;
      94002:data<=16'd12539;
      94003:data<=16'd10947;
      94004:data<=16'd11694;
      94005:data<=16'd11085;
      94006:data<=16'd9727;
      94007:data<=16'd9978;
      94008:data<=16'd9394;
      94009:data<=16'd9182;
      94010:data<=16'd10119;
      94011:data<=16'd9662;
      94012:data<=16'd8476;
      94013:data<=16'd8025;
      94014:data<=16'd7724;
      94015:data<=16'd6693;
      94016:data<=16'd6166;
      94017:data<=16'd6261;
      94018:data<=16'd5139;
      94019:data<=16'd5212;
      94020:data<=16'd5338;
      94021:data<=16'd3334;
      94022:data<=16'd4833;
      94023:data<=16'd3275;
      94024:data<=-16'd7476;
      94025:data<=-16'd12152;
      94026:data<=-16'd9793;
      94027:data<=-16'd10558;
      94028:data<=-16'd9464;
      94029:data<=-16'd8954;
      94030:data<=-16'd11103;
      94031:data<=-16'd8862;
      94032:data<=-16'd9682;
      94033:data<=-16'd15658;
      94034:data<=-16'd17203;
      94035:data<=-16'd16898;
      94036:data<=-16'd16201;
      94037:data<=-16'd13261;
      94038:data<=-16'd12640;
      94039:data<=-16'd13496;
      94040:data<=-16'd13083;
      94041:data<=-16'd12536;
      94042:data<=-16'd11917;
      94043:data<=-16'd11379;
      94044:data<=-16'd10818;
      94045:data<=-16'd10822;
      94046:data<=-16'd11236;
      94047:data<=-16'd10733;
      94048:data<=-16'd10777;
      94049:data<=-16'd9928;
      94050:data<=-16'd7468;
      94051:data<=-16'd7476;
      94052:data<=-16'd7746;
      94053:data<=-16'd6472;
      94054:data<=-16'd6666;
      94055:data<=-16'd6481;
      94056:data<=-16'd5868;
      94057:data<=-16'd6478;
      94058:data<=-16'd6138;
      94059:data<=-16'd5444;
      94060:data<=-16'd5720;
      94061:data<=-16'd6155;
      94062:data<=-16'd5335;
      94063:data<=-16'd3362;
      94064:data<=-16'd3331;
      94065:data<=-16'd3500;
      94066:data<=-16'd3140;
      94067:data<=-16'd4698;
      94068:data<=16'd256;
      94069:data<=16'd10986;
      94070:data<=16'd12897;
      94071:data<=16'd9931;
      94072:data<=16'd10199;
      94073:data<=16'd9523;
      94074:data<=16'd9306;
      94075:data<=16'd10122;
      94076:data<=16'd9270;
      94077:data<=16'd9224;
      94078:data<=16'd9285;
      94079:data<=16'd8766;
      94080:data<=16'd9012;
      94081:data<=16'd8410;
      94082:data<=16'd8100;
      94083:data<=16'd7959;
      94084:data<=16'd6308;
      94085:data<=16'd7357;
      94086:data<=16'd11492;
      94087:data<=16'd13207;
      94088:data<=16'd12314;
      94089:data<=16'd12134;
      94090:data<=16'd12800;
      94091:data<=16'd12527;
      94092:data<=16'd11670;
      94093:data<=16'd11244;
      94094:data<=16'd10393;
      94095:data<=16'd9077;
      94096:data<=16'd8346;
      94097:data<=16'd8296;
      94098:data<=16'd7874;
      94099:data<=16'd6904;
      94100:data<=16'd6881;
      94101:data<=16'd6508;
      94102:data<=16'd4739;
      94103:data<=16'd4325;
      94104:data<=16'd4610;
      94105:data<=16'd4053;
      94106:data<=16'd3592;
      94107:data<=16'd2908;
      94108:data<=16'd3002;
      94109:data<=16'd2529;
      94110:data<=16'd984;
      94111:data<=16'd2699;
      94112:data<=16'd960;
      94113:data<=-16'd9031;
      94114:data<=-16'd14815;
      94115:data<=-16'd14340;
      94116:data<=-16'd14894;
      94117:data<=-16'd14824;
      94118:data<=-16'd14659;
      94119:data<=-16'd14962;
      94120:data<=-16'd14160;
      94121:data<=-16'd14458;
      94122:data<=-16'd14040;
      94123:data<=-16'd12660;
      94124:data<=-16'd13086;
      94125:data<=-16'd12794;
      94126:data<=-16'd12392;
      94127:data<=-16'd12936;
      94128:data<=-16'd12334;
      94129:data<=-16'd12839;
      94130:data<=-16'd13758;
      94131:data<=-16'd12939;
      94132:data<=-16'd12687;
      94133:data<=-16'd12158;
      94134:data<=-16'd11168;
      94135:data<=-16'd11615;
      94136:data<=-16'd11665;
      94137:data<=-16'd10831;
      94138:data<=-16'd11453;
      94139:data<=-16'd14927;
      94140:data<=-16'd18454;
      94141:data<=-16'd18387;
      94142:data<=-16'd17796;
      94143:data<=-16'd18199;
      94144:data<=-16'd17139;
      94145:data<=-16'd16339;
      94146:data<=-16'd16104;
      94147:data<=-16'd15791;
      94148:data<=-16'd15688;
      94149:data<=-16'd14196;
      94150:data<=-16'd13776;
      94151:data<=-16'd14181;
      94152:data<=-16'd12696;
      94153:data<=-16'd13069;
      94154:data<=-16'd12736;
      94155:data<=-16'd11298;
      94156:data<=-16'd14832;
      94157:data<=-16'd12069;
      94158:data<=16'd129;
      94159:data<=16'd3849;
      94160:data<=16'd1184;
      94161:data<=16'd2329;
      94162:data<=16'd2602;
      94163:data<=16'd2147;
      94164:data<=16'd2640;
      94165:data<=16'd1701;
      94166:data<=16'd1492;
      94167:data<=16'd1933;
      94168:data<=16'd1193;
      94169:data<=16'd171;
      94170:data<=-16'd484;
      94171:data<=-16'd274;
      94172:data<=-16'd273;
      94173:data<=-16'd795;
      94174:data<=-16'd597;
      94175:data<=-16'd478;
      94176:data<=-16'd281;
      94177:data<=-16'd53;
      94178:data<=-16'd523;
      94179:data<=-16'd129;
      94180:data<=16'd390;
      94181:data<=-16'd127;
      94182:data<=-16'd607;
      94183:data<=-16'd1431;
      94184:data<=-16'd1945;
      94185:data<=-16'd1718;
      94186:data<=-16'd2067;
      94187:data<=-16'd2734;
      94188:data<=-16'd3084;
      94189:data<=-16'd1991;
      94190:data<=-16'd974;
      94191:data<=-16'd1771;
      94192:data<=16'd1157;
      94193:data<=16'd7094;
      94194:data<=16'd8062;
      94195:data<=16'd5749;
      94196:data<=16'd4000;
      94197:data<=16'd3315;
      94198:data<=16'd3770;
      94199:data<=16'd3287;
      94200:data<=16'd4153;
      94201:data<=16'd3871;
      94202:data<=-16'd4555;
      94203:data<=-16'd11661;
      94204:data<=-16'd10642;
      94205:data<=-16'd9853;
      94206:data<=-16'd9868;
      94207:data<=-16'd9053;
      94208:data<=-16'd9779;
      94209:data<=-16'd10185;
      94210:data<=-16'd10254;
      94211:data<=-16'd9893;
      94212:data<=-16'd8857;
      94213:data<=-16'd9400;
      94214:data<=-16'd9139;
      94215:data<=-16'd7843;
      94216:data<=-16'd7771;
      94217:data<=-16'd6924;
      94218:data<=-16'd6613;
      94219:data<=-16'd6902;
      94220:data<=-16'd5360;
      94221:data<=-16'd5151;
      94222:data<=-16'd6387;
      94223:data<=-16'd6560;
      94224:data<=-16'd6375;
      94225:data<=-16'd5715;
      94226:data<=-16'd5735;
      94227:data<=-16'd6190;
      94228:data<=-16'd5207;
      94229:data<=-16'd4466;
      94230:data<=-16'd4023;
      94231:data<=-16'd3547;
      94232:data<=-16'd3421;
      94233:data<=-16'd2431;
      94234:data<=-16'd2276;
      94235:data<=-16'd2895;
      94236:data<=-16'd3397;
      94237:data<=-16'd4696;
      94238:data<=-16'd3422;
      94239:data<=-16'd2011;
      94240:data<=-16'd3600;
      94241:data<=-16'd2652;
      94242:data<=-16'd2035;
      94243:data<=-16'd2745;
      94244:data<=-16'd1256;
      94245:data<=-16'd5292;
      94246:data<=-16'd7209;
      94247:data<=16'd2863;
      94248:data<=16'd7077;
      94249:data<=16'd2881;
      94250:data<=16'd3516;
      94251:data<=16'd4140;
      94252:data<=16'd3328;
      94253:data<=16'd4021;
      94254:data<=16'd3201;
      94255:data<=16'd3374;
      94256:data<=16'd3971;
      94257:data<=16'd3131;
      94258:data<=16'd3284;
      94259:data<=16'd2751;
      94260:data<=16'd2463;
      94261:data<=16'd3341;
      94262:data<=16'd2655;
      94263:data<=16'd2247;
      94264:data<=16'd1991;
      94265:data<=16'd1389;
      94266:data<=16'd2235;
      94267:data<=16'd1886;
      94268:data<=16'd1516;
      94269:data<=16'd2795;
      94270:data<=16'd2423;
      94271:data<=16'd2033;
      94272:data<=16'd2385;
      94273:data<=16'd1935;
      94274:data<=16'd2146;
      94275:data<=16'd1635;
      94276:data<=16'd611;
      94277:data<=16'd708;
      94278:data<=16'd467;
      94279:data<=16'd737;
      94280:data<=16'd1289;
      94281:data<=16'd1586;
      94282:data<=16'd2234;
      94283:data<=16'd1172;
      94284:data<=16'd584;
      94285:data<=16'd1221;
      94286:data<=16'd691;
      94287:data<=16'd1889;
      94288:data<=16'd1516;
      94289:data<=-16'd687;
      94290:data<=16'd1463;
      94291:data<=-16'd2695;
      94292:data<=-16'd13752;
      94293:data<=-16'd14885;
      94294:data<=-16'd11935;
      94295:data<=-16'd12722;
      94296:data<=-16'd11539;
      94297:data<=-16'd11230;
      94298:data<=-16'd9397;
      94299:data<=-16'd2936;
      94300:data<=-16'd432;
      94301:data<=-16'd887;
      94302:data<=-16'd513;
      94303:data<=-16'd1612;
      94304:data<=-16'd1541;
      94305:data<=-16'd704;
      94306:data<=-16'd1024;
      94307:data<=-16'd587;
      94308:data<=-16'd795;
      94309:data<=-16'd842;
      94310:data<=16'd832;
      94311:data<=16'd1368;
      94312:data<=16'd1171;
      94313:data<=16'd1383;
      94314:data<=16'd1128;
      94315:data<=16'd1318;
      94316:data<=16'd1862;
      94317:data<=16'd2096;
      94318:data<=16'd2161;
      94319:data<=16'd2170;
      94320:data<=16'd2752;
      94321:data<=16'd3146;
      94322:data<=16'd2823;
      94323:data<=16'd2954;
      94324:data<=16'd3189;
      94325:data<=16'd2974;
      94326:data<=16'd3008;
      94327:data<=16'd3598;
      94328:data<=16'd4652;
      94329:data<=16'd5970;
      94330:data<=16'd6379;
      94331:data<=16'd5137;
      94332:data<=16'd5113;
      94333:data<=16'd6261;
      94334:data<=16'd4852;
      94335:data<=16'd7350;
      94336:data<=16'd17004;
      94337:data<=16'd21256;
      94338:data<=16'd19297;
      94339:data<=16'd19658;
      94340:data<=16'd19012;
      94341:data<=16'd18190;
      94342:data<=16'd19866;
      94343:data<=16'd18654;
      94344:data<=16'd17042;
      94345:data<=16'd17417;
      94346:data<=16'd16120;
      94347:data<=16'd15535;
      94348:data<=16'd15245;
      94349:data<=16'd14101;
      94350:data<=16'd15218;
      94351:data<=16'd13314;
      94352:data<=16'd7010;
      94353:data<=16'd4763;
      94354:data<=16'd5636;
      94355:data<=16'd5668;
      94356:data<=16'd6328;
      94357:data<=16'd6423;
      94358:data<=16'd5780;
      94359:data<=16'd5773;
      94360:data<=16'd5192;
      94361:data<=16'd4895;
      94362:data<=16'd5524;
      94363:data<=16'd5131;
      94364:data<=16'd4808;
      94365:data<=16'd5377;
      94366:data<=16'd4535;
      94367:data<=16'd3938;
      94368:data<=16'd5554;
      94369:data<=16'd6024;
      94370:data<=16'd5071;
      94371:data<=16'd5015;
      94372:data<=16'd4892;
      94373:data<=16'd4807;
      94374:data<=16'd4358;
      94375:data<=16'd3529;
      94376:data<=16'd4684;
      94377:data<=16'd4528;
      94378:data<=16'd3159;
      94379:data<=16'd4833;
      94380:data<=16'd1011;
      94381:data<=-16'd8760;
      94382:data<=-16'd10293;
      94383:data<=-16'd7544;
      94384:data<=-16'd8971;
      94385:data<=-16'd8707;
      94386:data<=-16'd7210;
      94387:data<=-16'd7427;
      94388:data<=-16'd6871;
      94389:data<=-16'd6787;
      94390:data<=-16'd6495;
      94391:data<=-16'd5134;
      94392:data<=-16'd5598;
      94393:data<=-16'd6029;
      94394:data<=-16'd4517;
      94395:data<=-16'd2761;
      94396:data<=-16'd1644;
      94397:data<=-16'd2159;
      94398:data<=-16'd2802;
      94399:data<=-16'd2297;
      94400:data<=-16'd2532;
      94401:data<=-16'd2074;
      94402:data<=-16'd1266;
      94403:data<=-16'd2655;
      94404:data<=-16'd995;
      94405:data<=16'd4751;
      94406:data<=16'd6646;
      94407:data<=16'd6026;
      94408:data<=16'd7717;
      94409:data<=16'd8070;
      94410:data<=16'd7077;
      94411:data<=16'd7817;
      94412:data<=16'd7820;
      94413:data<=16'd6924;
      94414:data<=16'd6692;
      94415:data<=16'd6137;
      94416:data<=16'd6363;
      94417:data<=16'd6802;
      94418:data<=16'd6003;
      94419:data<=16'd5887;
      94420:data<=16'd5809;
      94421:data<=16'd6196;
      94422:data<=16'd8079;
      94423:data<=16'd7460;
      94424:data<=16'd8317;
      94425:data<=16'd15957;
      94426:data<=16'd21349;
      94427:data<=16'd20501;
      94428:data<=16'd19206;
      94429:data<=16'd17932;
      94430:data<=16'd17293;
      94431:data<=16'd17757;
      94432:data<=16'd16468;
      94433:data<=16'd15050;
      94434:data<=16'd15493;
      94435:data<=16'd16401;
      94436:data<=16'd16662;
      94437:data<=16'd15396;
      94438:data<=16'd13791;
      94439:data<=16'd13145;
      94440:data<=16'd12622;
      94441:data<=16'd12292;
      94442:data<=16'd11673;
      94443:data<=16'd10472;
      94444:data<=16'd10158;
      94445:data<=16'd10067;
      94446:data<=16'd9168;
      94447:data<=16'd9124;
      94448:data<=16'd10433;
      94449:data<=16'd10681;
      94450:data<=16'd9464;
      94451:data<=16'd8819;
      94452:data<=16'd8072;
      94453:data<=16'd7329;
      94454:data<=16'd7514;
      94455:data<=16'd6103;
      94456:data<=16'd5416;
      94457:data<=16'd6023;
      94458:data<=16'd980;
      94459:data<=-16'd4435;
      94460:data<=-16'd3742;
      94461:data<=-16'd3541;
      94462:data<=-16'd3060;
      94463:data<=-16'd1362;
      94464:data<=-16'd2537;
      94465:data<=-16'd2012;
      94466:data<=-16'd1927;
      94467:data<=-16'd3870;
      94468:data<=-16'd1212;
      94469:data<=-16'd4467;
      94470:data<=-16'd16318;
      94471:data<=-16'd19318;
      94472:data<=-16'd16932;
      94473:data<=-16'd18183;
      94474:data<=-16'd16821;
      94475:data<=-16'd14192;
      94476:data<=-16'd13884;
      94477:data<=-16'd13775;
      94478:data<=-16'd13399;
      94479:data<=-16'd12025;
      94480:data<=-16'd11667;
      94481:data<=-16'd12778;
      94482:data<=-16'd12070;
      94483:data<=-16'd11083;
      94484:data<=-16'd10894;
      94485:data<=-16'd11106;
      94486:data<=-16'd12064;
      94487:data<=-16'd10886;
      94488:data<=-16'd8772;
      94489:data<=-16'd8731;
      94490:data<=-16'd8625;
      94491:data<=-16'd8219;
      94492:data<=-16'd8069;
      94493:data<=-16'd7644;
      94494:data<=-16'd7665;
      94495:data<=-16'd7603;
      94496:data<=-16'd7371;
      94497:data<=-16'd6792;
      94498:data<=-16'd6388;
      94499:data<=-16'd7460;
      94500:data<=-16'd6719;
      94501:data<=-16'd4654;
      94502:data<=-16'd4980;
      94503:data<=-16'd4849;
      94504:data<=-16'd4235;
      94505:data<=-16'd4032;
      94506:data<=-16'd2692;
      94507:data<=-16'd3151;
      94508:data<=-16'd3536;
      94509:data<=-16'd3168;
      94510:data<=-16'd4842;
      94511:data<=-16'd986;
      94512:data<=16'd4790;
      94513:data<=16'd3980;
      94514:data<=16'd9570;
      94515:data<=16'd20410;
      94516:data<=16'd21114;
      94517:data<=16'd18481;
      94518:data<=16'd18192;
      94519:data<=16'd16393;
      94520:data<=16'd15920;
      94521:data<=16'd15558;
      94522:data<=16'd14164;
      94523:data<=16'd13966;
      94524:data<=16'd12842;
      94525:data<=16'd11890;
      94526:data<=16'd11826;
      94527:data<=16'd10358;
      94528:data<=16'd9541;
      94529:data<=16'd9770;
      94530:data<=16'd9615;
      94531:data<=16'd9094;
      94532:data<=16'd7494;
      94533:data<=16'd6757;
      94534:data<=16'd7386;
      94535:data<=16'd6777;
      94536:data<=16'd5996;
      94537:data<=16'd5745;
      94538:data<=16'd4728;
      94539:data<=16'd3896;
      94540:data<=16'd3413;
      94541:data<=16'd2002;
      94542:data<=16'd698;
      94543:data<=16'd981;
      94544:data<=16'd983;
      94545:data<=16'd71;
      94546:data<=-16'd2;
      94547:data<=-16'd828;
      94548:data<=-16'd1642;
      94549:data<=-16'd811;
      94550:data<=-16'd2235;
      94551:data<=-16'd3615;
      94552:data<=-16'd2326;
      94553:data<=-16'd3078;
      94554:data<=-16'd3659;
      94555:data<=-16'd4038;
      94556:data<=-16'd6105;
      94557:data<=-16'd3783;
      94558:data<=-16'd5694;
      94559:data<=-16'd17399;
      94560:data<=-16'd21755;
      94561:data<=-16'd19440;
      94562:data<=-16'd19926;
      94563:data<=-16'd17878;
      94564:data<=-16'd18853;
      94565:data<=-16'd25059;
      94566:data<=-16'd25901;
      94567:data<=-16'd24811;
      94568:data<=-16'd25513;
      94569:data<=-16'd24533;
      94570:data<=-16'd24190;
      94571:data<=-16'd23851;
      94572:data<=-16'd22573;
      94573:data<=-16'd22322;
      94574:data<=-16'd21673;
      94575:data<=-16'd21068;
      94576:data<=-16'd20724;
      94577:data<=-16'd19581;
      94578:data<=-16'd18886;
      94579:data<=-16'd18187;
      94580:data<=-16'd18268;
      94581:data<=-16'd19644;
      94582:data<=-16'd19317;
      94583:data<=-16'd17907;
      94584:data<=-16'd17064;
      94585:data<=-16'd16439;
      94586:data<=-16'd16316;
      94587:data<=-16'd15817;
      94588:data<=-16'd14956;
      94589:data<=-16'd14510;
      94590:data<=-16'd14634;
      94591:data<=-16'd14721;
      94592:data<=-16'd13013;
      94593:data<=-16'd12674;
      94594:data<=-16'd14489;
      94595:data<=-16'd13224;
      94596:data<=-16'd12198;
      94597:data<=-16'd12891;
      94598:data<=-16'd11270;
      94599:data<=-16'd11230;
      94600:data<=-16'd10854;
      94601:data<=-16'd9042;
      94602:data<=-16'd11306;
      94603:data<=-16'd6660;
      94604:data<=16'd5943;
      94605:data<=16'd8636;
      94606:data<=16'd5636;
      94607:data<=16'd5303;
      94608:data<=16'd3315;
      94609:data<=16'd2963;
      94610:data<=16'd3727;
      94611:data<=16'd3087;
      94612:data<=16'd4440;
      94613:data<=16'd4488;
      94614:data<=16'd3967;
      94615:data<=16'd4940;
      94616:data<=16'd3022;
      94617:data<=16'd4338;
      94618:data<=16'd10796;
      94619:data<=16'd12090;
      94620:data<=16'd9633;
      94621:data<=16'd8601;
      94622:data<=16'd8122;
      94623:data<=16'd8812;
      94624:data<=16'd8828;
      94625:data<=16'd7908;
      94626:data<=16'd8502;
      94627:data<=16'd8478;
      94628:data<=16'd7641;
      94629:data<=16'd7844;
      94630:data<=16'd7583;
      94631:data<=16'd6984;
      94632:data<=16'd6981;
      94633:data<=16'd5870;
      94634:data<=16'd3688;
      94635:data<=16'd3175;
      94636:data<=16'd4055;
      94637:data<=16'd3698;
      94638:data<=16'd2878;
      94639:data<=16'd2739;
      94640:data<=16'd2457;
      94641:data<=16'd2484;
      94642:data<=16'd2887;
      94643:data<=16'd3283;
      94644:data<=16'd3389;
      94645:data<=16'd3307;
      94646:data<=16'd4167;
      94647:data<=16'd837;
      94648:data<=-16'd9426;
      94649:data<=-16'd15584;
      94650:data<=-16'd14386;
      94651:data<=-16'd13693;
      94652:data<=-16'd13204;
      94653:data<=-16'd12240;
      94654:data<=-16'd12067;
      94655:data<=-16'd10742;
      94656:data<=-16'd10568;
      94657:data<=-16'd11103;
      94658:data<=-16'd9439;
      94659:data<=-16'd8966;
      94660:data<=-16'd9599;
      94661:data<=-16'd9676;
      94662:data<=-16'd10595;
      94663:data<=-16'd10014;
      94664:data<=-16'd8486;
      94665:data<=-16'd8343;
      94666:data<=-16'd7829;
      94667:data<=-16'd8062;
      94668:data<=-16'd8105;
      94669:data<=-16'd5947;
      94670:data<=-16'd7749;
      94671:data<=-16'd13392;
      94672:data<=-16'd14489;
      94673:data<=-16'd12968;
      94674:data<=-16'd13916;
      94675:data<=-16'd14233;
      94676:data<=-16'd13174;
      94677:data<=-16'd13027;
      94678:data<=-16'd12031;
      94679:data<=-16'd10924;
      94680:data<=-16'd11470;
      94681:data<=-16'd10658;
      94682:data<=-16'd9479;
      94683:data<=-16'd9462;
      94684:data<=-16'd7324;
      94685:data<=-16'd5835;
      94686:data<=-16'd7056;
      94687:data<=-16'd7571;
      94688:data<=-16'd8483;
      94689:data<=-16'd8056;
      94690:data<=-16'd6304;
      94691:data<=-16'd8069;
      94692:data<=-16'd4121;
      94693:data<=16'd7975;
      94694:data<=16'd11891;
      94695:data<=16'd8918;
      94696:data<=16'd9295;
      94697:data<=16'd9620;
      94698:data<=16'd9354;
      94699:data<=16'd9104;
      94700:data<=16'd7201;
      94701:data<=16'd7042;
      94702:data<=16'd7476;
      94703:data<=16'd6667;
      94704:data<=16'd7316;
      94705:data<=16'd7605;
      94706:data<=16'd7069;
      94707:data<=16'd7662;
      94708:data<=16'd7553;
      94709:data<=16'd6819;
      94710:data<=16'd6724;
      94711:data<=16'd7119;
      94712:data<=16'd7652;
      94713:data<=16'd6407;
      94714:data<=16'd4563;
      94715:data<=16'd4713;
      94716:data<=16'd5084;
      94717:data<=16'd5327;
      94718:data<=16'd6131;
      94719:data<=16'd5920;
      94720:data<=16'd5858;
      94721:data<=16'd6332;
      94722:data<=16'd5133;
      94723:data<=16'd5826;
      94724:data<=16'd11297;
      94725:data<=16'd14663;
      94726:data<=16'd12768;
      94727:data<=16'd11254;
      94728:data<=16'd10780;
      94729:data<=16'd9690;
      94730:data<=16'd9865;
      94731:data<=16'd10022;
      94732:data<=16'd9752;
      94733:data<=16'd10295;
      94734:data<=16'd9817;
      94735:data<=16'd10287;
      94736:data<=16'd10263;
      94737:data<=16'd3051;
      94738:data<=-16'd4323;
      94739:data<=-16'd4067;
      94740:data<=-16'd3045;
      94741:data<=-16'd3457;
      94742:data<=-16'd2373;
      94743:data<=-16'd2087;
      94744:data<=-16'd2400;
      94745:data<=-16'd2053;
      94746:data<=-16'd1867;
      94747:data<=-16'd1387;
      94748:data<=-16'd1083;
      94749:data<=-16'd1042;
      94750:data<=-16'd473;
      94751:data<=-16'd259;
      94752:data<=-16'd118;
      94753:data<=16'd1030;
      94754:data<=16'd2344;
      94755:data<=16'd2648;
      94756:data<=16'd2108;
      94757:data<=16'd1905;
      94758:data<=16'd2265;
      94759:data<=16'd2408;
      94760:data<=16'd2065;
      94761:data<=16'd1660;
      94762:data<=16'd1727;
      94763:data<=16'd1633;
      94764:data<=16'd1384;
      94765:data<=16'd2262;
      94766:data<=16'd3641;
      94767:data<=16'd4598;
      94768:data<=16'd4617;
      94769:data<=16'd3626;
      94770:data<=16'd3811;
      94771:data<=16'd4493;
      94772:data<=16'd4026;
      94773:data<=16'd4000;
      94774:data<=16'd3983;
      94775:data<=16'd4864;
      94776:data<=16'd5166;
      94777:data<=-16'd707;
      94778:data<=-16'd5163;
      94779:data<=-16'd2939;
      94780:data<=-16'd2995;
      94781:data<=-16'd367;
      94782:data<=16'd9030;
      94783:data<=16'd12134;
      94784:data<=16'd10154;
      94785:data<=16'd10736;
      94786:data<=16'd10411;
      94787:data<=16'd9835;
      94788:data<=16'd9606;
      94789:data<=16'd8936;
      94790:data<=16'd10113;
      94791:data<=16'd9908;
      94792:data<=16'd8774;
      94793:data<=16'd10342;
      94794:data<=16'd10422;
      94795:data<=16'd8851;
      94796:data<=16'd8962;
      94797:data<=16'd9209;
      94798:data<=16'd8912;
      94799:data<=16'd7949;
      94800:data<=16'd7219;
      94801:data<=16'd7774;
      94802:data<=16'd7562;
      94803:data<=16'd7313;
      94804:data<=16'd7773;
      94805:data<=16'd7432;
      94806:data<=16'd7928;
      94807:data<=16'd8924;
      94808:data<=16'd8690;
      94809:data<=16'd8587;
      94810:data<=16'd8520;
      94811:data<=16'd8017;
      94812:data<=16'd7656;
      94813:data<=16'd7585;
      94814:data<=16'd7370;
      94815:data<=16'd6220;
      94816:data<=16'd6241;
      94817:data<=16'd7007;
      94818:data<=16'd5520;
      94819:data<=16'd5635;
      94820:data<=16'd7435;
      94821:data<=16'd6672;
      94822:data<=16'd6607;
      94823:data<=16'd6971;
      94824:data<=16'd6575;
      94825:data<=16'd7544;
      94826:data<=16'd3052;
      94827:data<=-16'd5600;
      94828:data<=-16'd7664;
      94829:data<=-16'd6293;
      94830:data<=-16'd3765;
      94831:data<=16'd1924;
      94832:data<=16'd4173;
      94833:data<=16'd3539;
      94834:data<=16'd4222;
      94835:data<=16'd3479;
      94836:data<=16'd3008;
      94837:data<=16'd3695;
      94838:data<=16'd3130;
      94839:data<=16'd3207;
      94840:data<=16'd3300;
      94841:data<=16'd2328;
      94842:data<=16'd2535;
      94843:data<=16'd2728;
      94844:data<=16'd1944;
      94845:data<=16'd2024;
      94846:data<=16'd3119;
      94847:data<=16'd4320;
      94848:data<=16'd4636;
      94849:data<=16'd3715;
      94850:data<=16'd2761;
      94851:data<=16'd2984;
      94852:data<=16'd3845;
      94853:data<=16'd3612;
      94854:data<=16'd2511;
      94855:data<=16'd2115;
      94856:data<=16'd2452;
      94857:data<=16'd2570;
      94858:data<=16'd2068;
      94859:data<=16'd2541;
      94860:data<=16'd4287;
      94861:data<=16'd4593;
      94862:data<=16'd3706;
      94863:data<=16'd3160;
      94864:data<=16'd2968;
      94865:data<=16'd3304;
      94866:data<=16'd2623;
      94867:data<=16'd2214;
      94868:data<=16'd2804;
      94869:data<=16'd255;
      94870:data<=16'd1101;
      94871:data<=16'd10281;
      94872:data<=16'd15223;
      94873:data<=16'd14190;
      94874:data<=16'd15041;
      94875:data<=16'd14179;
      94876:data<=16'd11967;
      94877:data<=16'd11564;
      94878:data<=16'd10625;
      94879:data<=16'd10495;
      94880:data<=16'd9964;
      94881:data<=16'd8687;
      94882:data<=16'd9864;
      94883:data<=16'd7066;
      94884:data<=16'd85;
      94885:data<=-16'd717;
      94886:data<=16'd2014;
      94887:data<=16'd1858;
      94888:data<=16'd1084;
      94889:data<=16'd820;
      94890:data<=16'd622;
      94891:data<=16'd344;
      94892:data<=-16'd103;
      94893:data<=-16'd208;
      94894:data<=-16'd784;
      94895:data<=-16'd1196;
      94896:data<=-16'd626;
      94897:data<=-16'd616;
      94898:data<=-16'd555;
      94899:data<=16'd644;
      94900:data<=16'd1410;
      94901:data<=16'd673;
      94902:data<=-16'd549;
      94903:data<=-16'd966;
      94904:data<=-16'd980;
      94905:data<=-16'd931;
      94906:data<=-16'd1069;
      94907:data<=-16'd1891;
      94908:data<=-16'd1648;
      94909:data<=-16'd1377;
      94910:data<=-16'd2790;
      94911:data<=-16'd2466;
      94912:data<=-16'd1538;
      94913:data<=-16'd805;
      94914:data<=16'd2187;
      94915:data<=-16'd1530;
      94916:data<=-16'd12311;
      94917:data<=-16'd15151;
      94918:data<=-16'd12786;
      94919:data<=-16'd13251;
      94920:data<=-16'd12296;
      94921:data<=-16'd11615;
      94922:data<=-16'd11988;
      94923:data<=-16'd10483;
      94924:data<=-16'd10648;
      94925:data<=-16'd10593;
      94926:data<=-16'd8172;
      94927:data<=-16'd7817;
      94928:data<=-16'd7934;
      94929:data<=-16'd7242;
      94930:data<=-16'd7908;
      94931:data<=-16'd8273;
      94932:data<=-16'd7850;
      94933:data<=-16'd6858;
      94934:data<=-16'd6725;
      94935:data<=-16'd8657;
      94936:data<=-16'd6223;
      94937:data<=16'd525;
      94938:data<=16'd2726;
      94939:data<=16'd2196;
      94940:data<=16'd3192;
      94941:data<=16'd3005;
      94942:data<=16'd2399;
      94943:data<=16'd2522;
      94944:data<=16'd1867;
      94945:data<=16'd1709;
      94946:data<=16'd2200;
      94947:data<=16'd1818;
      94948:data<=16'd1365;
      94949:data<=16'd989;
      94950:data<=16'd205;
      94951:data<=16'd114;
      94952:data<=16'd462;
      94953:data<=16'd494;
      94954:data<=16'd776;
      94955:data<=16'd608;
      94956:data<=16'd273;
      94957:data<=16'd197;
      94958:data<=-16'd1604;
      94959:data<=-16'd857;
      94960:data<=16'd6526;
      94961:data<=16'd11828;
      94962:data<=16'd10913;
      94963:data<=16'd10125;
      94964:data<=16'd9538;
      94965:data<=16'd7677;
      94966:data<=16'd6623;
      94967:data<=16'd6082;
      94968:data<=16'd5885;
      94969:data<=16'd5245;
      94970:data<=16'd4175;
      94971:data<=16'd4690;
      94972:data<=16'd4363;
      94973:data<=16'd2939;
      94974:data<=16'd3363;
      94975:data<=16'd2898;
      94976:data<=16'd1720;
      94977:data<=16'd2364;
      94978:data<=16'd1359;
      94979:data<=-16'd881;
      94980:data<=-16'd1008;
      94981:data<=-16'd983;
      94982:data<=-16'd1908;
      94983:data<=-16'd2472;
      94984:data<=-16'd2185;
      94985:data<=-16'd1927;
      94986:data<=-16'd2992;
      94987:data<=-16'd3233;
      94988:data<=-16'd2206;
      94989:data<=-16'd4811;
      94990:data<=-16'd10387;
      94991:data<=-16'd13186;
      94992:data<=-16'd13606;
      94993:data<=-16'd13987;
      94994:data<=-16'd13004;
      94995:data<=-16'd11991;
      94996:data<=-16'd12765;
      94997:data<=-16'd12669;
      94998:data<=-16'd12125;
      94999:data<=-16'd12507;
      95000:data<=-16'd11394;
      95001:data<=-16'd11044;
      95002:data<=-16'd11359;
      95003:data<=-16'd8630;
      95004:data<=-16'd11382;
      95005:data<=-16'd21435;
      95006:data<=-16'd24958;
      95007:data<=-16'd23097;
      95008:data<=-16'd23830;
      95009:data<=-16'd23196;
      95010:data<=-16'd21209;
      95011:data<=-16'd20562;
      95012:data<=-16'd19890;
      95013:data<=-16'd19866;
      95014:data<=-16'd19455;
      95015:data<=-16'd18305;
      95016:data<=-16'd17902;
      95017:data<=-16'd16968;
      95018:data<=-16'd16906;
      95019:data<=-16'd17984;
      95020:data<=-16'd17437;
      95021:data<=-16'd16774;
      95022:data<=-16'd16152;
      95023:data<=-16'd15139;
      95024:data<=-16'd15515;
      95025:data<=-16'd14903;
      95026:data<=-16'd13573;
      95027:data<=-16'd13934;
      95028:data<=-16'd12947;
      95029:data<=-16'd11126;
      95030:data<=-16'd11217;
      95031:data<=-16'd11668;
      95032:data<=-16'd12019;
      95033:data<=-16'd11835;
      95034:data<=-16'd10672;
      95035:data<=-16'd9981;
      95036:data<=-16'd9485;
      95037:data<=-16'd9033;
      95038:data<=-16'd8640;
      95039:data<=-16'd7436;
      95040:data<=-16'd7057;
      95041:data<=-16'd7735;
      95042:data<=-16'd5325;
      95043:data<=16'd996;
      95044:data<=16'd4281;
      95045:data<=16'd1542;
      95046:data<=16'd206;
      95047:data<=16'd902;
      95048:data<=-16'd14;
      95049:data<=16'd4734;
      95050:data<=16'd13018;
      95051:data<=16'd13691;
      95052:data<=16'd12188;
      95053:data<=16'd13499;
      95054:data<=16'd12753;
      95055:data<=16'd11943;
      95056:data<=16'd12226;
      95057:data<=16'd11564;
      95058:data<=16'd10927;
      95059:data<=16'd9351;
      95060:data<=16'd8222;
      95061:data<=16'd8757;
      95062:data<=16'd7915;
      95063:data<=16'd7536;
      95064:data<=16'd8711;
      95065:data<=16'd8293;
      95066:data<=16'd7688;
      95067:data<=16'd7896;
      95068:data<=16'd7533;
      95069:data<=16'd7668;
      95070:data<=16'd8041;
      95071:data<=16'd6893;
      95072:data<=16'd4855;
      95073:data<=16'd4103;
      95074:data<=16'd4366;
      95075:data<=16'd3638;
      95076:data<=16'd3510;
      95077:data<=16'd4690;
      95078:data<=16'd4206;
      95079:data<=16'd3153;
      95080:data<=16'd3339;
      95081:data<=16'd2714;
      95082:data<=16'd2006;
      95083:data<=16'd2863;
      95084:data<=16'd2629;
      95085:data<=16'd399;
      95086:data<=-16'd519;
      95087:data<=-16'd214;
      95088:data<=-16'd713;
      95089:data<=-16'd303;
      95090:data<=16'd221;
      95091:data<=16'd56;
      95092:data<=16'd1657;
      95093:data<=-16'd644;
      95094:data<=-16'd8798;
      95095:data<=-16'd13244;
      95096:data<=-16'd16013;
      95097:data<=-16'd20901;
      95098:data<=-16'd20958;
      95099:data<=-16'd19511;
      95100:data<=-16'd20421;
      95101:data<=-16'd18650;
      95102:data<=-16'd17176;
      95103:data<=-16'd17356;
      95104:data<=-16'd15835;
      95105:data<=-16'd15192;
      95106:data<=-16'd14744;
      95107:data<=-16'd13521;
      95108:data<=-16'd13787;
      95109:data<=-16'd13056;
      95110:data<=-16'd11681;
      95111:data<=-16'd12091;
      95112:data<=-16'd12352;
      95113:data<=-16'd12352;
      95114:data<=-16'd12108;
      95115:data<=-16'd11059;
      95116:data<=-16'd10367;
      95117:data<=-16'd9583;
      95118:data<=-16'd9072;
      95119:data<=-16'd9027;
      95120:data<=-16'd8272;
      95121:data<=-16'd7859;
      95122:data<=-16'd7244;
      95123:data<=-16'd5987;
      95124:data<=-16'd6252;
      95125:data<=-16'd6905;
      95126:data<=-16'd6460;
      95127:data<=-16'd5918;
      95128:data<=-16'd5536;
      95129:data<=-16'd4796;
      95130:data<=-16'd3519;
      95131:data<=-16'd3168;
      95132:data<=-16'd3133;
      95133:data<=-16'd2308;
      95134:data<=-16'd3013;
      95135:data<=-16'd2359;
      95136:data<=-16'd338;
      95137:data<=-16'd2701;
      95138:data<=-16'd699;
      95139:data<=16'd8865;
      95140:data<=16'd11655;
      95141:data<=16'd9693;
      95142:data<=16'd10887;
      95143:data<=16'd10718;
      95144:data<=16'd10504;
      95145:data<=16'd11412;
      95146:data<=16'd10875;
      95147:data<=16'd10701;
      95148:data<=16'd10611;
      95149:data<=16'd13646;
      95150:data<=16'd19185;
      95151:data<=16'd17826;
      95152:data<=16'd14270;
      95153:data<=16'd15646;
      95154:data<=16'd15999;
      95155:data<=16'd15035;
      95156:data<=16'd14639;
      95157:data<=16'd13594;
      95158:data<=16'd14251;
      95159:data<=16'd14754;
      95160:data<=16'd13779;
      95161:data<=16'd13805;
      95162:data<=16'd13069;
      95163:data<=16'd12346;
      95164:data<=16'd13045;
      95165:data<=16'd12208;
      95166:data<=16'd11276;
      95167:data<=16'd11797;
      95168:data<=16'd11162;
      95169:data<=16'd10011;
      95170:data<=16'd9900;
      95171:data<=16'd9791;
      95172:data<=16'd9530;
      95173:data<=16'd9744;
      95174:data<=16'd9726;
      95175:data<=16'd9088;
      95176:data<=16'd8877;
      95177:data<=16'd9561;
      95178:data<=16'd10675;
      95179:data<=16'd10569;
      95180:data<=16'd9388;
      95181:data<=16'd10261;
      95182:data<=16'd9018;
      95183:data<=16'd1557;
      95184:data<=-16'd3336;
      95185:data<=-16'd3186;
      95186:data<=-16'd3791;
      95187:data<=-16'd2936;
      95188:data<=-16'd1830;
      95189:data<=-16'd2992;
      95190:data<=-16'd1814;
      95191:data<=-16'd70;
      95192:data<=-16'd77;
      95193:data<=16'd362;
      95194:data<=-16'd61;
      95195:data<=16'd18;
      95196:data<=16'd696;
      95197:data<=-16'd92;
      95198:data<=16'd505;
      95199:data<=16'd523;
      95200:data<=-16'd281;
      95201:data<=16'd1909;
      95202:data<=-16'd306;
      95203:data<=-16'd7050;
      95204:data<=-16'd7301;
      95205:data<=-16'd4545;
      95206:data<=-16'd4899;
      95207:data<=-16'd5095;
      95208:data<=-16'd4592;
      95209:data<=-16'd4067;
      95210:data<=-16'd3350;
      95211:data<=-16'd3069;
      95212:data<=-16'd2922;
      95213:data<=-16'd3125;
      95214:data<=-16'd2808;
      95215:data<=-16'd1501;
      95216:data<=-16'd1001;
      95217:data<=-16'd560;
      95218:data<=16'd1158;
      95219:data<=16'd1994;
      95220:data<=16'd876;
      95221:data<=16'd1099;
      95222:data<=16'd2689;
      95223:data<=16'd1413;
      95224:data<=16'd607;
      95225:data<=16'd2027;
      95226:data<=16'd382;
      95227:data<=16'd3087;
      95228:data<=16'd13195;
      95229:data<=16'd15910;
      95230:data<=16'd13345;
      95231:data<=16'd15471;
      95232:data<=16'd15738;
      95233:data<=16'd14101;
      95234:data<=16'd15206;
      95235:data<=16'd15226;
      95236:data<=16'd14158;
      95237:data<=16'd12948;
      95238:data<=16'd11555;
      95239:data<=16'd11872;
      95240:data<=16'd11785;
      95241:data<=16'd11045;
      95242:data<=16'd11075;
      95243:data<=16'd10821;
      95244:data<=16'd11706;
      95245:data<=16'd12539;
      95246:data<=16'd11762;
      95247:data<=16'd11902;
      95248:data<=16'd11585;
      95249:data<=16'd10780;
      95250:data<=16'd11306;
      95251:data<=16'd10759;
      95252:data<=16'd10489;
      95253:data<=16'd10520;
      95254:data<=16'd8387;
      95255:data<=16'd9975;
      95256:data<=16'd15388;
      95257:data<=16'd16789;
      95258:data<=16'd16443;
      95259:data<=16'd17306;
      95260:data<=16'd16211;
      95261:data<=16'd14784;
      95262:data<=16'd14613;
      95263:data<=16'd13761;
      95264:data<=16'd13509;
      95265:data<=16'd13981;
      95266:data<=16'd12501;
      95267:data<=16'd10909;
      95268:data<=16'd10687;
      95269:data<=16'd9821;
      95270:data<=16'd10692;
      95271:data<=16'd11800;
      95272:data<=16'd5564;
      95273:data<=-16'd2196;
      95274:data<=-16'd2704;
      95275:data<=-16'd2191;
      95276:data<=-16'd3322;
      95277:data<=-16'd2320;
      95278:data<=-16'd2299;
      95279:data<=-16'd3621;
      95280:data<=-16'd3445;
      95281:data<=-16'd3530;
      95282:data<=-16'd3566;
      95283:data<=-16'd2108;
      95284:data<=-16'd782;
      95285:data<=-16'd537;
      95286:data<=-16'd1165;
      95287:data<=-16'd1688;
      95288:data<=-16'd1365;
      95289:data<=-16'd1146;
      95290:data<=-16'd1375;
      95291:data<=-16'd1753;
      95292:data<=-16'd2135;
      95293:data<=-16'd2273;
      95294:data<=-16'd2551;
      95295:data<=-16'd2934;
      95296:data<=-16'd2922;
      95297:data<=-16'd1956;
      95298:data<=16'd20;
      95299:data<=16'd576;
      95300:data<=-16'd754;
      95301:data<=-16'd795;
      95302:data<=-16'd136;
      95303:data<=-16'd664;
      95304:data<=-16'd899;
      95305:data<=-16'd1274;
      95306:data<=-16'd1742;
      95307:data<=-16'd478;
      95308:data<=-16'd2378;
      95309:data<=-16'd9103;
      95310:data<=-16'd10572;
      95311:data<=-16'd6845;
      95312:data<=-16'd7494;
      95313:data<=-16'd8298;
      95314:data<=-16'd6505;
      95315:data<=-16'd8191;
      95316:data<=-16'd5877;
      95317:data<=16'd3554;
      95318:data<=16'd6652;
      95319:data<=16'd4329;
      95320:data<=16'd5118;
      95321:data<=16'd5247;
      95322:data<=16'd4276;
      95323:data<=16'd5084;
      95324:data<=16'd5799;
      95325:data<=16'd6313;
      95326:data<=16'd6076;
      95327:data<=16'd4793;
      95328:data<=16'd4431;
      95329:data<=16'd4084;
      95330:data<=16'd3447;
      95331:data<=16'd3568;
      95332:data<=16'd3600;
      95333:data<=16'd3318;
      95334:data<=16'd2601;
      95335:data<=16'd1807;
      95336:data<=16'd1783;
      95337:data<=16'd1985;
      95338:data<=16'd2767;
      95339:data<=16'd3553;
      95340:data<=16'd3248;
      95341:data<=16'd3052;
      95342:data<=16'd2475;
      95343:data<=16'd1659;
      95344:data<=16'd1939;
      95345:data<=16'd1363;
      95346:data<=16'd385;
      95347:data<=16'd725;
      95348:data<=16'd462;
      95349:data<=-16'd159;
      95350:data<=16'd652;
      95351:data<=16'd2171;
      95352:data<=16'd2353;
      95353:data<=16'd1155;
      95354:data<=16'd1460;
      95355:data<=16'd1895;
      95356:data<=16'd678;
      95357:data<=16'd1090;
      95358:data<=16'd1372;
      95359:data<=16'd470;
      95360:data<=16'd1086;
      95361:data<=-16'd1589;
      95362:data<=-16'd6169;
      95363:data<=-16'd5295;
      95364:data<=-16'd3457;
      95365:data<=-16'd3175;
      95366:data<=-16'd2187;
      95367:data<=-16'd3265;
      95368:data<=-16'd4367;
      95369:data<=-16'd3704;
      95370:data<=-16'd3944;
      95371:data<=-16'd3513;
      95372:data<=-16'd3063;
      95373:data<=-16'd3812;
      95374:data<=-16'd3333;
      95375:data<=-16'd3363;
      95376:data<=-16'd4458;
      95377:data<=-16'd4378;
      95378:data<=-16'd4649;
      95379:data<=-16'd5259;
      95380:data<=-16'd4755;
      95381:data<=-16'd4358;
      95382:data<=-16'd4498;
      95383:data<=-16'd4391;
      95384:data<=-16'd4282;
      95385:data<=-16'd4993;
      95386:data<=-16'd5385;
      95387:data<=-16'd4432;
      95388:data<=-16'd4303;
      95389:data<=-16'd5039;
      95390:data<=-16'd5169;
      95391:data<=-16'd5839;
      95392:data<=-16'd6338;
      95393:data<=-16'd5770;
      95394:data<=-16'd5630;
      95395:data<=-16'd5844;
      95396:data<=-16'd6117;
      95397:data<=-16'd6619;
      95398:data<=-16'd6733;
      95399:data<=-16'd6369;
      95400:data<=-16'd6313;
      95401:data<=-16'd6949;
      95402:data<=-16'd6457;
      95403:data<=-16'd6396;
      95404:data<=-16'd9254;
      95405:data<=-16'd7078;
      95406:data<=16'd1832;
      95407:data<=16'd5805;
      95408:data<=16'd4875;
      95409:data<=16'd4801;
      95410:data<=16'd3973;
      95411:data<=16'd3808;
      95412:data<=16'd4014;
      95413:data<=16'd3001;
      95414:data<=16'd2596;
      95415:data<=-16'd397;
      95416:data<=-16'd5063;
      95417:data<=-16'd6026;
      95418:data<=-16'd5994;
      95419:data<=-16'd6229;
      95420:data<=-16'd5662;
      95421:data<=-16'd5792;
      95422:data<=-16'd5463;
      95423:data<=-16'd5383;
      95424:data<=-16'd6009;
      95425:data<=-16'd5738;
      95426:data<=-16'd6431;
      95427:data<=-16'd6540;
      95428:data<=-16'd4993;
      95429:data<=-16'd5774;
      95430:data<=-16'd7339;
      95431:data<=-16'd7342;
      95432:data<=-16'd6939;
      95433:data<=-16'd6463;
      95434:data<=-16'd7147;
      95435:data<=-16'd7759;
      95436:data<=-16'd7292;
      95437:data<=-16'd7303;
      95438:data<=-16'd6657;
      95439:data<=-16'd6496;
      95440:data<=-16'd7056;
      95441:data<=-16'd5865;
      95442:data<=-16'd6047;
      95443:data<=-16'd7571;
      95444:data<=-16'd7985;
      95445:data<=-16'd8561;
      95446:data<=-16'd7260;
      95447:data<=-16'd6557;
      95448:data<=-16'd7982;
      95449:data<=-16'd6361;
      95450:data<=-16'd9162;
      95451:data<=-16'd18199;
      95452:data<=-16'd19946;
      95453:data<=-16'd17860;
      95454:data<=-16'd18836;
      95455:data<=-16'd17829;
      95456:data<=-16'd17397;
      95457:data<=-16'd19023;
      95458:data<=-16'd18779;
      95459:data<=-16'd18072;
      95460:data<=-16'd17051;
      95461:data<=-16'd15591;
      95462:data<=-16'd14968;
      95463:data<=-16'd14650;
      95464:data<=-16'd14625;
      95465:data<=-16'd13490;
      95466:data<=-16'd12475;
      95467:data<=-16'd12883;
      95468:data<=-16'd9793;
      95469:data<=-16'd5653;
      95470:data<=-16'd6096;
      95471:data<=-16'd6754;
      95472:data<=-16'd5899;
      95473:data<=-16'd5726;
      95474:data<=-16'd5297;
      95475:data<=-16'd5115;
      95476:data<=-16'd5197;
      95477:data<=-16'd4802;
      95478:data<=-16'd4046;
      95479:data<=-16'd2830;
      95480:data<=-16'd2825;
      95481:data<=-16'd3463;
      95482:data<=-16'd3362;
      95483:data<=-16'd4410;
      95484:data<=-16'd5369;
      95485:data<=-16'd4989;
      95486:data<=-16'd5143;
      95487:data<=-16'd5037;
      95488:data<=-16'd4358;
      95489:data<=-16'd3805;
      95490:data<=-16'd3140;
      95491:data<=-16'd2966;
      95492:data<=-16'd2713;
      95493:data<=-16'd2883;
      95494:data<=-16'd1883;
      95495:data<=16'd4702;
      95496:data<=16'd10619;
      95497:data<=16'd9608;
      95498:data<=16'd8636;
      95499:data<=16'd9621;
      95500:data<=16'd8805;
      95501:data<=16'd8502;
      95502:data<=16'd9086;
      95503:data<=16'd8980;
      95504:data<=16'd8937;
      95505:data<=16'd8379;
      95506:data<=16'd7420;
      95507:data<=16'd7332;
      95508:data<=16'd7685;
      95509:data<=16'd6795;
      95510:data<=16'd4773;
      95511:data<=16'd4432;
      95512:data<=16'd5184;
      95513:data<=16'd4830;
      95514:data<=16'd4919;
      95515:data<=16'd4814;
      95516:data<=16'd3839;
      95517:data<=16'd4340;
      95518:data<=16'd4543;
      95519:data<=16'd3833;
      95520:data<=16'd4481;
      95521:data<=16'd3175;
      95522:data<=-16'd1292;
      95523:data<=-16'd4149;
      95524:data<=-16'd4651;
      95525:data<=-16'd4987;
      95526:data<=-16'd4830;
      95527:data<=-16'd3915;
      95528:data<=-16'd3723;
      95529:data<=-16'd4212;
      95530:data<=-16'd3944;
      95531:data<=-16'd3295;
      95532:data<=-16'd2531;
      95533:data<=-16'd1794;
      95534:data<=-16'd1961;
      95535:data<=-16'd2208;
      95536:data<=-16'd3110;
      95537:data<=-16'd3824;
      95538:data<=-16'd1936;
      95539:data<=-16'd4466;
      95540:data<=-16'd13300;
      95541:data<=-16'd16597;
      95542:data<=-16'd14804;
      95543:data<=-16'd15382;
      95544:data<=-16'd14976;
      95545:data<=-16'd13417;
      95546:data<=-16'd13060;
      95547:data<=-16'd12102;
      95548:data<=-16'd11744;
      95549:data<=-16'd11970;
      95550:data<=-16'd11655;
      95551:data<=-16'd11653;
      95552:data<=-16'd10803;
      95553:data<=-16'd9947;
      95554:data<=-16'd10061;
      95555:data<=-16'd9567;
      95556:data<=-16'd9245;
      95557:data<=-16'd8596;
      95558:data<=-16'd7268;
      95559:data<=-16'd7069;
      95560:data<=-16'd6546;
      95561:data<=-16'd5940;
      95562:data<=-16'd6458;
      95563:data<=-16'd6244;
      95564:data<=-16'd6293;
      95565:data<=-16'd6608;
      95566:data<=-16'd5709;
      95567:data<=-16'd5351;
      95568:data<=-16'd4830;
      95569:data<=-16'd3926;
      95570:data<=-16'd4041;
      95571:data<=-16'd3142;
      95572:data<=-16'd2488;
      95573:data<=-16'd3145;
      95574:data<=-16'd854;
      95575:data<=16'd3089;
      95576:data<=16'd3886;
      95577:data<=16'd2726;
      95578:data<=16'd2966;
      95579:data<=16'd3755;
      95580:data<=16'd3139;
      95581:data<=16'd3712;
      95582:data<=16'd4596;
      95583:data<=16'd3453;
      95584:data<=16'd8094;
      95585:data<=16'd17089;
      95586:data<=16'd18048;
      95587:data<=16'd15753;
      95588:data<=16'd17026;
      95589:data<=16'd16553;
      95590:data<=16'd15890;
      95591:data<=16'd16480;
      95592:data<=16'd15013;
      95593:data<=16'd14659;
      95594:data<=16'd15396;
      95595:data<=16'd14277;
      95596:data<=16'd13712;
      95597:data<=16'd13746;
      95598:data<=16'd13295;
      95599:data<=16'd13373;
      95600:data<=16'd13103;
      95601:data<=16'd12703;
      95602:data<=16'd13408;
      95603:data<=16'd14239;
      95604:data<=16'd13960;
      95605:data<=16'd12944;
      95606:data<=16'd12663;
      95607:data<=16'd12803;
      95608:data<=16'd12298;
      95609:data<=16'd12037;
      95610:data<=16'd11905;
      95611:data<=16'd11555;
      95612:data<=16'd11594;
      95613:data<=16'd10865;
      95614:data<=16'd10041;
      95615:data<=16'd10939;
      95616:data<=16'd11379;
      95617:data<=16'd10837;
      95618:data<=16'd11309;
      95619:data<=16'd11341;
      95620:data<=16'd10775;
      95621:data<=16'd11376;
      95622:data<=16'd11174;
      95623:data<=16'd10178;
      95624:data<=16'd10454;
      95625:data<=16'd9879;
      95626:data<=16'd9009;
      95627:data<=16'd8445;
      95628:data<=16'd2247;
      95629:data<=-16'd6780;
      95630:data<=-16'd9520;
      95631:data<=-16'd9124;
      95632:data<=-16'd9829;
      95633:data<=-16'd9003;
      95634:data<=-16'd7890;
      95635:data<=-16'd8123;
      95636:data<=-16'd8144;
      95637:data<=-16'd7412;
      95638:data<=-16'd6463;
      95639:data<=-16'd6620;
      95640:data<=-16'd7024;
      95641:data<=-16'd5993;
      95642:data<=-16'd4545;
      95643:data<=-16'd2971;
      95644:data<=-16'd2194;
      95645:data<=-16'd2623;
      95646:data<=-16'd1988;
      95647:data<=-16'd1786;
      95648:data<=-16'd2534;
      95649:data<=-16'd1751;
      95650:data<=-16'd1589;
      95651:data<=-16'd2006;
      95652:data<=-16'd1171;
      95653:data<=-16'd1398;
      95654:data<=-16'd1583;
      95655:data<=-16'd335;
      95656:data<=16'd509;
      95657:data<=16'd1290;
      95658:data<=16'd1712;
      95659:data<=16'd1745;
      95660:data<=16'd1892;
      95661:data<=16'd1334;
      95662:data<=16'd1641;
      95663:data<=16'd2056;
      95664:data<=16'd1219;
      95665:data<=16'd1541;
      95666:data<=16'd1357;
      95667:data<=16'd546;
      95668:data<=16'd1619;
      95669:data<=16'd2246;
      95670:data<=16'd3745;
      95671:data<=16'd4965;
      95672:data<=16'd2449;
      95673:data<=16'd5938;
      95674:data<=16'd15517;
      95675:data<=16'd17183;
      95676:data<=16'd14681;
      95677:data<=16'd15822;
      95678:data<=16'd15622;
      95679:data<=16'd13925;
      95680:data<=16'd14904;
      95681:data<=16'd18269;
      95682:data<=16'd21158;
      95683:data<=16'd21026;
      95684:data<=16'd19590;
      95685:data<=16'd19073;
      95686:data<=16'd18692;
      95687:data<=16'd17984;
      95688:data<=16'd17048;
      95689:data<=16'd16407;
      95690:data<=16'd15716;
      95691:data<=16'd14592;
      95692:data<=16'd14252;
      95693:data<=16'd13298;
      95694:data<=16'd11759;
      95695:data<=16'd13016;
      95696:data<=16'd14533;
      95697:data<=16'd13358;
      95698:data<=16'd12531;
      95699:data<=16'd12668;
      95700:data<=16'd12167;
      95701:data<=16'd11441;
      95702:data<=16'd10712;
      95703:data<=16'd9906;
      95704:data<=16'd9263;
      95705:data<=16'd9003;
      95706:data<=16'd8523;
      95707:data<=16'd7511;
      95708:data<=16'd7632;
      95709:data<=16'd8857;
      95710:data<=16'd9166;
      95711:data<=16'd8445;
      95712:data<=16'd7705;
      95713:data<=16'd7533;
      95714:data<=16'd7127;
      95715:data<=16'd6328;
      95716:data<=16'd6449;
      95717:data<=16'd4206;
      95718:data<=-16'd2940;
      95719:data<=-16'd8816;
      95720:data<=-16'd9482;
      95721:data<=-16'd8040;
      95722:data<=-16'd6833;
      95723:data<=-16'd6592;
      95724:data<=-16'd6699;
      95725:data<=-16'd6106;
      95726:data<=-16'd5906;
      95727:data<=-16'd6296;
      95728:data<=-16'd5988;
      95729:data<=-16'd5462;
      95730:data<=-16'd5917;
      95731:data<=-16'd6328;
      95732:data<=-16'd5611;
      95733:data<=-16'd6296;
      95734:data<=-16'd8956;
      95735:data<=-16'd10105;
      95736:data<=-16'd10161;
      95737:data<=-16'd10317;
      95738:data<=-16'd9112;
      95739:data<=-16'd8422;
      95740:data<=-16'd9060;
      95741:data<=-16'd9021;
      95742:data<=-16'd9141;
      95743:data<=-16'd9159;
      95744:data<=-16'd8326;
      95745:data<=-16'd8349;
      95746:data<=-16'd8498;
      95747:data<=-16'd7756;
      95748:data<=-16'd6840;
      95749:data<=-16'd5621;
      95750:data<=-16'd4854;
      95751:data<=-16'd4808;
      95752:data<=-16'd4513;
      95753:data<=-16'd4193;
      95754:data<=-16'd4387;
      95755:data<=-16'd5072;
      95756:data<=-16'd4895;
      95757:data<=-16'd4340;
      95758:data<=-16'd5366;
      95759:data<=-16'd4940;
      95760:data<=-16'd3935;
      95761:data<=-16'd5601;
      95762:data<=-16'd1066;
      95763:data<=16'd9404;
      95764:data<=16'd11505;
      95765:data<=16'd9021;
      95766:data<=16'd10366;
      95767:data<=16'd9870;
      95768:data<=16'd8510;
      95769:data<=16'd9285;
      95770:data<=16'd8196;
      95771:data<=16'd7138;
      95772:data<=16'd7494;
      95773:data<=16'd6567;
      95774:data<=16'd6188;
      95775:data<=16'd7004;
      95776:data<=16'd7159;
      95777:data<=16'd6892;
      95778:data<=16'd6375;
      95779:data<=16'd5435;
      95780:data<=16'd4346;
      95781:data<=16'd3974;
      95782:data<=16'd4029;
      95783:data<=16'd3181;
      95784:data<=16'd3080;
      95785:data<=16'd3765;
      95786:data<=16'd3372;
      95787:data<=16'd5207;
      95788:data<=16'd9574;
      95789:data<=16'd11109;
      95790:data<=16'd10069;
      95791:data<=16'd9448;
      95792:data<=16'd8937;
      95793:data<=16'd8003;
      95794:data<=16'd7134;
      95795:data<=16'd7022;
      95796:data<=16'd6783;
      95797:data<=16'd5491;
      95798:data<=16'd4642;
      95799:data<=16'd4652;
      95800:data<=16'd4411;
      95801:data<=16'd3811;
      95802:data<=16'd3466;
      95803:data<=16'd3227;
      95804:data<=16'd1938;
      95805:data<=16'd1544;
      95806:data<=16'd2006;
      95807:data<=-16'd3471;
      95808:data<=-16'd11953;
      95809:data<=-16'd13423;
      95810:data<=-16'd11637;
      95811:data<=-16'd12087;
      95812:data<=-16'd11737;
      95813:data<=-16'd11389;
      95814:data<=-16'd12242;
      95815:data<=-16'd12313;
      95816:data<=-16'd12242;
      95817:data<=-16'd12334;
      95818:data<=-16'd12489;
      95819:data<=-16'd12851;
      95820:data<=-16'd12067;
      95821:data<=-16'd11122;
      95822:data<=-16'd11382;
      95823:data<=-16'd11330;
      95824:data<=-16'd10733;
      95825:data<=-16'd10671;
      95826:data<=-16'd10740;
      95827:data<=-16'd10486;
      95828:data<=-16'd10863;
      95829:data<=-16'd11870;
      95830:data<=-16'd11937;
      95831:data<=-16'd11696;
      95832:data<=-16'd11831;
      95833:data<=-16'd11091;
      95834:data<=-16'd10616;
      95835:data<=-16'd10819;
      95836:data<=-16'd10346;
      95837:data<=-16'd10746;
      95838:data<=-16'd11021;
      95839:data<=-16'd9292;
      95840:data<=-16'd10413;
      95841:data<=-16'd15393;
      95842:data<=-16'd17699;
      95843:data<=-16'd17027;
      95844:data<=-16'd17337;
      95845:data<=-16'd17030;
      95846:data<=-16'd15426;
      95847:data<=-16'd15215;
      95848:data<=-16'd14760;
      95849:data<=-16'd13841;
      95850:data<=-16'd14794;
      95851:data<=-16'd11359;
      95852:data<=-16'd1885;
      95853:data<=16'd2314;
      95854:data<=16'd320;
      95855:data<=-16'd143;
      95856:data<=-16'd347;
      95857:data<=-16'd1383;
      95858:data<=-16'd1175;
      95859:data<=-16'd807;
      95860:data<=-16'd687;
      95861:data<=-16'd957;
      95862:data<=-16'd1350;
      95863:data<=-16'd945;
      95864:data<=-16'd1127;
      95865:data<=-16'd1354;
      95866:data<=-16'd851;
      95867:data<=-16'd1838;
      95868:data<=-16'd3560;
      95869:data<=-16'd4259;
      95870:data<=-16'd4346;
      95871:data<=-16'd3805;
      95872:data<=-16'd3421;
      95873:data<=-16'd3497;
      95874:data<=-16'd3344;
      95875:data<=-16'd3113;
      95876:data<=-16'd2598;
      95877:data<=-16'd2440;
      95878:data<=-16'd2655;
      95879:data<=-16'd2121;
      95880:data<=-16'd2538;
      95881:data<=-16'd4026;
      95882:data<=-16'd4196;
      95883:data<=-16'd3717;
      95884:data<=-16'd3735;
      95885:data<=-16'd4358;
      95886:data<=-16'd4931;
      95887:data<=-16'd4200;
      95888:data<=-16'd3439;
      95889:data<=-16'd3206;
      95890:data<=-16'd2790;
      95891:data<=-16'd3149;
      95892:data<=-16'd3304;
      95893:data<=-16'd2046;
      95894:data<=16'd805;
      95895:data<=16'd3583;
      95896:data<=-16'd600;
      95897:data<=-16'd9829;
      95898:data<=-16'd12992;
      95899:data<=-16'd11658;
      95900:data<=-16'd11491;
      95901:data<=-16'd10287;
      95902:data<=-16'd9342;
      95903:data<=-16'd9962;
      95904:data<=-16'd9697;
      95905:data<=-16'd9106;
      95906:data<=-16'd8530;
      95907:data<=-16'd8379;
      95908:data<=-16'd9633;
      95909:data<=-16'd10016;
      95910:data<=-16'd9191;
      95911:data<=-16'd8787;
      95912:data<=-16'd8125;
      95913:data<=-16'd7412;
      95914:data<=-16'd7124;
      95915:data<=-16'd6748;
      95916:data<=-16'd6692;
      95917:data<=-16'd6648;
      95918:data<=-16'd5844;
      95919:data<=-16'd5015;
      95920:data<=-16'd5298;
      95921:data<=-16'd6313;
      95922:data<=-16'd6479;
      95923:data<=-16'd5938;
      95924:data<=-16'd5767;
      95925:data<=-16'd5497;
      95926:data<=-16'd5075;
      95927:data<=-16'd4837;
      95928:data<=-16'd4173;
      95929:data<=-16'd3609;
      95930:data<=-16'd3545;
      95931:data<=-16'd2819;
      95932:data<=-16'd2214;
      95933:data<=-16'd3008;
      95934:data<=-16'd3513;
      95935:data<=-16'd3530;
      95936:data<=-16'd4237;
      95937:data<=-16'd3682;
      95938:data<=-16'd2610;
      95939:data<=-16'd3336;
      95940:data<=-16'd819;
      95941:data<=16'd6930;
      95942:data<=16'd11914;
      95943:data<=16'd11430;
      95944:data<=16'd11054;
      95945:data<=16'd12013;
      95946:data<=16'd10079;
      95947:data<=16'd5130;
      95948:data<=16'd2126;
      95949:data<=16'd1679;
      95950:data<=16'd1384;
      95951:data<=16'd2030;
      95952:data<=16'd2799;
      95953:data<=16'd2634;
      95954:data<=16'd2969;
      95955:data<=16'd3083;
      95956:data<=16'd3171;
      95957:data<=16'd3570;
      95958:data<=16'd2878;
      95959:data<=16'd3213;
      95960:data<=16'd3680;
      95961:data<=16'd1691;
      95962:data<=16'd1431;
      95963:data<=16'd2537;
      95964:data<=16'd1674;
      95965:data<=16'd1923;
      95966:data<=16'd2651;
      95967:data<=16'd2046;
      95968:data<=16'd2591;
      95969:data<=16'd3080;
      95970:data<=16'd2522;
      95971:data<=16'd2529;
      95972:data<=16'd2684;
      95973:data<=16'd2455;
      95974:data<=16'd1463;
      95975:data<=16'd649;
      95976:data<=16'd937;
      95977:data<=16'd1104;
      95978:data<=16'd1886;
      95979:data<=16'd2362;
      95980:data<=16'd1612;
      95981:data<=16'd2593;
      95982:data<=16'd2523;
      95983:data<=16'd1128;
      95984:data<=16'd3139;
      95985:data<=16'd506;
      95986:data<=-16'd9182;
      95987:data<=-16'd13003;
      95988:data<=-16'd11728;
      95989:data<=-16'd12289;
      95990:data<=-16'd11492;
      95991:data<=-16'd10140;
      95992:data<=-16'd10216;
      95993:data<=-16'd9113;
      95994:data<=-16'd8099;
      95995:data<=-16'd8213;
      95996:data<=-16'd7412;
      95997:data<=-16'd6593;
      95998:data<=-16'd6824;
      95999:data<=-16'd5303;
      96000:data<=-16'd1607;
      96001:data<=16'd96;
      96002:data<=16'd109;
      96003:data<=16'd1213;
      96004:data<=16'd1274;
      96005:data<=16'd270;
      96006:data<=16'd467;
      96007:data<=16'd749;
      96008:data<=16'd930;
      96009:data<=16'd951;
      96010:data<=16'd481;
      96011:data<=16'd1127;
      96012:data<=16'd1953;
      96013:data<=16'd2032;
      96014:data<=16'd2211;
      96015:data<=16'd1889;
      96016:data<=16'd2215;
      96017:data<=16'd3283;
      96018:data<=16'd2952;
      96019:data<=16'd2364;
      96020:data<=16'd2364;
      96021:data<=16'd2508;
      96022:data<=16'd2846;
      96023:data<=16'd2863;
      96024:data<=16'd3412;
      96025:data<=16'd3513;
      96026:data<=16'd3186;
      96027:data<=16'd5318;
      96028:data<=16'd5841;
      96029:data<=16'd5410;
      96030:data<=16'd12283;
      96031:data<=16'd19388;
      96032:data<=16'd18907;
      96033:data<=16'd18107;
      96034:data<=16'd18383;
      96035:data<=16'd17059;
      96036:data<=16'd16953;
      96037:data<=16'd17054;
      96038:data<=16'd15719;
      96039:data<=16'd14930;
      96040:data<=16'd15565;
      96041:data<=16'd16533;
      96042:data<=16'd16304;
      96043:data<=16'd15769;
      96044:data<=16'd15822;
      96045:data<=16'd15420;
      96046:data<=16'd14737;
      96047:data<=16'd13746;
      96048:data<=16'd13129;
      96049:data<=16'd13402;
      96050:data<=16'd12830;
      96051:data<=16'd12706;
      96052:data<=16'd12228;
      96053:data<=16'd8420;
      96054:data<=16'd6087;
      96055:data<=16'd6840;
      96056:data<=16'd6401;
      96057:data<=16'd6032;
      96058:data<=16'd6220;
      96059:data<=16'd6147;
      96060:data<=16'd6663;
      96061:data<=16'd5903;
      96062:data<=16'd5225;
      96063:data<=16'd6273;
      96064:data<=16'd6169;
      96065:data<=16'd5498;
      96066:data<=16'd5850;
      96067:data<=16'd6704;
      96068:data<=16'd7169;
      96069:data<=16'd6766;
      96070:data<=16'd7733;
      96071:data<=16'd7820;
      96072:data<=16'd5947;
      96073:data<=16'd7409;
      96074:data<=16'd5059;
      96075:data<=-16'd4810;
      96076:data<=-16'd8150;
      96077:data<=-16'd6281;
      96078:data<=-16'd7876;
      96079:data<=-16'd7304;
      96080:data<=-16'd5109;
      96081:data<=-16'd4684;
      96082:data<=-16'd3594;
      96083:data<=-16'd3265;
      96084:data<=-16'd2984;
      96085:data<=-16'd2344;
      96086:data<=-16'd3310;
      96087:data<=-16'd3192;
      96088:data<=-16'd2766;
      96089:data<=-16'd3353;
      96090:data<=-16'd2684;
      96091:data<=-16'd2640;
      96092:data<=-16'd2877;
      96093:data<=-16'd1686;
      96094:data<=-16'd1017;
      96095:data<=-16'd378;
      96096:data<=-16'd56;
      96097:data<=-16'd246;
      96098:data<=16'd264;
      96099:data<=-16'd405;
      96100:data<=-16'd528;
      96101:data<=16'd588;
      96102:data<=-16'd334;
      96103:data<=-16'd202;
      96104:data<=16'd696;
      96105:data<=-16'd331;
      96106:data<=16'd2604;
      96107:data<=16'd7967;
      96108:data<=16'd8514;
      96109:data<=16'd7426;
      96110:data<=16'd8091;
      96111:data<=16'd7882;
      96112:data<=16'd6290;
      96113:data<=16'd6140;
      96114:data<=16'd6590;
      96115:data<=16'd4837;
      96116:data<=16'd4871;
      96117:data<=16'd6219;
      96118:data<=16'd4557;
      96119:data<=16'd8840;
      96120:data<=16'd19026;
      96121:data<=16'd20835;
      96122:data<=16'd18246;
      96123:data<=16'd19068;
      96124:data<=16'd18016;
      96125:data<=16'd15952;
      96126:data<=16'd15529;
      96127:data<=16'd14542;
      96128:data<=16'd13809;
      96129:data<=16'd13453;
      96130:data<=16'd13042;
      96131:data<=16'd12730;
      96132:data<=16'd12116;
      96133:data<=16'd12912;
      96134:data<=16'd13770;
      96135:data<=16'd12389;
      96136:data<=16'd11467;
      96137:data<=16'd11351;
      96138:data<=16'd10443;
      96139:data<=16'd9768;
      96140:data<=16'd9257;
      96141:data<=16'd8479;
      96142:data<=16'd8006;
      96143:data<=16'd8000;
      96144:data<=16'd7917;
      96145:data<=16'd7054;
      96146:data<=16'd6855;
      96147:data<=16'd7965;
      96148:data<=16'd8038;
      96149:data<=16'd7078;
      96150:data<=16'd6614;
      96151:data<=16'd6391;
      96152:data<=16'd6344;
      96153:data<=16'd6197;
      96154:data<=16'd5338;
      96155:data<=16'd4460;
      96156:data<=16'd4346;
      96157:data<=16'd4473;
      96158:data<=16'd4093;
      96159:data<=16'd2591;
      96160:data<=-16'd522;
      96161:data<=-16'd2205;
      96162:data<=-16'd714;
      96163:data<=-16'd3327;
      96164:data<=-16'd11565;
      96165:data<=-16'd15209;
      96166:data<=-16'd13638;
      96167:data<=-16'd13679;
      96168:data<=-16'd14064;
      96169:data<=-16'd13477;
      96170:data<=-16'd13553;
      96171:data<=-16'd13309;
      96172:data<=-16'd12425;
      96173:data<=-16'd11356;
      96174:data<=-16'd10184;
      96175:data<=-16'd9454;
      96176:data<=-16'd9150;
      96177:data<=-16'd9315;
      96178:data<=-16'd9612;
      96179:data<=-16'd9482;
      96180:data<=-16'd8980;
      96181:data<=-16'd7971;
      96182:data<=-16'd7771;
      96183:data<=-16'd8853;
      96184:data<=-16'd8960;
      96185:data<=-16'd8252;
      96186:data<=-16'd7676;
      96187:data<=-16'd6567;
      96188:data<=-16'd5883;
      96189:data<=-16'd5809;
      96190:data<=-16'd5363;
      96191:data<=-16'd5330;
      96192:data<=-16'd5902;
      96193:data<=-16'd5976;
      96194:data<=-16'd5356;
      96195:data<=-16'd5345;
      96196:data<=-16'd6229;
      96197:data<=-16'd6445;
      96198:data<=-16'd6296;
      96199:data<=-16'd5715;
      96200:data<=-16'd3988;
      96201:data<=-16'd3792;
      96202:data<=-16'd4215;
      96203:data<=-16'd3051;
      96204:data<=-16'd3612;
      96205:data<=-16'd4109;
      96206:data<=-16'd2984;
      96207:data<=-16'd4337;
      96208:data<=-16'd1350;
      96209:data<=16'd8537;
      96210:data<=16'd11018;
      96211:data<=16'd7101;
      96212:data<=16'd9859;
      96213:data<=16'd15003;
      96214:data<=16'd15493;
      96215:data<=16'd14678;
      96216:data<=16'd13987;
      96217:data<=16'd12889;
      96218:data<=16'd12192;
      96219:data<=16'd11292;
      96220:data<=16'd10328;
      96221:data<=16'd10073;
      96222:data<=16'd9729;
      96223:data<=16'd9104;
      96224:data<=16'd8616;
      96225:data<=16'd7802;
      96226:data<=16'd7125;
      96227:data<=16'd6965;
      96228:data<=16'd6291;
      96229:data<=16'd5630;
      96230:data<=16'd5636;
      96231:data<=16'd5194;
      96232:data<=16'd4620;
      96233:data<=16'd4394;
      96234:data<=16'd3591;
      96235:data<=16'd2567;
      96236:data<=16'd2232;
      96237:data<=16'd2567;
      96238:data<=16'd2637;
      96239:data<=16'd1701;
      96240:data<=16'd675;
      96241:data<=-16'd149;
      96242:data<=-16'd779;
      96243:data<=-16'd654;
      96244:data<=-16'd1068;
      96245:data<=-16'd1689;
      96246:data<=-16'd1239;
      96247:data<=-16'd1374;
      96248:data<=-16'd1556;
      96249:data<=-16'd1536;
      96250:data<=-16'd2623;
      96251:data<=-16'd2049;
      96252:data<=-16'd3169;
      96253:data<=-16'd11603;
      96254:data<=-16'd18357;
      96255:data<=-16'd17540;
      96256:data<=-16'd16821;
      96257:data<=-16'd17320;
      96258:data<=-16'd15916;
      96259:data<=-16'd15374;
      96260:data<=-16'd15719;
      96261:data<=-16'd14865;
      96262:data<=-16'd14305;
      96263:data<=-16'd13803;
      96264:data<=-16'd12566;
      96265:data<=-16'd14615;
      96266:data<=-16'd19920;
      96267:data<=-16'd21782;
      96268:data<=-16'd20624;
      96269:data<=-16'd20604;
      96270:data<=-16'd19735;
      96271:data<=-16'd18280;
      96272:data<=-16'd18098;
      96273:data<=-16'd17438;
      96274:data<=-16'd16971;
      96275:data<=-16'd16862;
      96276:data<=-16'd15775;
      96277:data<=-16'd15032;
      96278:data<=-16'd14424;
      96279:data<=-16'd14263;
      96280:data<=-16'd15344;
      96281:data<=-16'd15335;
      96282:data<=-16'd14929;
      96283:data<=-16'd15044;
      96284:data<=-16'd14102;
      96285:data<=-16'd13471;
      96286:data<=-16'd13132;
      96287:data<=-16'd12404;
      96288:data<=-16'd12392;
      96289:data<=-16'd12116;
      96290:data<=-16'd11991;
      96291:data<=-16'd11711;
      96292:data<=-16'd11166;
      96293:data<=-16'd13012;
      96294:data<=-16'd12569;
      96295:data<=-16'd10094;
      96296:data<=-16'd12622;
      96297:data<=-16'd9781;
      96298:data<=16'd1533;
      96299:data<=16'd4726;
      96300:data<=16'd2247;
      96301:data<=16'd3427;
      96302:data<=16'd2943;
      96303:data<=16'd1917;
      96304:data<=16'd3068;
      96305:data<=16'd2478;
      96306:data<=16'd1104;
      96307:data<=16'd293;
      96308:data<=-16'd197;
      96309:data<=16'd412;
      96310:data<=16'd890;
      96311:data<=16'd795;
      96312:data<=16'd455;
      96313:data<=16'd326;
      96314:data<=16'd1036;
      96315:data<=16'd993;
      96316:data<=16'd20;
      96317:data<=-16'd582;
      96318:data<=16'd287;
      96319:data<=16'd3506;
      96320:data<=16'd5410;
      96321:data<=16'd4411;
      96322:data<=16'd4361;
      96323:data<=16'd4704;
      96324:data<=16'd4175;
      96325:data<=16'd4202;
      96326:data<=16'd4131;
      96327:data<=16'd4123;
      96328:data<=16'd4255;
      96329:data<=16'd3971;
      96330:data<=16'd3900;
      96331:data<=16'd3142;
      96332:data<=16'd2253;
      96333:data<=16'd2094;
      96334:data<=16'd1565;
      96335:data<=16'd1721;
      96336:data<=16'd1780;
      96337:data<=16'd1263;
      96338:data<=16'd1992;
      96339:data<=16'd1140;
      96340:data<=16'd346;
      96341:data<=16'd1902;
      96342:data<=-16'd2616;
      96343:data<=-16'd10768;
      96344:data<=-16'd11825;
      96345:data<=-16'd10854;
      96346:data<=-16'd12587;
      96347:data<=-16'd12516;
      96348:data<=-16'd11304;
      96349:data<=-16'd10725;
      96350:data<=-16'd10003;
      96351:data<=-16'd9767;
      96352:data<=-16'd9726;
      96353:data<=-16'd8880;
      96354:data<=-16'd7897;
      96355:data<=-16'd7941;
      96356:data<=-16'd7971;
      96357:data<=-16'd7047;
      96358:data<=-16'd7021;
      96359:data<=-16'd7830;
      96360:data<=-16'd7903;
      96361:data<=-16'd7591;
      96362:data<=-16'd7042;
      96363:data<=-16'd6667;
      96364:data<=-16'd6446;
      96365:data<=-16'd5759;
      96366:data<=-16'd5375;
      96367:data<=-16'd4907;
      96368:data<=-16'd4722;
      96369:data<=-16'd5139;
      96370:data<=-16'd3876;
      96371:data<=-16'd4068;
      96372:data<=-16'd8548;
      96373:data<=-16'd11741;
      96374:data<=-16'd11756;
      96375:data<=-16'd11450;
      96376:data<=-16'd11088;
      96377:data<=-16'd10147;
      96378:data<=-16'd8831;
      96379:data<=-16'd8940;
      96380:data<=-16'd9189;
      96381:data<=-16'd7668;
      96382:data<=-16'd7735;
      96383:data<=-16'd7109;
      96384:data<=-16'd4971;
      96385:data<=-16'd7365;
      96386:data<=-16'd6102;
      96387:data<=16'd3330;
      96388:data<=16'd7043;
      96389:data<=16'd5338;
      96390:data<=16'd6507;
      96391:data<=16'd6937;
      96392:data<=16'd6354;
      96393:data<=16'd6590;
      96394:data<=16'd6467;
      96395:data<=16'd6843;
      96396:data<=16'd6716;
      96397:data<=16'd6222;
      96398:data<=16'd5968;
      96399:data<=16'd4437;
      96400:data<=16'd3738;
      96401:data<=16'd4282;
      96402:data<=16'd4302;
      96403:data<=16'd4764;
      96404:data<=16'd4531;
      96405:data<=16'd3629;
      96406:data<=16'd3758;
      96407:data<=16'd3748;
      96408:data<=16'd3990;
      96409:data<=16'd4485;
      96410:data<=16'd4140;
      96411:data<=16'd3902;
      96412:data<=16'd3284;
      96413:data<=16'd2851;
      96414:data<=16'd3560;
      96415:data<=16'd3633;
      96416:data<=16'd3562;
      96417:data<=16'd3532;
      96418:data<=16'd2949;
      96419:data<=16'd3442;
      96420:data<=16'd3993;
      96421:data<=16'd4181;
      96422:data<=16'd4751;
      96423:data<=16'd3990;
      96424:data<=16'd3785;
      96425:data<=16'd5839;
      96426:data<=16'd8257;
      96427:data<=16'd9909;
      96428:data<=16'd8772;
      96429:data<=16'd7988;
      96430:data<=16'd10041;
      96431:data<=16'd5785;
      96432:data<=-16'd3542;
      96433:data<=-16'd5676;
      96434:data<=-16'd3422;
      96435:data<=-16'd3201;
      96436:data<=-16'd3250;
      96437:data<=-16'd3660;
      96438:data<=-16'd3494;
      96439:data<=-16'd1806;
      96440:data<=-16'd1632;
      96441:data<=-16'd2305;
      96442:data<=-16'd1601;
      96443:data<=-16'd1068;
      96444:data<=-16'd1192;
      96445:data<=-16'd755;
      96446:data<=-16'd579;
      96447:data<=-16'd1254;
      96448:data<=-16'd905;
      96449:data<=16'd347;
      96450:data<=16'd667;
      96451:data<=16'd1307;
      96452:data<=16'd2714;
      96453:data<=16'd3115;
      96454:data<=16'd3196;
      96455:data<=16'd3624;
      96456:data<=16'd3435;
      96457:data<=16'd3001;
      96458:data<=16'd3228;
      96459:data<=16'd3768;
      96460:data<=16'd3621;
      96461:data<=16'd3319;
      96462:data<=16'd3657;
      96463:data<=16'd3656;
      96464:data<=16'd3990;
      96465:data<=16'd5359;
      96466:data<=16'd5821;
      96467:data<=16'd5577;
      96468:data<=16'd5718;
      96469:data<=16'd5835;
      96470:data<=16'd5968;
      96471:data<=16'd5462;
      96472:data<=16'd5247;
      96473:data<=16'd6081;
      96474:data<=16'd5369;
      96475:data<=16'd6366;
      96476:data<=16'd13409;
      96477:data<=16'd19103;
      96478:data<=16'd17223;
      96479:data<=16'd12968;
      96480:data<=16'd11588;
      96481:data<=16'd12126;
      96482:data<=16'd12108;
      96483:data<=16'd11608;
      96484:data<=16'd11059;
      96485:data<=16'd10175;
      96486:data<=16'd10342;
      96487:data<=16'd10995;
      96488:data<=16'd10087;
      96489:data<=16'd9183;
      96490:data<=16'd9401;
      96491:data<=16'd9952;
      96492:data<=16'd10722;
      96493:data<=16'd10812;
      96494:data<=16'd10117;
      96495:data<=16'd9394;
      96496:data<=16'd8904;
      96497:data<=16'd9294;
      96498:data<=16'd9283;
      96499:data<=16'd8260;
      96500:data<=16'd8616;
      96501:data<=16'd9514;
      96502:data<=16'd8617;
      96503:data<=16'd7503;
      96504:data<=16'd8040;
      96505:data<=16'd9256;
      96506:data<=16'd9297;
      96507:data<=16'd8640;
      96508:data<=16'd8439;
      96509:data<=16'd8156;
      96510:data<=16'd8290;
      96511:data<=16'd8275;
      96512:data<=16'd6884;
      96513:data<=16'd6479;
      96514:data<=16'd6728;
      96515:data<=16'd6050;
      96516:data<=16'd6581;
      96517:data<=16'd6613;
      96518:data<=16'd6194;
      96519:data<=16'd8279;
      96520:data<=16'd5295;
      96521:data<=-16'd4297;
      96522:data<=-16'd7712;
      96523:data<=-16'd5559;
      96524:data<=-16'd6478;
      96525:data<=-16'd6713;
      96526:data<=-16'd4902;
      96527:data<=-16'd5221;
      96528:data<=-16'd5195;
      96529:data<=-16'd4472;
      96530:data<=-16'd5274;
      96531:data<=-16'd2919;
      96532:data<=16'd2722;
      96533:data<=16'd4434;
      96534:data<=16'd3459;
      96535:data<=16'd4200;
      96536:data<=16'd4040;
      96537:data<=16'd2842;
      96538:data<=16'd3168;
      96539:data<=16'd3592;
      96540:data<=16'd3748;
      96541:data<=16'd4059;
      96542:data<=16'd3196;
      96543:data<=16'd2334;
      96544:data<=16'd3093;
      96545:data<=16'd4269;
      96546:data<=16'd4228;
      96547:data<=16'd3325;
      96548:data<=16'd3342;
      96549:data<=16'd3506;
      96550:data<=16'd2669;
      96551:data<=16'd2746;
      96552:data<=16'd3018;
      96553:data<=16'd2082;
      96554:data<=16'd1932;
      96555:data<=16'd1867;
      96556:data<=16'd1137;
      96557:data<=16'd1695;
      96558:data<=16'd2654;
      96559:data<=16'd3052;
      96560:data<=16'd2916;
      96561:data<=16'd2035;
      96562:data<=16'd2132;
      96563:data<=16'd2096;
      96564:data<=16'd2265;
      96565:data<=16'd7859;
      96566:data<=16'd14499;
      96567:data<=16'd14795;
      96568:data<=16'd13300;
      96569:data<=16'd13262;
      96570:data<=16'd12515;
      96571:data<=16'd12474;
      96572:data<=16'd12821;
      96573:data<=16'd11840;
      96574:data<=16'd11341;
      96575:data<=16'd11245;
      96576:data<=16'd10241;
      96577:data<=16'd9861;
      96578:data<=16'd9826;
      96579:data<=16'd8334;
      96580:data<=16'd7303;
      96581:data<=16'd7483;
      96582:data<=16'd6766;
      96583:data<=16'd6202;
      96584:data<=16'd5068;
      96585:data<=16'd1245;
      96586:data<=-16'd846;
      96587:data<=16'd52;
      96588:data<=-16'd8;
      96589:data<=16'd65;
      96590:data<=16'd582;
      96591:data<=16'd203;
      96592:data<=16'd161;
      96593:data<=-16'd277;
      96594:data<=-16'd729;
      96595:data<=-16'd610;
      96596:data<=-16'd1245;
      96597:data<=-16'd625;
      96598:data<=16'd514;
      96599:data<=16'd138;
      96600:data<=16'd602;
      96601:data<=16'd657;
      96602:data<=-16'd55;
      96603:data<=16'd385;
      96604:data<=-16'd156;
      96605:data<=-16'd375;
      96606:data<=16'd77;
      96607:data<=-16'd256;
      96608:data<=16'd963;
      96609:data<=-16'd2566;
      96610:data<=-16'd11822;
      96611:data<=-16'd13621;
      96612:data<=-16'd10662;
      96613:data<=-16'd11468;
      96614:data<=-16'd11412;
      96615:data<=-16'd10698;
      96616:data<=-16'd10965;
      96617:data<=-16'd10096;
      96618:data<=-16'd10325;
      96619:data<=-16'd10866;
      96620:data<=-16'd10232;
      96621:data<=-16'd10070;
      96622:data<=-16'd9726;
      96623:data<=-16'd9116;
      96624:data<=-16'd7962;
      96625:data<=-16'd6593;
      96626:data<=-16'd6719;
      96627:data<=-16'd6379;
      96628:data<=-16'd5604;
      96629:data<=-16'd5789;
      96630:data<=-16'd5371;
      96631:data<=-16'd5288;
      96632:data<=-16'd5460;
      96633:data<=-16'd5145;
      96634:data<=-16'd5779;
      96635:data<=-16'd6073;
      96636:data<=-16'd6108;
      96637:data<=-16'd4589;
      96638:data<=16'd687;
      96639:data<=16'd3389;
      96640:data<=16'd2347;
      96641:data<=16'd2538;
      96642:data<=16'd2126;
      96643:data<=16'd1897;
      96644:data<=16'd2447;
      96645:data<=16'd1325;
      96646:data<=16'd1154;
      96647:data<=16'd745;
      96648:data<=-16'd367;
      96649:data<=16'd544;
      96650:data<=-16'd197;
      96651:data<=-16'd429;
      96652:data<=16'd681;
      96653:data<=-16'd2029;
      96654:data<=16'd1039;
      96655:data<=16'd10939;
      96656:data<=16'd12489;
      96657:data<=16'd9523;
      96658:data<=16'd10166;
      96659:data<=16'd10093;
      96660:data<=16'd9324;
      96661:data<=16'd8748;
      96662:data<=16'd7993;
      96663:data<=16'd7615;
      96664:data<=16'd5786;
      96665:data<=16'd4422;
      96666:data<=16'd4373;
      96667:data<=16'd3275;
      96668:data<=16'd2908;
      96669:data<=16'd3198;
      96670:data<=16'd2928;
      96671:data<=16'd2904;
      96672:data<=16'd2091;
      96673:data<=16'd1583;
      96674:data<=16'd1836;
      96675:data<=16'd1087;
      96676:data<=16'd691;
      96677:data<=16'd82;
      96678:data<=-16'd1460;
      96679:data<=-16'd1739;
      96680:data<=-16'd1897;
      96681:data<=-16'd2387;
      96682:data<=-16'd1756;
      96683:data<=-16'd1234;
      96684:data<=-16'd1512;
      96685:data<=-16'd2161;
      96686:data<=-16'd2391;
      96687:data<=-16'd2040;
      96688:data<=-16'd2091;
      96689:data<=-16'd1989;
      96690:data<=-16'd3538;
      96691:data<=-16'd8049;
      96692:data<=-16'd10795;
      96693:data<=-16'd10624;
      96694:data<=-16'd10273;
      96695:data<=-16'd10055;
      96696:data<=-16'd9770;
      96697:data<=-16'd8422;
      96698:data<=-16'd9734;
      96699:data<=-16'd17126;
      96700:data<=-16'd21910;
      96701:data<=-16'd20342;
      96702:data<=-16'd19167;
      96703:data<=-16'd19182;
      96704:data<=-16'd19669;
      96705:data<=-16'd20407;
      96706:data<=-16'd19200;
      96707:data<=-16'd18515;
      96708:data<=-16'd18534;
      96709:data<=-16'd17123;
      96710:data<=-16'd16795;
      96711:data<=-16'd16583;
      96712:data<=-16'd15132;
      96713:data<=-16'd14974;
      96714:data<=-16'd14759;
      96715:data<=-16'd13778;
      96716:data<=-16'd13670;
      96717:data<=-16'd13486;
      96718:data<=-16'd13471;
      96719:data<=-16'd13737;
      96720:data<=-16'd13063;
      96721:data<=-16'd12214;
      96722:data<=-16'd11491;
      96723:data<=-16'd11089;
      96724:data<=-16'd11630;
      96725:data<=-16'd11784;
      96726:data<=-16'd11144;
      96727:data<=-16'd10807;
      96728:data<=-16'd10572;
      96729:data<=-16'd9966;
      96730:data<=-16'd9890;
      96731:data<=-16'd10605;
      96732:data<=-16'd10317;
      96733:data<=-16'd9388;
      96734:data<=-16'd9351;
      96735:data<=-16'd8846;
      96736:data<=-16'd8422;
      96737:data<=-16'd8783;
      96738:data<=-16'd8214;
      96739:data<=-16'd8062;
      96740:data<=-16'd7585;
      96741:data<=-16'd6258;
      96742:data<=-16'd7732;
      96743:data<=-16'd5137;
      96744:data<=16'd5844;
      96745:data<=16'd12216;
      96746:data<=16'd11303;
      96747:data<=16'd11191;
      96748:data<=16'd10680;
      96749:data<=16'd9855;
      96750:data<=16'd10245;
      96751:data<=16'd9480;
      96752:data<=16'd8836;
      96753:data<=16'd8625;
      96754:data<=16'd8090;
      96755:data<=16'd8123;
      96756:data<=16'd6898;
      96757:data<=16'd5201;
      96758:data<=16'd4687;
      96759:data<=16'd3940;
      96760:data<=16'd4117;
      96761:data<=16'd4466;
      96762:data<=16'd3290;
      96763:data<=16'd3109;
      96764:data<=16'd3441;
      96765:data<=16'd3254;
      96766:data<=16'd3653;
      96767:data<=16'd3272;
      96768:data<=16'd3113;
      96769:data<=16'd3974;
      96770:data<=16'd2981;
      96771:data<=16'd1406;
      96772:data<=16'd1375;
      96773:data<=16'd1278;
      96774:data<=16'd1060;
      96775:data<=16'd1542;
      96776:data<=16'd1838;
      96777:data<=16'd1562;
      96778:data<=16'd1718;
      96779:data<=16'd2249;
      96780:data<=16'd2185;
      96781:data<=16'd2278;
      96782:data<=16'd2472;
      96783:data<=16'd1629;
      96784:data<=16'd253;
      96785:data<=-16'd975;
      96786:data<=-16'd719;
      96787:data<=-16'd1037;
      96788:data<=-16'd7004;
      96789:data<=-16'd13347;
      96790:data<=-16'd13251;
      96791:data<=-16'd11800;
      96792:data<=-16'd11515;
      96793:data<=-16'd10499;
      96794:data<=-16'd10484;
      96795:data<=-16'd10084;
      96796:data<=-16'd9315;
      96797:data<=-16'd12477;
      96798:data<=-16'd16860;
      96799:data<=-16'd17424;
      96800:data<=-16'd15834;
      96801:data<=-16'd14678;
      96802:data<=-16'd13725;
      96803:data<=-16'd12868;
      96804:data<=-16'd12248;
      96805:data<=-16'd11435;
      96806:data<=-16'd10947;
      96807:data<=-16'd10499;
      96808:data<=-16'd8997;
      96809:data<=-16'd8698;
      96810:data<=-16'd10398;
      96811:data<=-16'd10592;
      96812:data<=-16'd9362;
      96813:data<=-16'd9222;
      96814:data<=-16'd9524;
      96815:data<=-16'd8846;
      96816:data<=-16'd7721;
      96817:data<=-16'd7410;
      96818:data<=-16'd6998;
      96819:data<=-16'd6005;
      96820:data<=-16'd5894;
      96821:data<=-16'd5788;
      96822:data<=-16'd5650;
      96823:data<=-16'd6115;
      96824:data<=-16'd5650;
      96825:data<=-16'd5973;
      96826:data<=-16'd6672;
      96827:data<=-16'd5072;
      96828:data<=-16'd4434;
      96829:data<=-16'd4131;
      96830:data<=-16'd3338;
      96831:data<=-16'd5115;
      96832:data<=-16'd1353;
      96833:data<=16'd8757;
      96834:data<=16'd11617;
      96835:data<=16'd9740;
      96836:data<=16'd10006;
      96837:data<=16'd8733;
      96838:data<=16'd8231;
      96839:data<=16'd9012;
      96840:data<=16'd7577;
      96841:data<=16'd7480;
      96842:data<=16'd8602;
      96843:data<=16'd7800;
      96844:data<=16'd7007;
      96845:data<=16'd6695;
      96846:data<=16'd6432;
      96847:data<=16'd7021;
      96848:data<=16'd7127;
      96849:data<=16'd5768;
      96850:data<=16'd6029;
      96851:data<=16'd10029;
      96852:data<=16'd12622;
      96853:data<=16'd11122;
      96854:data<=16'd10608;
      96855:data<=16'd11324;
      96856:data<=16'd10643;
      96857:data<=16'd10110;
      96858:data<=16'd9835;
      96859:data<=16'd9864;
      96860:data<=16'd10516;
      96861:data<=16'd10334;
      96862:data<=16'd10011;
      96863:data<=16'd10003;
      96864:data<=16'd9847;
      96865:data<=16'd9752;
      96866:data<=16'd9230;
      96867:data<=16'd9429;
      96868:data<=16'd9464;
      96869:data<=16'd7840;
      96870:data<=16'd8032;
      96871:data<=16'd9065;
      96872:data<=16'd8396;
      96873:data<=16'd8514;
      96874:data<=16'd7838;
      96875:data<=16'd7238;
      96876:data<=16'd9009;
      96877:data<=16'd5412;
      96878:data<=-16'd2714;
      96879:data<=-16'd4757;
      96880:data<=-16'd3096;
      96881:data<=-16'd3298;
      96882:data<=-16'd3095;
      96883:data<=-16'd2088;
      96884:data<=-16'd1691;
      96885:data<=-16'd1436;
      96886:data<=-16'd974;
      96887:data<=-16'd1031;
      96888:data<=-16'd1583;
      96889:data<=-16'd731;
      96890:data<=16'd1384;
      96891:data<=16'd2202;
      96892:data<=16'd1610;
      96893:data<=16'd1748;
      96894:data<=16'd2673;
      96895:data<=16'd2681;
      96896:data<=16'd2793;
      96897:data<=16'd3553;
      96898:data<=16'd2917;
      96899:data<=16'd2547;
      96900:data<=16'd2878;
      96901:data<=16'd1964;
      96902:data<=16'd2623;
      96903:data<=16'd2749;
      96904:data<=-16'd1239;
      96905:data<=-16'd3266;
      96906:data<=-16'd2645;
      96907:data<=-16'd3089;
      96908:data<=-16'd2184;
      96909:data<=-16'd1158;
      96910:data<=-16'd1303;
      96911:data<=-16'd925;
      96912:data<=-16'd1272;
      96913:data<=-16'd785;
      96914:data<=16'd247;
      96915:data<=-16'd414;
      96916:data<=16'd429;
      96917:data<=16'd1741;
      96918:data<=16'd1918;
      96919:data<=16'd2584;
      96920:data<=16'd1330;
      96921:data<=16'd3386;
      96922:data<=16'd12420;
      96923:data<=16'd16991;
      96924:data<=16'd15424;
      96925:data<=16'd15200;
      96926:data<=16'd15045;
      96927:data<=16'd14380;
      96928:data<=16'd13814;
      96929:data<=16'd13098;
      96930:data<=16'd13885;
      96931:data<=16'd13938;
      96932:data<=16'd13144;
      96933:data<=16'd13776;
      96934:data<=16'd13238;
      96935:data<=16'd11905;
      96936:data<=16'd11568;
      96937:data<=16'd10778;
      96938:data<=16'd10237;
      96939:data<=16'd9962;
      96940:data<=16'd9135;
      96941:data<=16'd8581;
      96942:data<=16'd8830;
      96943:data<=16'd10654;
      96944:data<=16'd11894;
      96945:data<=16'd10657;
      96946:data<=16'd9761;
      96947:data<=16'd9270;
      96948:data<=16'd8655;
      96949:data<=16'd9294;
      96950:data<=16'd9365;
      96951:data<=16'd8648;
      96952:data<=16'd8146;
      96953:data<=16'd7360;
      96954:data<=16'd7053;
      96955:data<=16'd7235;
      96956:data<=16'd9700;
      96957:data<=16'd14084;
      96958:data<=16'd14912;
      96959:data<=16'd14048;
      96960:data<=16'd13957;
      96961:data<=16'd12513;
      96962:data<=16'd12739;
      96963:data<=16'd12637;
      96964:data<=16'd10534;
      96965:data<=16'd11459;
      96966:data<=16'd7620;
      96967:data<=-16'd2766;
      96968:data<=-16'd5096;
      96969:data<=-16'd1982;
      96970:data<=-16'd2064;
      96971:data<=-16'd1398;
      96972:data<=-16'd769;
      96973:data<=-16'd1720;
      96974:data<=-16'd1623;
      96975:data<=-16'd1325;
      96976:data<=-16'd1286;
      96977:data<=-16'd1874;
      96978:data<=-16'd2599;
      96979:data<=-16'd2023;
      96980:data<=-16'd2153;
      96981:data<=-16'd2340;
      96982:data<=-16'd896;
      96983:data<=16'd230;
      96984:data<=16'd863;
      96985:data<=16'd757;
      96986:data<=16'd64;
      96987:data<=16'd438;
      96988:data<=16'd217;
      96989:data<=-16'd664;
      96990:data<=-16'd397;
      96991:data<=-16'd14;
      96992:data<=16'd56;
      96993:data<=-16'd514;
      96994:data<=-16'd1348;
      96995:data<=-16'd907;
      96996:data<=-16'd196;
      96997:data<=16'd176;
      96998:data<=16'd203;
      96999:data<=-16'd124;
      97000:data<=16'd288;
      97001:data<=16'd130;
      97002:data<=-16'd299;
      97003:data<=16'd311;
      97004:data<=-16'd49;
      97005:data<=-16'd32;
      97006:data<=16'd209;
      97007:data<=-16'd1380;
      97008:data<=-16'd999;
      97009:data<=-16'd619;
      97010:data<=-16'd1803;
      97011:data<=16'd2534;
      97012:data<=16'd7755;
      97013:data<=16'd7078;
      97014:data<=16'd6363;
      97015:data<=16'd6608;
      97016:data<=16'd5662;
      97017:data<=16'd5103;
      97018:data<=16'd4523;
      97019:data<=16'd4435;
      97020:data<=16'd4053;
      97021:data<=16'd2977;
      97022:data<=16'd4235;
      97023:data<=16'd5771;
      97024:data<=16'd5413;
      97025:data<=16'd4861;
      97026:data<=16'd3808;
      97027:data<=16'd3290;
      97028:data<=16'd3375;
      97029:data<=16'd2546;
      97030:data<=16'd2396;
      97031:data<=16'd2275;
      97032:data<=16'd1572;
      97033:data<=16'd1773;
      97034:data<=16'd1474;
      97035:data<=16'd1333;
      97036:data<=16'd2255;
      97037:data<=16'd2353;
      97038:data<=16'd2693;
      97039:data<=16'd3175;
      97040:data<=16'd2281;
      97041:data<=16'd1653;
      97042:data<=16'd1580;
      97043:data<=16'd1196;
      97044:data<=16'd670;
      97045:data<=16'd466;
      97046:data<=16'd828;
      97047:data<=16'd604;
      97048:data<=16'd641;
      97049:data<=16'd1580;
      97050:data<=16'd1545;
      97051:data<=16'd1654;
      97052:data<=16'd1418;
      97053:data<=16'd365;
      97054:data<=16'd1072;
      97055:data<=-16'd2520;
      97056:data<=-16'd11649;
      97057:data<=-16'd14486;
      97058:data<=-16'd12336;
      97059:data<=-16'd12807;
      97060:data<=-16'd12571;
      97061:data<=-16'd11423;
      97062:data<=-16'd10351;
      97063:data<=-16'd6514;
      97064:data<=-16'd2799;
      97065:data<=-16'd2079;
      97066:data<=-16'd2502;
      97067:data<=-16'd2601;
      97068:data<=-16'd2466;
      97069:data<=-16'd3037;
      97070:data<=-16'd3372;
      97071:data<=-16'd2795;
      97072:data<=-16'd2799;
      97073:data<=-16'd3078;
      97074:data<=-16'd3510;
      97075:data<=-16'd3748;
      97076:data<=-16'd2537;
      97077:data<=-16'd2319;
      97078:data<=-16'd3491;
      97079:data<=-16'd3251;
      97080:data<=-16'd2854;
      97081:data<=-16'd3224;
      97082:data<=-16'd3501;
      97083:data<=-16'd4061;
      97084:data<=-16'd4238;
      97085:data<=-16'd4214;
      97086:data<=-16'd4443;
      97087:data<=-16'd4229;
      97088:data<=-16'd4748;
      97089:data<=-16'd6002;
      97090:data<=-16'd6484;
      97091:data<=-16'd6690;
      97092:data<=-16'd6837;
      97093:data<=-16'd6733;
      97094:data<=-16'd6419;
      97095:data<=-16'd5940;
      97096:data<=-16'd5768;
      97097:data<=-16'd5259;
      97098:data<=-16'd5277;
      97099:data<=-16'd5389;
      97100:data<=-16'd109;
      97101:data<=16'd7136;
      97102:data<=16'd6981;
      97103:data<=16'd3968;
      97104:data<=16'd4320;
      97105:data<=16'd4111;
      97106:data<=16'd3260;
      97107:data<=16'd3600;
      97108:data<=16'd2875;
      97109:data<=16'd2127;
      97110:data<=16'd2461;
      97111:data<=16'd2405;
      97112:data<=16'd2328;
      97113:data<=16'd1801;
      97114:data<=16'd1014;
      97115:data<=16'd866;
      97116:data<=-16'd2064;
      97117:data<=-16'd7233;
      97118:data<=-16'd8567;
      97119:data<=-16'd7313;
      97120:data<=-16'd7462;
      97121:data<=-16'd7771;
      97122:data<=-16'd7676;
      97123:data<=-16'd7347;
      97124:data<=-16'd6799;
      97125:data<=-16'd7181;
      97126:data<=-16'd6966;
      97127:data<=-16'd5830;
      97128:data<=-16'd6343;
      97129:data<=-16'd7392;
      97130:data<=-16'd7797;
      97131:data<=-16'd8270;
      97132:data<=-16'd7861;
      97133:data<=-16'd7301;
      97134:data<=-16'd7283;
      97135:data<=-16'd6819;
      97136:data<=-16'd6646;
      97137:data<=-16'd6420;
      97138:data<=-16'd6128;
      97139:data<=-16'd6536;
      97140:data<=-16'd6005;
      97141:data<=-16'd6531;
      97142:data<=-16'd8378;
      97143:data<=-16'd7077;
      97144:data<=-16'd8834;
      97145:data<=-16'd17482;
      97146:data<=-16'd21444;
      97147:data<=-16'd19429;
      97148:data<=-16'd19450;
      97149:data<=-16'd19209;
      97150:data<=-16'd17734;
      97151:data<=-16'd17785;
      97152:data<=-16'd16936;
      97153:data<=-16'd15300;
      97154:data<=-16'd15259;
      97155:data<=-16'd15737;
      97156:data<=-16'd16016;
      97157:data<=-16'd15781;
      97158:data<=-16'd14515;
      97159:data<=-16'd13828;
      97160:data<=-16'd14120;
      97161:data<=-16'd13400;
      97162:data<=-16'd12355;
      97163:data<=-16'd12422;
      97164:data<=-16'd11947;
      97165:data<=-16'd11060;
      97166:data<=-16'd10674;
      97167:data<=-16'd9805;
      97168:data<=-16'd10013;
      97169:data<=-16'd9549;
      97170:data<=-16'd5084;
      97171:data<=-16'd2649;
      97172:data<=-16'd3983;
      97173:data<=-16'd3209;
      97174:data<=-16'd2253;
      97175:data<=-16'd2466;
      97176:data<=-16'd1762;
      97177:data<=-16'd2056;
      97178:data<=-16'd2137;
      97179:data<=-16'd1582;
      97180:data<=-16'd2358;
      97181:data<=-16'd2590;
      97182:data<=-16'd3331;
      97183:data<=-16'd4162;
      97184:data<=-16'd2783;
      97185:data<=-16'd2990;
      97186:data<=-16'd3109;
      97187:data<=-16'd1754;
      97188:data<=-16'd3263;
      97189:data<=16'd103;
      97190:data<=16'd9835;
      97191:data<=16'd12236;
      97192:data<=16'd9855;
      97193:data<=16'd10874;
      97194:data<=16'd10147;
      97195:data<=16'd7511;
      97196:data<=16'd7145;
      97197:data<=16'd7174;
      97198:data<=16'd6461;
      97199:data<=16'd6184;
      97200:data<=16'd6617;
      97201:data<=16'd6948;
      97202:data<=16'd6766;
      97203:data<=16'd6602;
      97204:data<=16'd6256;
      97205:data<=16'd6114;
      97206:data<=16'd6479;
      97207:data<=16'd5950;
      97208:data<=16'd4501;
      97209:data<=16'd3638;
      97210:data<=16'd3838;
      97211:data<=16'd3829;
      97212:data<=16'd2936;
      97213:data<=16'd2787;
      97214:data<=16'd3198;
      97215:data<=16'd2986;
      97216:data<=16'd3031;
      97217:data<=16'd3219;
      97218:data<=16'd3359;
      97219:data<=16'd3381;
      97220:data<=16'd3039;
      97221:data<=16'd3081;
      97222:data<=16'd334;
      97223:data<=-16'd5021;
      97224:data<=-16'd6114;
      97225:data<=-16'd5228;
      97226:data<=-16'd5979;
      97227:data<=-16'd4928;
      97228:data<=-16'd4367;
      97229:data<=-16'd4736;
      97230:data<=-16'd3585;
      97231:data<=-16'd3906;
      97232:data<=-16'd3491;
      97233:data<=-16'd3991;
      97234:data<=-16'd11922;
      97235:data<=-16'd18102;
      97236:data<=-16'd17051;
      97237:data<=-16'd16836;
      97238:data<=-16'd16525;
      97239:data<=-16'd14248;
      97240:data<=-16'd13526;
      97241:data<=-16'd12845;
      97242:data<=-16'd11768;
      97243:data<=-16'd11356;
      97244:data<=-16'd10704;
      97245:data<=-16'd10202;
      97246:data<=-16'd9589;
      97247:data<=-16'd9498;
      97248:data<=-16'd10583;
      97249:data<=-16'd10589;
      97250:data<=-16'd9655;
      97251:data<=-16'd9247;
      97252:data<=-16'd8880;
      97253:data<=-16'd8385;
      97254:data<=-16'd7589;
      97255:data<=-16'd6589;
      97256:data<=-16'd5829;
      97257:data<=-16'd5644;
      97258:data<=-16'd5888;
      97259:data<=-16'd5143;
      97260:data<=-16'd4378;
      97261:data<=-16'd5046;
      97262:data<=-16'd5532;
      97263:data<=-16'd5492;
      97264:data<=-16'd4751;
      97265:data<=-16'd3592;
      97266:data<=-16'd3764;
      97267:data<=-16'd3325;
      97268:data<=-16'd2246;
      97269:data<=-16'd2517;
      97270:data<=-16'd2391;
      97271:data<=-16'd2379;
      97272:data<=-16'd1304;
      97273:data<=16'd849;
      97274:data<=-16'd1633;
      97275:data<=-16'd2353;
      97276:data<=16'd2834;
      97277:data<=16'd4131;
      97278:data<=16'd7517;
      97279:data<=16'd17129;
      97280:data<=16'd18973;
      97281:data<=16'd16537;
      97282:data<=16'd18116;
      97283:data<=16'd17243;
      97284:data<=16'd15640;
      97285:data<=16'd16075;
      97286:data<=16'd14945;
      97287:data<=16'd14566;
      97288:data<=16'd15062;
      97289:data<=16'd14152;
      97290:data<=16'd13421;
      97291:data<=16'd13170;
      97292:data<=16'd13176;
      97293:data<=16'd13198;
      97294:data<=16'd13151;
      97295:data<=16'd13435;
      97296:data<=16'd12888;
      97297:data<=16'd12377;
      97298:data<=16'd12181;
      97299:data<=16'd11110;
      97300:data<=16'd11532;
      97301:data<=16'd12743;
      97302:data<=16'd12581;
      97303:data<=16'd12783;
      97304:data<=16'd12258;
      97305:data<=16'd11072;
      97306:data<=16'd11441;
      97307:data<=16'd11492;
      97308:data<=16'd11013;
      97309:data<=16'd10499;
      97310:data<=16'd9589;
      97311:data<=16'd10151;
      97312:data<=16'd10163;
      97313:data<=16'd8575;
      97314:data<=16'd9197;
      97315:data<=16'd10584;
      97316:data<=16'd10257;
      97317:data<=16'd10017;
      97318:data<=16'd10184;
      97319:data<=16'd9549;
      97320:data<=16'd8445;
      97321:data<=16'd9207;
      97322:data<=16'd8942;
      97323:data<=16'd1918;
      97324:data<=-16'd5100;
      97325:data<=-16'd5583;
      97326:data<=-16'd5257;
      97327:data<=-16'd4487;
      97328:data<=-16'd2534;
      97329:data<=-16'd4949;
      97330:data<=-16'd8284;
      97331:data<=-16'd7642;
      97332:data<=-16'd6819;
      97333:data<=-16'd6734;
      97334:data<=-16'd6037;
      97335:data<=-16'd5897;
      97336:data<=-16'd5870;
      97337:data<=-16'd5204;
      97338:data<=-16'd4899;
      97339:data<=-16'd5224;
      97340:data<=-16'd4523;
      97341:data<=-16'd2590;
      97342:data<=-16'd1867;
      97343:data<=-16'd2099;
      97344:data<=-16'd1340;
      97345:data<=-16'd943;
      97346:data<=-16'd1585;
      97347:data<=-16'd1445;
      97348:data<=-16'd990;
      97349:data<=-16'd1333;
      97350:data<=-16'd954;
      97351:data<=-16'd199;
      97352:data<=-16'd901;
      97353:data<=-16'd652;
      97354:data<=16'd1539;
      97355:data<=16'd2594;
      97356:data<=16'd2717;
      97357:data<=16'd2622;
      97358:data<=16'd2064;
      97359:data<=16'd2588;
      97360:data<=16'd2931;
      97361:data<=16'd2772;
      97362:data<=16'd3237;
      97363:data<=16'd2256;
      97364:data<=16'd2312;
      97365:data<=16'd3428;
      97366:data<=16'd1277;
      97367:data<=16'd4661;
      97368:data<=16'd15477;
      97369:data<=16'd18657;
      97370:data<=16'd15964;
      97371:data<=16'd16700;
      97372:data<=16'd16222;
      97373:data<=16'd14756;
      97374:data<=16'd15217;
      97375:data<=16'd13981;
      97376:data<=16'd12759;
      97377:data<=16'd13265;
      97378:data<=16'd12639;
      97379:data<=16'd12073;
      97380:data<=16'd12337;
      97381:data<=16'd12148;
      97382:data<=16'd14070;
      97383:data<=16'd18174;
      97384:data<=16'd19161;
      97385:data<=16'd17018;
      97386:data<=16'd16407;
      97387:data<=16'd16698;
      97388:data<=16'd15970;
      97389:data<=16'd15406;
      97390:data<=16'd14885;
      97391:data<=16'd14324;
      97392:data<=16'd13872;
      97393:data<=16'd13173;
      97394:data<=16'd13847;
      97395:data<=16'd14892;
      97396:data<=16'd14061;
      97397:data<=16'd13118;
      97398:data<=16'd12213;
      97399:data<=16'd11077;
      97400:data<=16'd11100;
      97401:data<=16'd10543;
      97402:data<=16'd9597;
      97403:data<=16'd10035;
      97404:data<=16'd9905;
      97405:data<=16'd8950;
      97406:data<=16'd8396;
      97407:data<=16'd8740;
      97408:data<=16'd9984;
      97409:data<=16'd9247;
      97410:data<=16'd8103;
      97411:data<=16'd8960;
      97412:data<=16'd4394;
      97413:data<=-16'd4692;
      97414:data<=-16'd6858;
      97415:data<=-16'd4913;
      97416:data<=-16'd5594;
      97417:data<=-16'd5316;
      97418:data<=-16'd4716;
      97419:data<=-16'd5827;
      97420:data<=-16'd4793;
      97421:data<=-16'd2667;
      97422:data<=-16'd2432;
      97423:data<=-16'd2605;
      97424:data<=-16'd3043;
      97425:data<=-16'd3738;
      97426:data<=-16'd3767;
      97427:data<=-16'd3692;
      97428:data<=-16'd3504;
      97429:data<=-16'd3795;
      97430:data<=-16'd4034;
      97431:data<=-16'd2898;
      97432:data<=-16'd3410;
      97433:data<=-16'd3993;
      97434:data<=-16'd1024;
      97435:data<=-16'd1918;
      97436:data<=-16'd7558;
      97437:data<=-16'd8572;
      97438:data<=-16'd7492;
      97439:data<=-16'd8422;
      97440:data<=-16'd7932;
      97441:data<=-16'd7356;
      97442:data<=-16'd7310;
      97443:data<=-16'd6683;
      97444:data<=-16'd7383;
      97445:data<=-16'd7417;
      97446:data<=-16'd5729;
      97447:data<=-16'd4528;
      97448:data<=-16'd3773;
      97449:data<=-16'd4311;
      97450:data<=-16'd4661;
      97451:data<=-16'd3529;
      97452:data<=-16'd4355;
      97453:data<=-16'd4695;
      97454:data<=-16'd3397;
      97455:data<=-16'd4957;
      97456:data<=-16'd3034;
      97457:data<=16'd5526;
      97458:data<=16'd9652;
      97459:data<=16'd8316;
      97460:data<=16'd8877;
      97461:data<=16'd9996;
      97462:data<=16'd9233;
      97463:data<=16'd8216;
      97464:data<=16'd7956;
      97465:data<=16'd7973;
      97466:data<=16'd7429;
      97467:data<=16'd6334;
      97468:data<=16'd5197;
      97469:data<=16'd5086;
      97470:data<=16'd5944;
      97471:data<=16'd5413;
      97472:data<=16'd4235;
      97473:data<=16'd5339;
      97474:data<=16'd7664;
      97475:data<=16'd8666;
      97476:data<=16'd7976;
      97477:data<=16'd7083;
      97478:data<=16'd6880;
      97479:data<=16'd6458;
      97480:data<=16'd5814;
      97481:data<=16'd4831;
      97482:data<=16'd3533;
      97483:data<=16'd3647;
      97484:data<=16'd3935;
      97485:data<=16'd3271;
      97486:data<=16'd3145;
      97487:data<=16'd2772;
      97488:data<=16'd4131;
      97489:data<=16'd7730;
      97490:data<=16'd7460;
      97491:data<=16'd5445;
      97492:data<=16'd6143;
      97493:data<=16'd5706;
      97494:data<=16'd5078;
      97495:data<=16'd5348;
      97496:data<=16'd4049;
      97497:data<=16'd4034;
      97498:data<=16'd3753;
      97499:data<=16'd2196;
      97500:data<=16'd3579;
      97501:data<=16'd784;
      97502:data<=-16'd7935;
      97503:data<=-16'd10713;
      97504:data<=-16'd9417;
      97505:data<=-16'd10207;
      97506:data<=-16'd9749;
      97507:data<=-16'd9163;
      97508:data<=-16'd9338;
      97509:data<=-16'd8542;
      97510:data<=-16'd8943;
      97511:data<=-16'd9260;
      97512:data<=-16'd8211;
      97513:data<=-16'd8830;
      97514:data<=-16'd10381;
      97515:data<=-16'd10658;
      97516:data<=-16'd10342;
      97517:data<=-16'd10401;
      97518:data<=-16'd10510;
      97519:data<=-16'd9902;
      97520:data<=-16'd9735;
      97521:data<=-16'd10017;
      97522:data<=-16'd9122;
      97523:data<=-16'd8731;
      97524:data<=-16'd9185;
      97525:data<=-16'd8801;
      97526:data<=-16'd9468;
      97527:data<=-16'd10860;
      97528:data<=-16'd10301;
      97529:data<=-16'd9658;
      97530:data<=-16'd9999;
      97531:data<=-16'd9280;
      97532:data<=-16'd8548;
      97533:data<=-16'd9259;
      97534:data<=-16'd9524;
      97535:data<=-16'd9085;
      97536:data<=-16'd8977;
      97537:data<=-16'd8055;
      97538:data<=-16'd7506;
      97539:data<=-16'd8719;
      97540:data<=-16'd9256;
      97541:data<=-16'd10175;
      97542:data<=-16'd12722;
      97543:data<=-16'd13573;
      97544:data<=-16'd13473;
      97545:data<=-16'd12170;
      97546:data<=-16'd6264;
      97547:data<=-16'd957;
      97548:data<=-16'd725;
      97549:data<=-16'd1465;
      97550:data<=-16'd1571;
      97551:data<=-16'd1618;
      97552:data<=-16'd1615;
      97553:data<=-16'd2705;
      97554:data<=-16'd3956;
      97555:data<=-16'd4276;
      97556:data<=-16'd3971;
      97557:data<=-16'd3359;
      97558:data<=-16'd3509;
      97559:data<=-16'd3946;
      97560:data<=-16'd3883;
      97561:data<=-16'd3932;
      97562:data<=-16'd3603;
      97563:data<=-16'd3330;
      97564:data<=-16'd3510;
      97565:data<=-16'd3156;
      97566:data<=-16'd3733;
      97567:data<=-16'd5447;
      97568:data<=-16'd5861;
      97569:data<=-16'd5539;
      97570:data<=-16'd5483;
      97571:data<=-16'd5098;
      97572:data<=-16'd5078;
      97573:data<=-16'd5524;
      97574:data<=-16'd5147;
      97575:data<=-16'd4769;
      97576:data<=-16'd5782;
      97577:data<=-16'd5994;
      97578:data<=-16'd4770;
      97579:data<=-16'd5386;
      97580:data<=-16'd6699;
      97581:data<=-16'd6479;
      97582:data<=-16'd6575;
      97583:data<=-16'd6273;
      97584:data<=-16'd5389;
      97585:data<=-16'd5541;
      97586:data<=-16'd5335;
      97587:data<=-16'd5833;
      97588:data<=-16'd6172;
      97589:data<=-16'd3950;
      97590:data<=-16'd6326;
      97591:data<=-16'd13582;
      97592:data<=-16'd16102;
      97593:data<=-16'd16119;
      97594:data<=-16'd16230;
      97595:data<=-16'd12847;
      97596:data<=-16'd10561;
      97597:data<=-16'd10924;
      97598:data<=-16'd9674;
      97599:data<=-16'd8933;
      97600:data<=-16'd9368;
      97601:data<=-16'd8727;
      97602:data<=-16'd8116;
      97603:data<=-16'd7755;
      97604:data<=-16'd7245;
      97605:data<=-16'd7318;
      97606:data<=-16'd8316;
      97607:data<=-16'd9906;
      97608:data<=-16'd10079;
      97609:data<=-16'd8595;
      97610:data<=-16'd7908;
      97611:data<=-16'd7947;
      97612:data<=-16'd7603;
      97613:data<=-16'd7442;
      97614:data<=-16'd7160;
      97615:data<=-16'd5943;
      97616:data<=-16'd5012;
      97617:data<=-16'd5068;
      97618:data<=-16'd4410;
      97619:data<=-16'd4303;
      97620:data<=-16'd6402;
      97621:data<=-16'd6689;
      97622:data<=-16'd4940;
      97623:data<=-16'd5016;
      97624:data<=-16'd4993;
      97625:data<=-16'd4434;
      97626:data<=-16'd5074;
      97627:data<=-16'd4610;
      97628:data<=-16'd3783;
      97629:data<=-16'd3953;
      97630:data<=-16'd3606;
      97631:data<=-16'd3509;
      97632:data<=-16'd3200;
      97633:data<=-16'd3556;
      97634:data<=-16'd5336;
      97635:data<=-16'd1506;
      97636:data<=16'd6285;
      97637:data<=16'd7865;
      97638:data<=16'd6493;
      97639:data<=16'd6909;
      97640:data<=16'd6158;
      97641:data<=16'd5877;
      97642:data<=16'd6416;
      97643:data<=16'd5814;
      97644:data<=16'd5993;
      97645:data<=16'd5861;
      97646:data<=16'd4499;
      97647:data<=16'd3529;
      97648:data<=16'd1202;
      97649:data<=-16'd1078;
      97650:data<=-16'd462;
      97651:data<=16'd35;
      97652:data<=-16'd320;
      97653:data<=-16'd44;
      97654:data<=-16'd611;
      97655:data<=-16'd1077;
      97656:data<=-16'd146;
      97657:data<=16'd557;
      97658:data<=16'd576;
      97659:data<=-16'd209;
      97660:data<=-16'd1626;
      97661:data<=-16'd2071;
      97662:data<=-16'd1415;
      97663:data<=-16'd675;
      97664:data<=-16'd907;
      97665:data<=-16'd1724;
      97666:data<=-16'd905;
      97667:data<=16'd187;
      97668:data<=-16'd456;
      97669:data<=-16'd481;
      97670:data<=16'd159;
      97671:data<=16'd138;
      97672:data<=16'd279;
      97673:data<=-16'd1004;
      97674:data<=-16'd2708;
      97675:data<=-16'd1574;
      97676:data<=-16'd887;
      97677:data<=-16'd1612;
      97678:data<=-16'd675;
      97679:data<=-16'd2690;
      97680:data<=-16'd9415;
      97681:data<=-16'd12815;
      97682:data<=-16'd11388;
      97683:data<=-16'd10290;
      97684:data<=-16'd10058;
      97685:data<=-16'd10103;
      97686:data<=-16'd10763;
      97687:data<=-16'd10766;
      97688:data<=-16'd10207;
      97689:data<=-16'd9881;
      97690:data<=-16'd9085;
      97691:data<=-16'd7873;
      97692:data<=-16'd6922;
      97693:data<=-16'd6570;
      97694:data<=-16'd6775;
      97695:data<=-16'd6476;
      97696:data<=-16'd5745;
      97697:data<=-16'd5474;
      97698:data<=-16'd4993;
      97699:data<=-16'd4942;
      97700:data<=-16'd6034;
      97701:data<=-16'd5098;
      97702:data<=-16'd1539;
      97703:data<=16'd232;
      97704:data<=-16'd74;
      97705:data<=16'd657;
      97706:data<=16'd1676;
      97707:data<=16'd1829;
      97708:data<=16'd1924;
      97709:data<=16'd1856;
      97710:data<=16'd2056;
      97711:data<=16'd2353;
      97712:data<=16'd1762;
      97713:data<=16'd1841;
      97714:data<=16'd2578;
      97715:data<=16'd2461;
      97716:data<=16'd2246;
      97717:data<=16'd1729;
      97718:data<=16'd2385;
      97719:data<=16'd4728;
      97720:data<=16'd4269;
      97721:data<=16'd3256;
      97722:data<=16'd4225;
      97723:data<=16'd3162;
      97724:data<=16'd5899;
      97725:data<=16'd14546;
      97726:data<=16'd17482;
      97727:data<=16'd15758;
      97728:data<=16'd16422;
      97729:data<=16'd16374;
      97730:data<=16'd15344;
      97731:data<=16'd15111;
      97732:data<=16'd15215;
      97733:data<=16'd15618;
      97734:data<=16'd14645;
      97735:data<=16'd13596;
      97736:data<=16'd13203;
      97737:data<=16'd11635;
      97738:data<=16'd12281;
      97739:data<=16'd14706;
      97740:data<=16'd14584;
      97741:data<=16'd14352;
      97742:data<=16'd14402;
      97743:data<=16'd13000;
      97744:data<=16'd12378;
      97745:data<=16'd12205;
      97746:data<=16'd12058;
      97747:data<=16'd12800;
      97748:data<=16'd12339;
      97749:data<=16'd10995;
      97750:data<=16'd10546;
      97751:data<=16'd10270;
      97752:data<=16'd11488;
      97753:data<=16'd13729;
      97754:data<=16'd11794;
      97755:data<=16'd7427;
      97756:data<=16'd7104;
      97757:data<=16'd8094;
      97758:data<=16'd6805;
      97759:data<=16'd6206;
      97760:data<=16'd6097;
      97761:data<=16'd5780;
      97762:data<=16'd6408;
      97763:data<=16'd6078;
      97764:data<=16'd5380;
      97765:data<=16'd5510;
      97766:data<=16'd5832;
      97767:data<=16'd7558;
      97768:data<=16'd6579;
      97769:data<=16'd126;
      97770:data<=-16'd4397;
      97771:data<=-16'd4264;
      97772:data<=-16'd3356;
      97773:data<=-16'd3174;
      97774:data<=-16'd3674;
      97775:data<=-16'd3665;
      97776:data<=-16'd3805;
      97777:data<=-16'd4300;
      97778:data<=-16'd2511;
      97779:data<=16'd20;
      97780:data<=16'd998;
      97781:data<=16'd710;
      97782:data<=-16'd167;
      97783:data<=16'd651;
      97784:data<=16'd1280;
      97785:data<=-16'd522;
      97786:data<=-16'd1127;
      97787:data<=-16'd244;
      97788:data<=16'd296;
      97789:data<=16'd138;
      97790:data<=-16'd699;
      97791:data<=16'd698;
      97792:data<=16'd2517;
      97793:data<=16'd1864;
      97794:data<=16'd2064;
      97795:data<=16'd2206;
      97796:data<=16'd1623;
      97797:data<=16'd2544;
      97798:data<=16'd2593;
      97799:data<=16'd2672;
      97800:data<=16'd3298;
      97801:data<=16'd2264;
      97802:data<=16'd2381;
      97803:data<=16'd2672;
      97804:data<=16'd2381;
      97805:data<=16'd3985;
      97806:data<=16'd4161;
      97807:data<=16'd5257;
      97808:data<=16'd8822;
      97809:data<=16'd8352;
      97810:data<=16'd8025;
      97811:data<=16'd9065;
      97812:data<=16'd6264;
      97813:data<=16'd8539;
      97814:data<=16'd16597;
      97815:data<=16'd18892;
      97816:data<=16'd17232;
      97817:data<=16'd16126;
      97818:data<=16'd15770;
      97819:data<=16'd17215;
      97820:data<=16'd17202;
      97821:data<=16'd15383;
      97822:data<=16'd14806;
      97823:data<=16'd14415;
      97824:data<=16'd14204;
      97825:data<=16'd14266;
      97826:data<=16'd13555;
      97827:data<=16'd13160;
      97828:data<=16'd12525;
      97829:data<=16'd11406;
      97830:data<=16'd11418;
      97831:data<=16'd11345;
      97832:data<=16'd10531;
      97833:data<=16'd10495;
      97834:data<=16'd10969;
      97835:data<=16'd10965;
      97836:data<=16'd10111;
      97837:data<=16'd9144;
      97838:data<=16'd9103;
      97839:data<=16'd8866;
      97840:data<=16'd7837;
      97841:data<=16'd7009;
      97842:data<=16'd6234;
      97843:data<=16'd5753;
      97844:data<=16'd5849;
      97845:data<=16'd6018;
      97846:data<=16'd6586;
      97847:data<=16'd6393;
      97848:data<=16'd5147;
      97849:data<=16'd5718;
      97850:data<=16'd6869;
      97851:data<=16'd5538;
      97852:data<=16'd4026;
      97853:data<=16'd4197;
      97854:data<=16'd4050;
      97855:data<=16'd3039;
      97856:data<=16'd2980;
      97857:data<=16'd2350;
      97858:data<=-16'd2093;
      97859:data<=-16'd6384;
      97860:data<=-16'd7066;
      97861:data<=-16'd8440;
      97862:data<=-16'd10276;
      97863:data<=-16'd10144;
      97864:data<=-16'd10314;
      97865:data<=-16'd9932;
      97866:data<=-16'd9085;
      97867:data<=-16'd9773;
      97868:data<=-16'd9744;
      97869:data<=-16'd9433;
      97870:data<=-16'd9614;
      97871:data<=-16'd8129;
      97872:data<=-16'd6478;
      97873:data<=-16'd5550;
      97874:data<=-16'd5380;
      97875:data<=-16'd6575;
      97876:data<=-16'd6305;
      97877:data<=-16'd5372;
      97878:data<=-16'd6272;
      97879:data<=-16'd6485;
      97880:data<=-16'd6067;
      97881:data<=-16'd6464;
      97882:data<=-16'd6523;
      97883:data<=-16'd6417;
      97884:data<=-16'd6241;
      97885:data<=-16'd5244;
      97886:data<=-16'd3436;
      97887:data<=-16'd2414;
      97888:data<=-16'd3092;
      97889:data<=-16'd3046;
      97890:data<=-16'd2346;
      97891:data<=-16'd2604;
      97892:data<=-16'd2773;
      97893:data<=-16'd3742;
      97894:data<=-16'd4793;
      97895:data<=-16'd4029;
      97896:data<=-16'd3145;
      97897:data<=-16'd1997;
      97898:data<=-16'd1219;
      97899:data<=-16'd1378;
      97900:data<=-16'd757;
      97901:data<=-16'd1642;
      97902:data<=-16'd144;
      97903:data<=16'd7319;
      97904:data<=16'd10364;
      97905:data<=16'd8499;
      97906:data<=16'd8561;
      97907:data<=16'd7106;
      97908:data<=16'd6234;
      97909:data<=16'd7233;
      97910:data<=16'd5661;
      97911:data<=16'd5844;
      97912:data<=16'd7712;
      97913:data<=16'd7383;
      97914:data<=16'd8426;
      97915:data<=16'd10084;
      97916:data<=16'd10137;
      97917:data<=16'd9646;
      97918:data<=16'd8592;
      97919:data<=16'd8225;
      97920:data<=16'd7497;
      97921:data<=16'd6451;
      97922:data<=16'd6893;
      97923:data<=16'd5977;
      97924:data<=16'd5413;
      97925:data<=16'd6757;
      97926:data<=16'd5638;
      97927:data<=16'd4494;
      97928:data<=16'd4634;
      97929:data<=16'd3243;
      97930:data<=16'd2963;
      97931:data<=16'd3019;
      97932:data<=16'd1851;
      97933:data<=16'd1786;
      97934:data<=16'd1530;
      97935:data<=16'd1128;
      97936:data<=16'd1192;
      97937:data<=-16'd39;
      97938:data<=-16'd1342;
      97939:data<=-16'd1935;
      97940:data<=-16'd1989;
      97941:data<=-16'd2226;
      97942:data<=-16'd3344;
      97943:data<=-16'd3002;
      97944:data<=-16'd3372;
      97945:data<=-16'd4637;
      97946:data<=-16'd2581;
      97947:data<=-16'd5330;
      97948:data<=-16'd14408;
      97949:data<=-16'd16589;
      97950:data<=-16'd14304;
      97951:data<=-16'd14871;
      97952:data<=-16'd14756;
      97953:data<=-16'd14465;
      97954:data<=-16'd14777;
      97955:data<=-16'd14648;
      97956:data<=-16'd15300;
      97957:data<=-16'd14857;
      97958:data<=-16'd13741;
      97959:data<=-16'd13295;
      97960:data<=-16'd12105;
      97961:data<=-16'd12340;
      97962:data<=-16'd13365;
      97963:data<=-16'd12451;
      97964:data<=-16'd12304;
      97965:data<=-16'd13109;
      97966:data<=-16'd13567;
      97967:data<=-16'd15314;
      97968:data<=-16'd16756;
      97969:data<=-16'd16272;
      97970:data<=-16'd16126;
      97971:data<=-16'd16832;
      97972:data<=-16'd16099;
      97973:data<=-16'd14216;
      97974:data<=-16'd13887;
      97975:data<=-16'd14211;
      97976:data<=-16'd13403;
      97977:data<=-16'd13179;
      97978:data<=-16'd13803;
      97979:data<=-16'd13646;
      97980:data<=-16'd12657;
      97981:data<=-16'd12067;
      97982:data<=-16'd12211;
      97983:data<=-16'd11251;
      97984:data<=-16'd9897;
      97985:data<=-16'd10100;
      97986:data<=-16'd10119;
      97987:data<=-16'd10060;
      97988:data<=-16'd10249;
      97989:data<=-16'd9385;
      97990:data<=-16'd9535;
      97991:data<=-16'd8147;
      97992:data<=-16'd2223;
      97993:data<=16'd1369;
      97994:data<=16'd843;
      97995:data<=16'd829;
      97996:data<=16'd693;
      97997:data<=16'd549;
      97998:data<=16'd1054;
      97999:data<=16'd1045;
      98000:data<=16'd1560;
      98001:data<=16'd1850;
      98002:data<=16'd1127;
      98003:data<=16'd943;
      98004:data<=16'd405;
      98005:data<=-16'd647;
      98006:data<=-16'd886;
      98007:data<=-16'd1224;
      98008:data<=-16'd1600;
      98009:data<=-16'd1160;
      98010:data<=-16'd1002;
      98011:data<=-16'd1271;
      98012:data<=-16'd805;
      98013:data<=-16'd258;
      98014:data<=-16'd443;
      98015:data<=-16'd578;
      98016:data<=-16'd611;
      98017:data<=-16'd867;
      98018:data<=-16'd1851;
      98019:data<=-16'd3180;
      98020:data<=-16'd1459;
      98021:data<=16'd1610;
      98022:data<=16'd1187;
      98023:data<=16'd886;
      98024:data<=16'd2073;
      98025:data<=16'd1163;
      98026:data<=16'd814;
      98027:data<=16'd1193;
      98028:data<=16'd870;
      98029:data<=16'd2144;
      98030:data<=16'd1324;
      98031:data<=-16'd1609;
      98032:data<=-16'd1300;
      98033:data<=-16'd1372;
      98034:data<=-16'd2344;
      98035:data<=-16'd1257;
      98036:data<=-16'd4220;
      98037:data<=-16'd10803;
      98038:data<=-16'd12836;
      98039:data<=-16'd11479;
      98040:data<=-16'd10919;
      98041:data<=-16'd10546;
      98042:data<=-16'd9755;
      98043:data<=-16'd9195;
      98044:data<=-16'd9909;
      98045:data<=-16'd11606;
      98046:data<=-16'd11306;
      98047:data<=-16'd9074;
      98048:data<=-16'd8853;
      98049:data<=-16'd9439;
      98050:data<=-16'd8360;
      98051:data<=-16'd8414;
      98052:data<=-16'd8607;
      98053:data<=-16'd7382;
      98054:data<=-16'd8296;
      98055:data<=-16'd8801;
      98056:data<=-16'd6510;
      98057:data<=-16'd6246;
      98058:data<=-16'd7413;
      98059:data<=-16'd7533;
      98060:data<=-16'd7806;
      98061:data<=-16'd7401;
      98062:data<=-16'd6654;
      98063:data<=-16'd5987;
      98064:data<=-16'd4620;
      98065:data<=-16'd4064;
      98066:data<=-16'd4038;
      98067:data<=-16'd4229;
      98068:data<=-16'd4764;
      98069:data<=-16'd3489;
      98070:data<=-16'd3099;
      98071:data<=-16'd5127;
      98072:data<=-16'd5063;
      98073:data<=-16'd5104;
      98074:data<=-16'd7620;
      98075:data<=-16'd8006;
      98076:data<=-16'd7119;
      98077:data<=-16'd7333;
      98078:data<=-16'd6951;
      98079:data<=-16'd7069;
      98080:data<=-16'd5624;
      98081:data<=16'd980;
      98082:data<=16'd6284;
      98083:data<=16'd5520;
      98084:data<=16'd3971;
      98085:data<=16'd3855;
      98086:data<=16'd3579;
      98087:data<=16'd3582;
      98088:data<=16'd3375;
      98089:data<=16'd3471;
      98090:data<=16'd4449;
      98091:data<=16'd4093;
      98092:data<=16'd3297;
      98093:data<=16'd3753;
      98094:data<=16'd3234;
      98095:data<=16'd2255;
      98096:data<=16'd3306;
      98097:data<=16'd4314;
      98098:data<=16'd2842;
      98099:data<=16'd1155;
      98100:data<=16'd1559;
      98101:data<=16'd2176;
      98102:data<=16'd2043;
      98103:data<=16'd2538;
      98104:data<=16'd2814;
      98105:data<=16'd2264;
      98106:data<=16'd1823;
      98107:data<=16'd1692;
      98108:data<=16'd2429;
      98109:data<=16'd3174;
      98110:data<=16'd2150;
      98111:data<=16'd450;
      98112:data<=16'd320;
      98113:data<=16'd1535;
      98114:data<=16'd1096;
      98115:data<=-16'd205;
      98116:data<=16'd1166;
      98117:data<=16'd1953;
      98118:data<=16'd617;
      98119:data<=16'd926;
      98120:data<=16'd1061;
      98121:data<=16'd628;
      98122:data<=16'd1630;
      98123:data<=16'd1930;
      98124:data<=16'd1572;
      98125:data<=-16'd2071;
      98126:data<=-16'd8937;
      98127:data<=-16'd8727;
      98128:data<=-16'd4199;
      98129:data<=-16'd4798;
      98130:data<=-16'd5357;
      98131:data<=-16'd4152;
      98132:data<=-16'd4285;
      98133:data<=-16'd3328;
      98134:data<=-16'd2719;
      98135:data<=-16'd2732;
      98136:data<=-16'd1351;
      98137:data<=-16'd1324;
      98138:data<=-16'd1847;
      98139:data<=-16'd1037;
      98140:data<=-16'd1057;
      98141:data<=-16'd1394;
      98142:data<=-16'd1162;
      98143:data<=-16'd1028;
      98144:data<=-16'd415;
      98145:data<=16'd130;
      98146:data<=-16'd244;
      98147:data<=-16'd626;
      98148:data<=-16'd514;
      98149:data<=16'd102;
      98150:data<=16'd2018;
      98151:data<=16'd3952;
      98152:data<=16'd3961;
      98153:data<=16'd4432;
      98154:data<=16'd5369;
      98155:data<=16'd4343;
      98156:data<=16'd4728;
      98157:data<=16'd6073;
      98158:data<=16'd4928;
      98159:data<=16'd4861;
      98160:data<=16'd5154;
      98161:data<=16'd3533;
      98162:data<=16'd3744;
      98163:data<=16'd4963;
      98164:data<=16'd6472;
      98165:data<=16'd8367;
      98166:data<=16'd7301;
      98167:data<=16'd6393;
      98168:data<=16'd6162;
      98169:data<=16'd4978;
      98170:data<=16'd10151;
      98171:data<=16'd17484;
      98172:data<=16'd17570;
      98173:data<=16'd16625;
      98174:data<=16'd16818;
      98175:data<=16'd15209;
      98176:data<=16'd15379;
      98177:data<=16'd16621;
      98178:data<=16'd16390;
      98179:data<=16'd14568;
      98180:data<=16'd11841;
      98181:data<=16'd10988;
      98182:data<=16'd10393;
      98183:data<=16'd9103;
      98184:data<=16'd9853;
      98185:data<=16'd10208;
      98186:data<=16'd9714;
      98187:data<=16'd9926;
      98188:data<=16'd8696;
      98189:data<=16'd8249;
      98190:data<=16'd9859;
      98191:data<=16'd10404;
      98192:data<=16'd10513;
      98193:data<=16'd10448;
      98194:data<=16'd9580;
      98195:data<=16'd9091;
      98196:data<=16'd8469;
      98197:data<=16'd7527;
      98198:data<=16'd6805;
      98199:data<=16'd6561;
      98200:data<=16'd6925;
      98201:data<=16'd6830;
      98202:data<=16'd6423;
      98203:data<=16'd6446;
      98204:data<=16'd7608;
      98205:data<=16'd9350;
      98206:data<=16'd8372;
      98207:data<=16'd7034;
      98208:data<=16'd7877;
      98209:data<=16'd6713;
      98210:data<=16'd5506;
      98211:data<=16'd5692;
      98212:data<=16'd4708;
      98213:data<=16'd6191;
      98214:data<=16'd4814;
      98215:data<=-16'd3694;
      98216:data<=-16'd6169;
      98217:data<=-16'd2406;
      98218:data<=-16'd2159;
      98219:data<=-16'd2058;
      98220:data<=-16'd1506;
      98221:data<=-16'd2422;
      98222:data<=-16'd1823;
      98223:data<=-16'd1463;
      98224:data<=-16'd2773;
      98225:data<=-16'd3287;
      98226:data<=-16'd2294;
      98227:data<=-16'd1742;
      98228:data<=-16'd2088;
      98229:data<=-16'd185;
      98230:data<=16'd1262;
      98231:data<=-16'd525;
      98232:data<=16'd1014;
      98233:data<=16'd5025;
      98234:data<=16'd5341;
      98235:data<=16'd3880;
      98236:data<=16'd3060;
      98237:data<=16'd3805;
      98238:data<=16'd4156;
      98239:data<=16'd2594;
      98240:data<=16'd3486;
      98241:data<=16'd4699;
      98242:data<=16'd3941;
      98243:data<=16'd5060;
      98244:data<=16'd5565;
      98245:data<=16'd5861;
      98246:data<=16'd7150;
      98247:data<=16'd5495;
      98248:data<=16'd5450;
      98249:data<=16'd6476;
      98250:data<=16'd3774;
      98251:data<=16'd3650;
      98252:data<=16'd4878;
      98253:data<=16'd4161;
      98254:data<=16'd4675;
      98255:data<=16'd3720;
      98256:data<=16'd4405;
      98257:data<=16'd6678;
      98258:data<=16'd4273;
      98259:data<=16'd7494;
      98260:data<=16'd16507;
      98261:data<=16'd17186;
      98262:data<=16'd14680;
      98263:data<=16'd14647;
      98264:data<=16'd13436;
      98265:data<=16'd12754;
      98266:data<=16'd12737;
      98267:data<=16'd12665;
      98268:data<=16'd11662;
      98269:data<=16'd10016;
      98270:data<=16'd11335;
      98271:data<=16'd12014;
      98272:data<=16'd11118;
      98273:data<=16'd11820;
      98274:data<=16'd10066;
      98275:data<=16'd8781;
      98276:data<=16'd9896;
      98277:data<=16'd7773;
      98278:data<=16'd7512;
      98279:data<=16'd9453;
      98280:data<=16'd7636;
      98281:data<=16'd6504;
      98282:data<=16'd6311;
      98283:data<=16'd6875;
      98284:data<=16'd12060;
      98285:data<=16'd15896;
      98286:data<=16'd12765;
      98287:data<=16'd5009;
      98288:data<=16'd714;
      98289:data<=16'd3250;
      98290:data<=16'd2781;
      98291:data<=16'd373;
      98292:data<=16'd1994;
      98293:data<=16'd2690;
      98294:data<=16'd6940;
      98295:data<=16'd10063;
      98296:data<=16'd4382;
      98297:data<=16'd10343;
      98298:data<=16'd22436;
      98299:data<=16'd12886;
      98300:data<=-16'd4502;
      98301:data<=-16'd11438;
      98302:data<=-16'd11532;
      98303:data<=-16'd8871;
      98304:data<=-16'd10684;
      98305:data<=-16'd15597;
      98306:data<=-16'd20039;
      98307:data<=-16'd23575;
      98308:data<=-16'd16474;
      98309:data<=-16'd9024;
      98310:data<=-16'd14936;
      98311:data<=-16'd18339;
      98312:data<=-16'd15740;
      98313:data<=-16'd14230;
      98314:data<=-16'd11163;
      98315:data<=-16'd13928;
      98316:data<=-16'd18360;
      98317:data<=-16'd12154;
      98318:data<=-16'd6472;
      98319:data<=-16'd11496;
      98320:data<=-16'd21737;
      98321:data<=-16'd26480;
      98322:data<=-16'd21023;
      98323:data<=-16'd15095;
      98324:data<=-16'd11814;
      98325:data<=-16'd10912;
      98326:data<=-16'd18603;
      98327:data<=-16'd21851;
      98328:data<=-16'd12146;
      98329:data<=-16'd9056;
      98330:data<=-16'd15596;
      98331:data<=-16'd15168;
      98332:data<=-16'd9518;
      98333:data<=-16'd8787;
      98334:data<=-16'd8889;
      98335:data<=-16'd7089;
      98336:data<=-16'd10596;
      98337:data<=-16'd12730;
      98338:data<=-16'd6300;
      98339:data<=-16'd7820;
      98340:data<=-16'd19408;
      98341:data<=-16'd21294;
      98342:data<=-16'd15690;
      98343:data<=-16'd15803;
      98344:data<=-16'd17044;
      98345:data<=-16'd14765;
      98346:data<=-16'd16069;
      98347:data<=-16'd18120;
      98348:data<=-16'd9915;
      98349:data<=16'd522;
      98350:data<=16'd3454;
      98351:data<=16'd5037;
      98352:data<=16'd3257;
      98353:data<=-16'd3859;
      98354:data<=-16'd7104;
      98355:data<=-16'd5694;
      98356:data<=-16'd2740;
      98357:data<=16'd966;
      98358:data<=16'd2890;
      98359:data<=-16'd361;
      98360:data<=-16'd8573;
      98361:data<=-16'd8472;
      98362:data<=-16'd713;
      98363:data<=-16'd2746;
      98364:data<=-16'd5157;
      98365:data<=-16'd1807;
      98366:data<=-16'd4047;
      98367:data<=-16'd183;
      98368:data<=16'd9109;
      98369:data<=16'd7544;
      98370:data<=16'd5413;
      98371:data<=16'd8005;
      98372:data<=16'd7071;
      98373:data<=16'd2857;
      98374:data<=16'd664;
      98375:data<=16'd5436;
      98376:data<=16'd6625;
      98377:data<=16'd2908;
      98378:data<=16'd7885;
      98379:data<=16'd5651;
      98380:data<=-16'd7239;
      98381:data<=-16'd7577;
      98382:data<=-16'd3435;
      98383:data<=-16'd1729;
      98384:data<=16'd3404;
      98385:data<=16'd305;
      98386:data<=-16'd8804;
      98387:data<=-16'd12965;
      98388:data<=-16'd12313;
      98389:data<=-16'd7595;
      98390:data<=-16'd3127;
      98391:data<=16'd1322;
      98392:data<=-16'd1380;
      98393:data<=-16'd15743;
      98394:data<=-16'd16577;
      98395:data<=-16'd7752;
      98396:data<=-16'd13141;
      98397:data<=-16'd12972;
      98398:data<=-16'd4444;
      98399:data<=-16'd7709;
      98400:data<=-16'd8698;
      98401:data<=-16'd4021;
      98402:data<=-16'd7216;
      98403:data<=-16'd8066;
      98404:data<=-16'd787;
      98405:data<=16'd1080;
      98406:data<=-16'd7767;
      98407:data<=-16'd14524;
      98408:data<=-16'd10454;
      98409:data<=-16'd4103;
      98410:data<=-16'd1124;
      98411:data<=-16'd1459;
      98412:data<=-16'd4391;
      98413:data<=-16'd3142;
      98414:data<=16'd1233;
      98415:data<=16'd2701;
      98416:data<=16'd1897;
      98417:data<=16'd1215;
      98418:data<=16'd5456;
      98419:data<=16'd7887;
      98420:data<=16'd514;
      98421:data<=-16'd1181;
      98422:data<=16'd3824;
      98423:data<=16'd341;
      98424:data<=-16'd1936;
      98425:data<=16'd1293;
      98426:data<=-16'd1407;
      98427:data<=-16'd3342;
      98428:data<=16'd1941;
      98429:data<=16'd6419;
      98430:data<=16'd6637;
      98431:data<=16'd5150;
      98432:data<=16'd5328;
      98433:data<=16'd6953;
      98434:data<=16'd4047;
      98435:data<=-16'd2382;
      98436:data<=-16'd1730;
      98437:data<=16'd6000;
      98438:data<=16'd9050;
      98439:data<=16'd7553;
      98440:data<=16'd9709;
      98441:data<=16'd13223;
      98442:data<=16'd13164;
      98443:data<=16'd11694;
      98444:data<=16'd12104;
      98445:data<=16'd10337;
      98446:data<=16'd4905;
      98447:data<=16'd7555;
      98448:data<=16'd15053;
      98449:data<=16'd11888;
      98450:data<=16'd8317;
      98451:data<=16'd12132;
      98452:data<=16'd12759;
      98453:data<=16'd13608;
      98454:data<=16'd15074;
      98455:data<=16'd11220;
      98456:data<=16'd9988;
      98457:data<=16'd11634;
      98458:data<=16'd11370;
      98459:data<=16'd11981;
      98460:data<=16'd11030;
      98461:data<=16'd6473;
      98462:data<=16'd1903;
      98463:data<=16'd3638;
      98464:data<=16'd8978;
      98465:data<=16'd6972;
      98466:data<=16'd7650;
      98467:data<=16'd13718;
      98468:data<=16'd8560;
      98469:data<=16'd7782;
      98470:data<=16'd15700;
      98471:data<=16'd7759;
      98472:data<=16'd735;
      98473:data<=16'd5271;
      98474:data<=16'd1554;
      98475:data<=16'd2247;
      98476:data<=16'd9489;
      98477:data<=16'd3243;
      98478:data<=-16'd632;
      98479:data<=16'd7944;
      98480:data<=16'd8675;
      98481:data<=16'd926;
      98482:data<=-16'd1278;
      98483:data<=-16'd970;
      98484:data<=-16'd2094;
      98485:data<=16'd855;
      98486:data<=-16'd235;
      98487:data<=-16'd7401;
      98488:data<=-16'd2963;
      98489:data<=16'd2726;
      98490:data<=-16'd3882;
      98491:data<=-16'd3653;
      98492:data<=16'd224;
      98493:data<=-16'd4892;
      98494:data<=-16'd4514;
      98495:data<=16'd2065;
      98496:data<=16'd2910;
      98497:data<=-16'd1677;
      98498:data<=-16'd3553;
      98499:data<=16'd1183;
      98500:data<=16'd402;
      98501:data<=-16'd1460;
      98502:data<=16'd10073;
      98503:data<=16'd13885;
      98504:data<=16'd2353;
      98505:data<=-16'd943;
      98506:data<=16'd3347;
      98507:data<=16'd4278;
      98508:data<=16'd2061;
      98509:data<=16'd819;
      98510:data<=16'd5395;
      98511:data<=16'd6836;
      98512:data<=-16'd65;
      98513:data<=-16'd4144;
      98514:data<=-16'd4564;
      98515:data<=-16'd7673;
      98516:data<=-16'd7555;
      98517:data<=16'd1448;
      98518:data<=16'd4438;
      98519:data<=-16'd5488;
      98520:data<=-16'd6754;
      98521:data<=-16'd1149;
      98522:data<=-16'd4975;
      98523:data<=-16'd7092;
      98524:data<=-16'd7285;
      98525:data<=-16'd7859;
      98526:data<=16'd208;
      98527:data<=16'd3516;
      98528:data<=16'd1977;
      98529:data<=16'd5611;
      98530:data<=16'd4050;
      98531:data<=16'd4049;
      98532:data<=16'd6673;
      98533:data<=16'd476;
      98534:data<=-16'd1616;
      98535:data<=-16'd338;
      98536:data<=-16'd2393;
      98537:data<=16'd1618;
      98538:data<=16'd3668;
      98539:data<=16'd854;
      98540:data<=16'd472;
      98541:data<=-16'd831;
      98542:data<=-16'd230;
      98543:data<=-16'd438;
      98544:data<=-16'd3782;
      98545:data<=-16'd1700;
      98546:data<=-16'd382;
      98547:data<=-16'd4202;
      98548:data<=-16'd5723;
      98549:data<=-16'd3547;
      98550:data<=-16'd2232;
      98551:data<=-16'd8158;
      98552:data<=-16'd12612;
      98553:data<=-16'd8387;
      98554:data<=-16'd6476;
      98555:data<=-16'd5040;
      98556:data<=-16'd3222;
      98557:data<=-16'd5557;
      98558:data<=-16'd5482;
      98559:data<=-16'd9310;
      98560:data<=-16'd12668;
      98561:data<=-16'd6862;
      98562:data<=-16'd9489;
      98563:data<=-16'd10890;
      98564:data<=-16'd2422;
      98565:data<=-16'd7591;
      98566:data<=-16'd13273;
      98567:data<=-16'd8232;
      98568:data<=-16'd10554;
      98569:data<=-16'd13687;
      98570:data<=-16'd17105;
      98571:data<=-16'd26835;
      98572:data<=-16'd28056;
      98573:data<=-16'd22474;
      98574:data<=-16'd22789;
      98575:data<=-16'd26567;
      98576:data<=-16'd25795;
      98577:data<=-16'd23623;
      98578:data<=-16'd26735;
      98579:data<=-16'd23760;
      98580:data<=-16'd19560;
      98581:data<=-16'd27200;
      98582:data<=-16'd24861;
      98583:data<=-16'd16556;
      98584:data<=-16'd22418;
      98585:data<=-16'd23325;
      98586:data<=-16'd21047;
      98587:data<=-16'd24683;
      98588:data<=-16'd20359;
      98589:data<=-16'd17766;
      98590:data<=-16'd18409;
      98591:data<=-16'd16001;
      98592:data<=-16'd22063;
      98593:data<=-16'd24002;
      98594:data<=-16'd18700;
      98595:data<=-16'd20959;
      98596:data<=-16'd17250;
      98597:data<=-16'd8728;
      98598:data<=-16'd9564;
      98599:data<=-16'd12375;
      98600:data<=-16'd15117;
      98601:data<=-16'd14533;
      98602:data<=-16'd7978;
      98603:data<=-16'd4855;
      98604:data<=-16'd3785;
      98605:data<=-16'd4529;
      98606:data<=-16'd8179;
      98607:data<=-16'd6529;
      98608:data<=-16'd4623;
      98609:data<=-16'd5937;
      98610:data<=-16'd2370;
      98611:data<=16'd284;
      98612:data<=-16'd5553;
      98613:data<=-16'd9163;
      98614:data<=-16'd1145;
      98615:data<=16'd6018;
      98616:data<=16'd5175;
      98617:data<=16'd8407;
      98618:data<=16'd10181;
      98619:data<=16'd6774;
      98620:data<=16'd13543;
      98621:data<=16'd17964;
      98622:data<=16'd9168;
      98623:data<=16'd4382;
      98624:data<=16'd3096;
      98625:data<=16'd3591;
      98626:data<=16'd8915;
      98627:data<=16'd8181;
      98628:data<=16'd9262;
      98629:data<=16'd15800;
      98630:data<=16'd12148;
      98631:data<=16'd9036;
      98632:data<=16'd13197;
      98633:data<=16'd11156;
      98634:data<=16'd13150;
      98635:data<=16'd25504;
      98636:data<=16'd28652;
      98637:data<=16'd20019;
      98638:data<=16'd16352;
      98639:data<=16'd19930;
      98640:data<=16'd22301;
      98641:data<=16'd24768;
      98642:data<=16'd26714;
      98643:data<=16'd20818;
      98644:data<=16'd13019;
      98645:data<=16'd12844;
      98646:data<=16'd19026;
      98647:data<=16'd25058;
      98648:data<=16'd22465;
      98649:data<=16'd16037;
      98650:data<=16'd16991;
      98651:data<=16'd19444;
      98652:data<=16'd19403;
      98653:data<=16'd21318;
      98654:data<=16'd19902;
      98655:data<=16'd13250;
      98656:data<=16'd10783;
      98657:data<=16'd16530;
      98658:data<=16'd21284;
      98659:data<=16'd16939;
      98660:data<=16'd9562;
      98661:data<=16'd4579;
      98662:data<=16'd2340;
      98663:data<=16'd3703;
      98664:data<=16'd1703;
      98665:data<=-16'd863;
      98666:data<=16'd7110;
      98667:data<=16'd14299;
      98668:data<=16'd12733;
      98669:data<=16'd11684;
      98670:data<=16'd8217;
      98671:data<=16'd3228;
      98672:data<=16'd6381;
      98673:data<=16'd8552;
      98674:data<=16'd4490;
      98675:data<=16'd6335;
      98676:data<=16'd8410;
      98677:data<=16'd1430;
      98678:data<=16'd1844;
      98679:data<=16'd8834;
      98680:data<=16'd5177;
      98681:data<=16'd7001;
      98682:data<=16'd15778;
      98683:data<=16'd7471;
      98684:data<=16'd1736;
      98685:data<=16'd10890;
      98686:data<=16'd9632;
      98687:data<=16'd6211;
      98688:data<=16'd10213;
      98689:data<=16'd6249;
      98690:data<=16'd3045;
      98691:data<=16'd7808;
      98692:data<=16'd9280;
      98693:data<=16'd6028;
      98694:data<=16'd3633;
      98695:data<=16'd8786;
      98696:data<=16'd14750;
      98697:data<=16'd10258;
      98698:data<=16'd5835;
      98699:data<=16'd8244;
      98700:data<=16'd10564;
      98701:data<=16'd7031;
      98702:data<=-16'd2496;
      98703:data<=-16'd3051;
      98704:data<=16'd5883;
      98705:data<=16'd8977;
      98706:data<=16'd12897;
      98707:data<=16'd16381;
      98708:data<=16'd10850;
      98709:data<=16'd9871;
      98710:data<=16'd10912;
      98711:data<=16'd3953;
      98712:data<=16'd1224;
      98713:data<=16'd7174;
      98714:data<=16'd12373;
      98715:data<=16'd9535;
      98716:data<=16'd4799;
      98717:data<=16'd7247;
      98718:data<=16'd7118;
      98719:data<=16'd4636;
      98720:data<=16'd6310;
      98721:data<=16'd1870;
      98722:data<=16'd1105;
      98723:data<=16'd8705;
      98724:data<=16'd4052;
      98725:data<=-16'd2828;
      98726:data<=-16'd1415;
      98727:data<=-16'd4585;
      98728:data<=-16'd5503;
      98729:data<=-16'd2309;
      98730:data<=-16'd3204;
      98731:data<=-16'd2372;
      98732:data<=-16'd2181;
      98733:data<=-16'd2714;
      98734:data<=16'd227;
      98735:data<=-16'd2649;
      98736:data<=-16'd6161;
      98737:data<=-16'd2408;
      98738:data<=-16'd5068;
      98739:data<=-16'd13499;
      98740:data<=-16'd13453;
      98741:data<=-16'd8231;
      98742:data<=-16'd4828;
      98743:data<=-16'd3080;
      98744:data<=-16'd5776;
      98745:data<=-16'd9824;
      98746:data<=-16'd8375;
      98747:data<=-16'd10292;
      98748:data<=-16'd19074;
      98749:data<=-16'd21191;
      98750:data<=-16'd17902;
      98751:data<=-16'd15629;
      98752:data<=-16'd14037;
      98753:data<=-16'd19465;
      98754:data<=-16'd23572;
      98755:data<=-16'd19274;
      98756:data<=-16'd19509;
      98757:data<=-16'd18331;
      98758:data<=-16'd14571;
      98759:data<=-16'd21268;
      98760:data<=-16'd21743;
      98761:data<=-16'd15544;
      98762:data<=-16'd20566;
      98763:data<=-16'd18128;
      98764:data<=-16'd8210;
      98765:data<=-16'd13684;
      98766:data<=-16'd20118;
      98767:data<=-16'd15987;
      98768:data<=-16'd9976;
      98769:data<=-16'd2823;
      98770:data<=-16'd2775;
      98771:data<=-16'd12049;
      98772:data<=-16'd14145;
      98773:data<=-16'd8129;
      98774:data<=-16'd6736;
      98775:data<=-16'd8943;
      98776:data<=-16'd7413;
      98777:data<=-16'd4493;
      98778:data<=-16'd5254;
      98779:data<=-16'd7415;
      98780:data<=-16'd6990;
      98781:data<=-16'd5513;
      98782:data<=-16'd5365;
      98783:data<=-16'd3921;
      98784:data<=-16'd2390;
      98785:data<=-16'd3968;
      98786:data<=-16'd2167;
      98787:data<=-16'd1466;
      98788:data<=-16'd8085;
      98789:data<=-16'd4799;
      98790:data<=16'd793;
      98791:data<=-16'd8828;
      98792:data<=-16'd7063;
      98793:data<=16'd7010;
      98794:data<=16'd6570;
      98795:data<=16'd4846;
      98796:data<=16'd7169;
      98797:data<=16'd4952;
      98798:data<=16'd4896;
      98799:data<=16'd2126;
      98800:data<=16'd3510;
      98801:data<=16'd11473;
      98802:data<=16'd4943;
      98803:data<=-16'd473;
      98804:data<=16'd5181;
      98805:data<=16'd206;
      98806:data<=-16'd3559;
      98807:data<=16'd652;
      98808:data<=16'd1400;
      98809:data<=16'd4943;
      98810:data<=16'd2823;
      98811:data<=-16'd4490;
      98812:data<=-16'd1152;
      98813:data<=16'd905;
      98814:data<=16'd229;
      98815:data<=16'd3112;
      98816:data<=-16'd1962;
      98817:data<=-16'd5315;
      98818:data<=16'd302;
      98819:data<=-16'd241;
      98820:data<=-16'd4058;
      98821:data<=-16'd1930;
      98822:data<=16'd1290;
      98823:data<=16'd569;
      98824:data<=-16'd817;
      98825:data<=16'd1068;
      98826:data<=16'd384;
      98827:data<=-16'd1337;
      98828:data<=16'd2231;
      98829:data<=16'd2924;
      98830:data<=16'd3058;
      98831:data<=16'd7988;
      98832:data<=16'd4775;
      98833:data<=-16'd340;
      98834:data<=16'd6153;
      98835:data<=16'd6337;
      98836:data<=-16'd7474;
      98837:data<=-16'd14352;
      98838:data<=-16'd10693;
      98839:data<=-16'd8836;
      98840:data<=-16'd7703;
      98841:data<=-16'd7391;
      98842:data<=-16'd12584;
      98843:data<=-16'd14287;
      98844:data<=-16'd8907;
      98845:data<=-16'd6566;
      98846:data<=-16'd8320;
      98847:data<=-16'd8660;
      98848:data<=-16'd6655;
      98849:data<=-16'd7103;
      98850:data<=-16'd10096;
      98851:data<=-16'd5253;
      98852:data<=16'd1830;
      98853:data<=-16'd940;
      98854:data<=-16'd3301;
      98855:data<=-16'd1051;
      98856:data<=-16'd2275;
      98857:data<=-16'd4687;
      98858:data<=-16'd3685;
      98859:data<=16'd696;
      98860:data<=16'd1618;
      98861:data<=-16'd1178;
      98862:data<=-16'd341;
      98863:data<=-16'd3189;
      98864:data<=-16'd4848;
      98865:data<=16'd3523;
      98866:data<=16'd3988;
      98867:data<=16'd2685;
      98868:data<=16'd10448;
      98869:data<=16'd8188;
      98870:data<=16'd4858;
      98871:data<=16'd6428;
      98872:data<=-16'd1090;
      98873:data<=16'd1233;
      98874:data<=16'd11497;
      98875:data<=16'd8408;
      98876:data<=16'd7051;
      98877:data<=16'd10319;
      98878:data<=16'd11036;
      98879:data<=16'd13458;
      98880:data<=16'd10545;
      98881:data<=16'd12202;
      98882:data<=16'd23461;
      98883:data<=16'd21687;
      98884:data<=16'd13609;
      98885:data<=16'd15377;
      98886:data<=16'd17837;
      98887:data<=16'd18824;
      98888:data<=16'd20735;
      98889:data<=16'd20236;
      98890:data<=16'd16997;
      98891:data<=16'd14095;
      98892:data<=16'd15778;
      98893:data<=16'd18057;
      98894:data<=16'd18257;
      98895:data<=16'd19459;
      98896:data<=16'd17264;
      98897:data<=16'd14683;
      98898:data<=16'd16986;
      98899:data<=16'd16651;
      98900:data<=16'd15308;
      98901:data<=16'd16713;
      98902:data<=16'd16600;
      98903:data<=16'd19358;
      98904:data<=16'd23770;
      98905:data<=16'd22557;
      98906:data<=16'd21484;
      98907:data<=16'd22896;
      98908:data<=16'd21989;
      98909:data<=16'd20192;
      98910:data<=16'd18143;
      98911:data<=16'd17843;
      98912:data<=16'd21805;
      98913:data<=16'd20409;
      98914:data<=16'd12962;
      98915:data<=16'd14415;
      98916:data<=16'd18086;
      98917:data<=16'd12974;
      98918:data<=16'd13443;
      98919:data<=16'd17003;
      98920:data<=16'd10754;
      98921:data<=16'd9066;
      98922:data<=16'd12828;
      98923:data<=16'd10520;
      98924:data<=16'd10419;
      98925:data<=16'd6805;
      98926:data<=-16'd5389;
      98927:data<=-16'd7636;
      98928:data<=-16'd2455;
      98929:data<=-16'd878;
      98930:data<=16'd667;
      98931:data<=-16'd2370;
      98932:data<=-16'd6848;
      98933:data<=-16'd5265;
      98934:data<=-16'd5604;
      98935:data<=-16'd5768;
      98936:data<=-16'd1914;
      98937:data<=-16'd3653;
      98938:data<=-16'd8822;
      98939:data<=-16'd8969;
      98940:data<=-16'd5638;
      98941:data<=-16'd5817;
      98942:data<=-16'd10680;
      98943:data<=-16'd8868;
      98944:data<=-16'd4276;
      98945:data<=-16'd11614;
      98946:data<=-16'd17438;
      98947:data<=-16'd13235;
      98948:data<=-16'd12850;
      98949:data<=-16'd13212;
      98950:data<=-16'd10351;
      98951:data<=-16'd10322;
      98952:data<=-16'd9050;
      98953:data<=-16'd7941;
      98954:data<=-16'd11506;
      98955:data<=-16'd15875;
      98956:data<=-16'd18674;
      98957:data<=-16'd15555;
      98958:data<=-16'd9887;
      98959:data<=-16'd11169;
      98960:data<=-16'd13846;
      98961:data<=-16'd13452;
      98962:data<=-16'd11960;
      98963:data<=-16'd8868;
      98964:data<=-16'd10601;
      98965:data<=-16'd16049;
      98966:data<=-16'd16093;
      98967:data<=-16'd12825;
      98968:data<=-16'd10313;
      98969:data<=-16'd11361;
      98970:data<=-16'd13267;
      98971:data<=-16'd8472;
      98972:data<=-16'd5201;
      98973:data<=-16'd9397;
      98974:data<=-16'd13476;
      98975:data<=-16'd16829;
      98976:data<=-16'd16307;
      98977:data<=-16'd10290;
      98978:data<=-16'd8481;
      98979:data<=-16'd10637;
      98980:data<=-16'd11435;
      98981:data<=-16'd11655;
      98982:data<=-16'd11056;
      98983:data<=-16'd9059;
      98984:data<=-16'd6434;
      98985:data<=-16'd8067;
      98986:data<=-16'd10836;
      98987:data<=-16'd6191;
      98988:data<=-16'd6155;
      98989:data<=-16'd14011;
      98990:data<=-16'd14839;
      98991:data<=-16'd14680;
      98992:data<=-16'd13626;
      98993:data<=-16'd5359;
      98994:data<=-16'd9304;
      98995:data<=-16'd18766;
      98996:data<=-16'd10116;
      98997:data<=-16'd3375;
      98998:data<=-16'd11118;
      98999:data<=-16'd13671;
      99000:data<=-16'd9688;
      99001:data<=-16'd7351;
      99002:data<=-16'd5466;
      99003:data<=-16'd6393;
      99004:data<=-16'd9647;
      99005:data<=-16'd10534;
      99006:data<=-16'd10056;
      99007:data<=-16'd9418;
      99008:data<=-16'd8163;
      99009:data<=-16'd8766;
      99010:data<=-16'd12242;
      99011:data<=-16'd14634;
      99012:data<=-16'd12120;
      99013:data<=-16'd9809;
      99014:data<=-16'd15330;
      99015:data<=-16'd21456;
      99016:data<=-16'd20269;
      99017:data<=-16'd19564;
      99018:data<=-16'd20900;
      99019:data<=-16'd17666;
      99020:data<=-16'd14434;
      99021:data<=-16'd17452;
      99022:data<=-16'd20425;
      99023:data<=-16'd13944;
      99024:data<=-16'd8598;
      99025:data<=-16'd16695;
      99026:data<=-16'd19097;
      99027:data<=-16'd11065;
      99028:data<=-16'd13188;
      99029:data<=-16'd14684;
      99030:data<=-16'd8014;
      99031:data<=-16'd10088;
      99032:data<=-16'd13776;
      99033:data<=-16'd10310;
      99034:data<=-16'd6587;
      99035:data<=-16'd5683;
      99036:data<=-16'd7976;
      99037:data<=-16'd2522;
      99038:data<=16'd8040;
      99039:data<=16'd6761;
      99040:data<=16'd3171;
      99041:data<=16'd1627;
      99042:data<=-16'd1806;
      99043:data<=16'd2576;
      99044:data<=16'd6005;
      99045:data<=16'd6199;
      99046:data<=16'd11179;
      99047:data<=16'd9549;
      99048:data<=16'd8381;
      99049:data<=16'd11866;
      99050:data<=16'd7767;
      99051:data<=16'd9169;
      99052:data<=16'd13362;
      99053:data<=16'd9721;
      99054:data<=16'd11486;
      99055:data<=16'd10301;
      99056:data<=16'd6479;
      99057:data<=16'd13831;
      99058:data<=16'd14289;
      99059:data<=16'd10040;
      99060:data<=16'd16234;
      99061:data<=16'd19024;
      99062:data<=16'd18007;
      99063:data<=16'd19535;
      99064:data<=16'd20409;
      99065:data<=16'd23813;
      99066:data<=16'd23390;
      99067:data<=16'd15898;
      99068:data<=16'd11580;
      99069:data<=16'd12487;
      99070:data<=16'd16901;
      99071:data<=16'd22515;
      99072:data<=16'd24331;
      99073:data<=16'd21796;
      99074:data<=16'd18415;
      99075:data<=16'd16710;
      99076:data<=16'd15644;
      99077:data<=16'd18377;
      99078:data<=16'd22444;
      99079:data<=16'd17673;
      99080:data<=16'd13524;
      99081:data<=16'd16525;
      99082:data<=16'd16680;
      99083:data<=16'd17452;
      99084:data<=16'd18249;
      99085:data<=16'd16892;
      99086:data<=16'd19317;
      99087:data<=16'd13470;
      99088:data<=16'd4026;
      99089:data<=16'd9244;
      99090:data<=16'd14724;
      99091:data<=16'd14427;
      99092:data<=16'd15697;
      99093:data<=16'd13073;
      99094:data<=16'd11664;
      99095:data<=16'd13972;
      99096:data<=16'd16387;
      99097:data<=16'd18773;
      99098:data<=16'd13045;
      99099:data<=16'd8395;
      99100:data<=16'd13609;
      99101:data<=16'd13342;
      99102:data<=16'd9888;
      99103:data<=16'd5656;
      99104:data<=-16'd7080;
      99105:data<=-16'd11773;
      99106:data<=-16'd6975;
      99107:data<=-16'd9365;
      99108:data<=-16'd9730;
      99109:data<=-16'd3428;
      99110:data<=-16'd1447;
      99111:data<=-16'd2311;
      99112:data<=-16'd2009;
      99113:data<=-16'd845;
      99114:data<=16'd1083;
      99115:data<=16'd526;
      99116:data<=-16'd1068;
      99117:data<=16'd541;
      99118:data<=16'd80;
      99119:data<=-16'd3078;
      99120:data<=-16'd640;
      99121:data<=16'd2265;
      99122:data<=16'd194;
      99123:data<=-16'd491;
      99124:data<=-16'd1154;
      99125:data<=-16'd1629;
      99126:data<=-16'd155;
      99127:data<=-16'd1463;
      99128:data<=16'd1151;
      99129:data<=16'd4801;
      99130:data<=16'd115;
      99131:data<=16'd1007;
      99132:data<=16'd3844;
      99133:data<=-16'd2338;
      99134:data<=-16'd535;
      99135:data<=16'd5501;
      99136:data<=16'd3870;
      99137:data<=16'd5066;
      99138:data<=16'd5668;
      99139:data<=16'd2226;
      99140:data<=16'd1365;
      99141:data<=-16'd53;
      99142:data<=-16'd513;
      99143:data<=-16'd537;
      99144:data<=-16'd3641;
      99145:data<=-16'd3541;
      99146:data<=-16'd1233;
      99147:data<=-16'd196;
      99148:data<=16'd2314;
      99149:data<=16'd5914;
      99150:data<=16'd7250;
      99151:data<=16'd3225;
      99152:data<=16'd1304;
      99153:data<=16'd3858;
      99154:data<=16'd1572;
      99155:data<=16'd2863;
      99156:data<=16'd5715;
      99157:data<=-16'd3582;
      99158:data<=-16'd4930;
      99159:data<=16'd5636;
      99160:data<=16'd5242;
      99161:data<=16'd699;
      99162:data<=-16'd1522;
      99163:data<=-16'd4284;
      99164:data<=16'd484;
      99165:data<=16'd4532;
      99166:data<=16'd550;
      99167:data<=-16'd2525;
      99168:data<=-16'd3667;
      99169:data<=-16'd3365;
      99170:data<=-16'd1795;
      99171:data<=16'd1615;
      99172:data<=16'd8399;
      99173:data<=16'd6267;
      99174:data<=-16'd1862;
      99175:data<=16'd2211;
      99176:data<=16'd5137;
      99177:data<=-16'd2290;
      99178:data<=-16'd2848;
      99179:data<=-16'd3794;
      99180:data<=-16'd10881;
      99181:data<=-16'd5086;
      99182:data<=16'd3421;
      99183:data<=-16'd1192;
      99184:data<=-16'd4678;
      99185:data<=-16'd4563;
      99186:data<=-16'd2784;
      99187:data<=16'd3882;
      99188:data<=16'd807;
      99189:data<=-16'd7201;
      99190:data<=-16'd3498;
      99191:data<=-16'd1125;
      99192:data<=-16'd5470;
      99193:data<=-16'd9723;
      99194:data<=-16'd14451;
      99195:data<=-16'd13869;
      99196:data<=-16'd11837;
      99197:data<=-16'd13411;
      99198:data<=-16'd14765;
      99199:data<=-16'd20677;
      99200:data<=-16'd21558;
      99201:data<=-16'd12207;
      99202:data<=-16'd10343;
      99203:data<=-16'd12057;
      99204:data<=-16'd12414;
      99205:data<=-16'd15958;
      99206:data<=-16'd13591;
      99207:data<=-16'd13535;
      99208:data<=-16'd18201;
      99209:data<=-16'd13944;
      99210:data<=-16'd11737;
      99211:data<=-16'd11568;
      99212:data<=-16'd7826;
      99213:data<=-16'd13568;
      99214:data<=-16'd17754;
      99215:data<=-16'd13318;
      99216:data<=-16'd12772;
      99217:data<=-16'd12763;
      99218:data<=-16'd13855;
      99219:data<=-16'd13746;
      99220:data<=-16'd9254;
      99221:data<=-16'd12968;
      99222:data<=-16'd15582;
      99223:data<=-16'd11705;
      99224:data<=-16'd13388;
      99225:data<=-16'd10064;
      99226:data<=-16'd7529;
      99227:data<=-16'd13452;
      99228:data<=-16'd6886;
      99229:data<=-16'd2452;
      99230:data<=-16'd13153;
      99231:data<=-16'd12975;
      99232:data<=-16'd8604;
      99233:data<=-16'd14073;
      99234:data<=-16'd15945;
      99235:data<=-16'd13750;
      99236:data<=-16'd10683;
      99237:data<=-16'd7618;
      99238:data<=-16'd7366;
      99239:data<=-16'd3225;
      99240:data<=-16'd434;
      99241:data<=-16'd4646;
      99242:data<=-16'd6645;
      99243:data<=-16'd9421;
      99244:data<=-16'd11012;
      99245:data<=-16'd3576;
      99246:data<=-16'd1403;
      99247:data<=-16'd5039;
      99248:data<=-16'd513;
      99249:data<=16'd2073;
      99250:data<=-16'd2068;
      99251:data<=-16'd1707;
      99252:data<=16'd258;
      99253:data<=-16'd1979;
      99254:data<=-16'd3021;
      99255:data<=16'd907;
      99256:data<=16'd3342;
      99257:data<=16'd341;
      99258:data<=16'd437;
      99259:data<=16'd4391;
      99260:data<=16'd5655;
      99261:data<=16'd6197;
      99262:data<=16'd4584;
      99263:data<=16'd2611;
      99264:data<=16'd4296;
      99265:data<=16'd2264;
      99266:data<=16'd1989;
      99267:data<=16'd7426;
      99268:data<=16'd6690;
      99269:data<=16'd7630;
      99270:data<=16'd11970;
      99271:data<=16'd7720;
      99272:data<=16'd6123;
      99273:data<=16'd8572;
      99274:data<=16'd7932;
      99275:data<=16'd10731;
      99276:data<=16'd9776;
      99277:data<=16'd6034;
      99278:data<=16'd7289;
      99279:data<=16'd5818;
      99280:data<=16'd8301;
      99281:data<=16'd11447;
      99282:data<=16'd3756;
      99283:data<=16'd3472;
      99284:data<=16'd9297;
      99285:data<=16'd7300;
      99286:data<=16'd7294;
      99287:data<=16'd7470;
      99288:data<=16'd6701;
      99289:data<=16'd9154;
      99290:data<=16'd8516;
      99291:data<=16'd9700;
      99292:data<=16'd10164;
      99293:data<=16'd6777;
      99294:data<=16'd10094;
      99295:data<=16'd10340;
      99296:data<=16'd7169;
      99297:data<=16'd11362;
      99298:data<=16'd10624;
      99299:data<=16'd8646;
      99300:data<=16'd11800;
      99301:data<=16'd9917;
      99302:data<=16'd9356;
      99303:data<=16'd10845;
      99304:data<=16'd12078;
      99305:data<=16'd18189;
      99306:data<=16'd19296;
      99307:data<=16'd18034;
      99308:data<=16'd20051;
      99309:data<=16'd17346;
      99310:data<=16'd17584;
      99311:data<=16'd19135;
      99312:data<=16'd15945;
      99313:data<=16'd17634;
      99314:data<=16'd16496;
      99315:data<=16'd11758;
      99316:data<=16'd14408;
      99317:data<=16'd16211;
      99318:data<=16'd16204;
      99319:data<=16'd15091;
      99320:data<=16'd11094;
      99321:data<=16'd13417;
      99322:data<=16'd14575;
      99323:data<=16'd11947;
      99324:data<=16'd14433;
      99325:data<=16'd12548;
      99326:data<=16'd11938;
      99327:data<=16'd20412;
      99328:data<=16'd22394;
      99329:data<=16'd20635;
      99330:data<=16'd21902;
      99331:data<=16'd20051;
      99332:data<=16'd18698;
      99333:data<=16'd18395;
      99334:data<=16'd17567;
      99335:data<=16'd17632;
      99336:data<=16'd15834;
      99337:data<=16'd15409;
      99338:data<=16'd16384;
      99339:data<=16'd14678;
      99340:data<=16'd13600;
      99341:data<=16'd13238;
      99342:data<=16'd12709;
      99343:data<=16'd12319;
      99344:data<=16'd11183;
      99345:data<=16'd11077;
      99346:data<=16'd9596;
      99347:data<=16'd8595;
      99348:data<=16'd11494;
      99349:data<=16'd10944;
      99350:data<=16'd9145;
      99351:data<=16'd10208;
      99352:data<=16'd8020;
      99353:data<=16'd6343;
      99354:data<=16'd6896;
      99355:data<=16'd5715;
      99356:data<=16'd5281;
      99357:data<=16'd3168;
      99358:data<=16'd1002;
      99359:data<=16'd2980;
      99360:data<=16'd3219;
      99361:data<=16'd2135;
      99362:data<=16'd1466;
      99363:data<=-16'd836;
      99364:data<=-16'd1598;
      99365:data<=-16'd2761;
      99366:data<=-16'd4114;
      99367:data<=-16'd3063;
      99368:data<=-16'd4632;
      99369:data<=-16'd4129;
      99370:data<=-16'd1204;
      99371:data<=-16'd9808;
      99372:data<=-16'd23008;
      99373:data<=-16'd25370;
      99374:data<=-16'd22774;
      99375:data<=-16'd22946;
      99376:data<=-16'd23736;
      99377:data<=-16'd23919;
      99378:data<=-16'd24463;
      99379:data<=-16'd24075;
      99380:data<=-16'd21857;
      99381:data<=-16'd20171;
      99382:data<=-16'd19766;
      99383:data<=-16'd20299;
      99384:data<=-16'd21425;
      99385:data<=-16'd21117;
      99386:data<=-16'd20228;
      99387:data<=-16'd19462;
      99388:data<=-16'd18598;
      99389:data<=-16'd19801;
      99390:data<=-16'd20760;
      99391:data<=-16'd19952;
      99392:data<=-16'd19497;
      99393:data<=-16'd17596;
      99394:data<=-16'd16449;
      99395:data<=-16'd18046;
      99396:data<=-16'd17870;
      99397:data<=-16'd17233;
      99398:data<=-16'd17708;
      99399:data<=-16'd17629;
      99400:data<=-16'd18049;
      99401:data<=-16'd16315;
      99402:data<=-16'd13505;
      99403:data<=-16'd15012;
      99404:data<=-16'd17192;
      99405:data<=-16'd16830;
      99406:data<=-16'd15476;
      99407:data<=-16'd13444;
      99408:data<=-16'd12736;
      99409:data<=-16'd13697;
      99410:data<=-16'd14766;
      99411:data<=-16'd14863;
      99412:data<=-16'd13091;
      99413:data<=-16'd12707;
      99414:data<=-16'd13797;
      99415:data<=-16'd10872;
      99416:data<=-16'd5303;
      99417:data<=-16'd2434;
      99418:data<=-16'd2641;
      99419:data<=-16'd2998;
      99420:data<=-16'd2312;
      99421:data<=-16'd2070;
      99422:data<=-16'd1979;
      99423:data<=-16'd2184;
      99424:data<=-16'd3266;
      99425:data<=-16'd3001;
      99426:data<=-16'd2690;
      99427:data<=-16'd3040;
      99428:data<=-16'd1845;
      99429:data<=-16'd2613;
      99430:data<=-16'd4930;
      99431:data<=-16'd4208;
      99432:data<=-16'd3550;
      99433:data<=-16'd4361;
      99434:data<=-16'd3676;
      99435:data<=-16'd1521;
      99436:data<=-16'd842;
      99437:data<=-16'd3309;
      99438:data<=-16'd1991;
      99439:data<=16'd4364;
      99440:data<=16'd5338;
      99441:data<=16'd3409;
      99442:data<=16'd3917;
      99443:data<=16'd1938;
      99444:data<=16'd981;
      99445:data<=16'd2704;
      99446:data<=16'd1868;
      99447:data<=16'd1791;
      99448:data<=16'd2217;
      99449:data<=16'd323;
      99450:data<=-16'd203;
      99451:data<=-16'd549;
      99452:data<=-16'd970;
      99453:data<=16'd470;
      99454:data<=16'd274;
      99455:data<=16'd153;
      99456:data<=16'd1131;
      99457:data<=-16'd799;
      99458:data<=-16'd520;
      99459:data<=16'd2813;
      99460:data<=-16'd946;
      99461:data<=-16'd9128;
      99462:data<=-16'd11326;
      99463:data<=-16'd9680;
      99464:data<=-16'd9031;
      99465:data<=-16'd7442;
      99466:data<=-16'd5741;
      99467:data<=-16'd6722;
      99468:data<=-16'd7228;
      99469:data<=-16'd5128;
      99470:data<=-16'd3456;
      99471:data<=-16'd2890;
      99472:data<=-16'd2314;
      99473:data<=-16'd2059;
      99474:data<=-16'd1671;
      99475:data<=-16'd884;
      99476:data<=-16'd67;
      99477:data<=16'd643;
      99478:data<=16'd658;
      99479:data<=16'd705;
      99480:data<=16'd1152;
      99481:data<=16'd522;
      99482:data<=16'd832;
      99483:data<=16'd3601;
      99484:data<=16'd4548;
      99485:data<=16'd4153;
      99486:data<=16'd5592;
      99487:data<=16'd4356;
      99488:data<=16'd1783;
      99489:data<=16'd4567;
      99490:data<=16'd6774;
      99491:data<=16'd4731;
      99492:data<=16'd4915;
      99493:data<=16'd5142;
      99494:data<=16'd3257;
      99495:data<=16'd4457;
      99496:data<=16'd6325;
      99497:data<=16'd5953;
      99498:data<=16'd6360;
      99499:data<=16'd6584;
      99500:data<=16'd5714;
      99501:data<=16'd5389;
      99502:data<=16'd5386;
      99503:data<=16'd6692;
      99504:data<=16'd9835;
      99505:data<=16'd11593;
      99506:data<=16'd9990;
      99507:data<=16'd8000;
      99508:data<=16'd8439;
      99509:data<=16'd9244;
      99510:data<=16'd9492;
      99511:data<=16'd10272;
      99512:data<=16'd9796;
      99513:data<=16'd8878;
      99514:data<=16'd8903;
      99515:data<=16'd8117;
      99516:data<=16'd9412;
      99517:data<=16'd12730;
      99518:data<=16'd11920;
      99519:data<=16'd9374;
      99520:data<=16'd8778;
      99521:data<=16'd8187;
      99522:data<=16'd9251;
      99523:data<=16'd10828;
      99524:data<=16'd9444;
      99525:data<=16'd8523;
      99526:data<=16'd9066;
      99527:data<=16'd8551;
      99528:data<=16'd8299;
      99529:data<=16'd8818;
      99530:data<=16'd9418;
      99531:data<=16'd9753;
      99532:data<=16'd9374;
      99533:data<=16'd9438;
      99534:data<=16'd8702;
      99535:data<=16'd7198;
      99536:data<=16'd8937;
      99537:data<=16'd10392;
      99538:data<=16'd8169;
      99539:data<=16'd7746;
      99540:data<=16'd8296;
      99541:data<=16'd7294;
      99542:data<=16'd8554;
      99543:data<=16'd9583;
      99544:data<=16'd8669;
      99545:data<=16'd9341;
      99546:data<=16'd8637;
      99547:data<=16'd6962;
      99548:data<=16'd7879;
      99549:data<=16'd5667;
      99550:data<=-16'd359;
      99551:data<=-16'd3049;
      99552:data<=-16'd2641;
      99553:data<=-16'd2370;
      99554:data<=-16'd1976;
      99555:data<=-16'd767;
      99556:data<=16'd247;
      99557:data<=-16'd149;
      99558:data<=-16'd52;
      99559:data<=16'd698;
      99560:data<=16'd44;
      99561:data<=-16'd111;
      99562:data<=16'd274;
      99563:data<=-16'd643;
      99564:data<=-16'd969;
      99565:data<=-16'd549;
      99566:data<=-16'd443;
      99567:data<=-16'd778;
      99568:data<=-16'd1754;
      99569:data<=-16'd1304;
      99570:data<=-16'd1535;
      99571:data<=-16'd4561;
      99572:data<=-16'd2723;
      99573:data<=16'd4008;
      99574:data<=16'd5703;
      99575:data<=16'd3723;
      99576:data<=16'd3504;
      99577:data<=16'd3139;
      99578:data<=16'd2249;
      99579:data<=16'd2184;
      99580:data<=16'd2226;
      99581:data<=16'd2231;
      99582:data<=16'd1283;
      99583:data<=-16'd1075;
      99584:data<=-16'd1632;
      99585:data<=-16'd243;
      99586:data<=-16'd887;
      99587:data<=-16'd1747;
      99588:data<=-16'd519;
      99589:data<=-16'd1310;
      99590:data<=-16'd3033;
      99591:data<=-16'd1836;
      99592:data<=-16'd1569;
      99593:data<=-16'd2529;
      99594:data<=16'd863;
      99595:data<=16'd6299;
      99596:data<=16'd7468;
      99597:data<=16'd5515;
      99598:data<=16'd4431;
      99599:data<=16'd3639;
      99600:data<=16'd3257;
      99601:data<=16'd4520;
      99602:data<=16'd3615;
      99603:data<=16'd631;
      99604:data<=16'd699;
      99605:data<=16'd1592;
      99606:data<=16'd1149;
      99607:data<=16'd1216;
      99608:data<=-16'd176;
      99609:data<=-16'd1911;
      99610:data<=-16'd1309;
      99611:data<=-16'd949;
      99612:data<=-16'd1369;
      99613:data<=-16'd1574;
      99614:data<=-16'd1630;
      99615:data<=-16'd1663;
      99616:data<=-16'd3536;
      99617:data<=-16'd5071;
      99618:data<=-16'd4005;
      99619:data<=-16'd3973;
      99620:data<=-16'd3964;
      99621:data<=-16'd2619;
      99622:data<=-16'd3921;
      99623:data<=-16'd5689;
      99624:data<=-16'd5009;
      99625:data<=-16'd4683;
      99626:data<=-16'd4722;
      99627:data<=-16'd4404;
      99628:data<=-16'd4731;
      99629:data<=-16'd5550;
      99630:data<=-16'd6613;
      99631:data<=-16'd6913;
      99632:data<=-16'd6957;
      99633:data<=-16'd7696;
      99634:data<=-16'd6579;
      99635:data<=-16'd5691;
      99636:data<=-16'd8511;
      99637:data<=-16'd9163;
      99638:data<=-16'd8235;
      99639:data<=-16'd15571;
      99640:data<=-16'd24965;
      99641:data<=-16'd24932;
      99642:data<=-16'd22944;
      99643:data<=-16'd25062;
      99644:data<=-16'd24501;
      99645:data<=-16'd21946;
      99646:data<=-16'd21490;
      99647:data<=-16'd20319;
      99648:data<=-16'd19373;
      99649:data<=-16'd20688;
      99650:data<=-16'd20797;
      99651:data<=-16'd19180;
      99652:data<=-16'd18154;
      99653:data<=-16'd17496;
      99654:data<=-16'd16745;
      99655:data<=-16'd16409;
      99656:data<=-16'd16536;
      99657:data<=-16'd16083;
      99658:data<=-16'd14979;
      99659:data<=-16'd14425;
      99660:data<=-16'd13749;
      99661:data<=-16'd13168;
      99662:data<=-16'd14225;
      99663:data<=-16'd14692;
      99664:data<=-16'd12930;
      99665:data<=-16'd11276;
      99666:data<=-16'd10718;
      99667:data<=-16'd10762;
      99668:data<=-16'd10925;
      99669:data<=-16'd10266;
      99670:data<=-16'd9232;
      99671:data<=-16'd8783;
      99672:data<=-16'd8859;
      99673:data<=-16'd8918;
      99674:data<=-16'd7592;
      99675:data<=-16'd4990;
      99676:data<=-16'd3383;
      99677:data<=-16'd3125;
      99678:data<=-16'd3189;
      99679:data<=-16'd3046;
      99680:data<=-16'd1880;
      99681:data<=-16'd1398;
      99682:data<=-16'd1999;
      99683:data<=16'd2176;
      99684:data<=16'd9985;
      99685:data<=16'd12242;
      99686:data<=16'd10416;
      99687:data<=16'd10310;
      99688:data<=16'd10499;
      99689:data<=16'd11318;
      99690:data<=16'd12656;
      99691:data<=16'd12213;
      99692:data<=16'd12422;
      99693:data<=16'd12750;
      99694:data<=16'd11195;
      99695:data<=16'd11345;
      99696:data<=16'd12607;
      99697:data<=16'd12190;
      99698:data<=16'd11532;
      99699:data<=16'd11012;
      99700:data<=16'd11141;
      99701:data<=16'd11373;
      99702:data<=16'd10499;
      99703:data<=16'd11479;
      99704:data<=16'd12624;
      99705:data<=16'd11213;
      99706:data<=16'd13051;
      99707:data<=16'd17594;
      99708:data<=16'd18682;
      99709:data<=16'd18885;
      99710:data<=16'd19688;
      99711:data<=16'd18445;
      99712:data<=16'd17105;
      99713:data<=16'd16750;
      99714:data<=16'd16069;
      99715:data<=16'd16028;
      99716:data<=16'd16769;
      99717:data<=16'd16962;
      99718:data<=16'd16202;
      99719:data<=16'd14882;
      99720:data<=16'd14275;
      99721:data<=16'd14519;
      99722:data<=16'd14512;
      99723:data<=16'd14783;
      99724:data<=16'd14751;
      99725:data<=16'd13435;
      99726:data<=16'd13059;
      99727:data<=16'd11626;
      99728:data<=16'd5829;
      99729:data<=16'd2135;
      99730:data<=16'd3624;
      99731:data<=16'd3674;
      99732:data<=16'd2144;
      99733:data<=16'd2132;
      99734:data<=16'd1723;
      99735:data<=16'd1563;
      99736:data<=16'd2961;
      99737:data<=16'd3626;
      99738:data<=16'd3168;
      99739:data<=16'd3213;
      99740:data<=16'd3432;
      99741:data<=16'd3055;
      99742:data<=16'd3430;
      99743:data<=16'd4505;
      99744:data<=16'd4446;
      99745:data<=16'd4347;
      99746:data<=16'd4332;
      99747:data<=16'd3482;
      99748:data<=16'd4407;
      99749:data<=16'd5864;
      99750:data<=16'd4699;
      99751:data<=16'd3906;
      99752:data<=16'd4538;
      99753:data<=16'd4325;
      99754:data<=16'd3870;
      99755:data<=16'd4087;
      99756:data<=16'd4761;
      99757:data<=16'd4969;
      99758:data<=16'd4441;
      99759:data<=16'd4040;
      99760:data<=16'd3451;
      99761:data<=16'd3300;
      99762:data<=16'd3811;
      99763:data<=16'd3560;
      99764:data<=16'd3395;
      99765:data<=16'd3751;
      99766:data<=16'd4135;
      99767:data<=16'd4161;
      99768:data<=16'd3701;
      99769:data<=16'd5395;
      99770:data<=16'd5680;
      99771:data<=16'd2326;
      99772:data<=16'd6109;
      99773:data<=16'd12419;
      99774:data<=16'd7876;
      99775:data<=16'd3421;
      99776:data<=16'd5045;
      99777:data<=16'd3723;
      99778:data<=16'd2734;
      99779:data<=16'd3835;
      99780:data<=16'd2992;
      99781:data<=16'd2155;
      99782:data<=16'd872;
      99783:data<=16'd35;
      99784:data<=16'd769;
      99785:data<=-16'd370;
      99786:data<=-16'd1089;
      99787:data<=-16'd549;
      99788:data<=-16'd2159;
      99789:data<=-16'd3636;
      99790:data<=-16'd4146;
      99791:data<=-16'd4799;
      99792:data<=-16'd4576;
      99793:data<=-16'd4259;
      99794:data<=-16'd4027;
      99795:data<=-16'd4775;
      99796:data<=-16'd6943;
      99797:data<=-16'd7407;
      99798:data<=-16'd6792;
      99799:data<=-16'd6660;
      99800:data<=-16'd5749;
      99801:data<=-16'd5721;
      99802:data<=-16'd7465;
      99803:data<=-16'd8743;
      99804:data<=-16'd8081;
      99805:data<=-16'd6517;
      99806:data<=-16'd6646;
      99807:data<=-16'd7244;
      99808:data<=-16'd6989;
      99809:data<=-16'd7896;
      99810:data<=-16'd8557;
      99811:data<=-16'd8199;
      99812:data<=-16'd8129;
      99813:data<=-16'd7655;
      99814:data<=-16'd8454;
      99815:data<=-16'd9447;
      99816:data<=-16'd8997;
      99817:data<=-16'd12974;
      99818:data<=-16'd19083;
      99819:data<=-16'd19036;
      99820:data<=-16'd17073;
      99821:data<=-16'd17942;
      99822:data<=-16'd18492;
      99823:data<=-16'd17975;
      99824:data<=-16'd17755;
      99825:data<=-16'd17634;
      99826:data<=-16'd16768;
      99827:data<=-16'd15869;
      99828:data<=-16'd16404;
      99829:data<=-16'd17053;
      99830:data<=-16'd16725;
      99831:data<=-16'd16105;
      99832:data<=-16'd15206;
      99833:data<=-16'd14314;
      99834:data<=-16'd13756;
      99835:data<=-16'd14366;
      99836:data<=-16'd15396;
      99837:data<=-16'd14001;
      99838:data<=-16'd12983;
      99839:data<=-16'd13778;
      99840:data<=-16'd10222;
      99841:data<=-16'd4748;
      99842:data<=-16'd4494;
      99843:data<=-16'd5447;
      99844:data<=-16'd4249;
      99845:data<=-16'd4306;
      99846:data<=-16'd4649;
      99847:data<=-16'd3313;
      99848:data<=-16'd3344;
      99849:data<=-16'd5171;
      99850:data<=-16'd5541;
      99851:data<=-16'd5259;
      99852:data<=-16'd5598;
      99853:data<=-16'd4808;
      99854:data<=-16'd4508;
      99855:data<=-16'd5709;
      99856:data<=-16'd5641;
      99857:data<=-16'd4928;
      99858:data<=-16'd4434;
      99859:data<=-16'd3902;
      99860:data<=-16'd4466;
      99861:data<=-16'd2652;
      99862:data<=16'd2757;
      99863:data<=16'd5338;
      99864:data<=16'd4410;
      99865:data<=16'd4109;
      99866:data<=16'd4334;
      99867:data<=16'd4191;
      99868:data<=16'd3542;
      99869:data<=16'd2849;
      99870:data<=16'd2869;
      99871:data<=16'd2689;
      99872:data<=16'd2485;
      99873:data<=16'd2881;
      99874:data<=16'd2381;
      99875:data<=16'd834;
      99876:data<=16'd194;
      99877:data<=16'd920;
      99878:data<=16'd999;
      99879:data<=-16'd94;
      99880:data<=-16'd62;
      99881:data<=16'd1004;
      99882:data<=16'd1307;
      99883:data<=16'd1045;
      99884:data<=16'd731;
      99885:data<=16'd1107;
      99886:data<=16'd1486;
      99887:data<=16'd716;
      99888:data<=16'd1580;
      99889:data<=16'd3827;
      99890:data<=16'd3902;
      99891:data<=16'd3748;
      99892:data<=16'd3902;
      99893:data<=16'd2519;
      99894:data<=16'd2911;
      99895:data<=16'd5313;
      99896:data<=16'd6081;
      99897:data<=16'd5702;
      99898:data<=16'd5163;
      99899:data<=16'd4807;
      99900:data<=16'd4968;
      99901:data<=16'd5216;
      99902:data<=16'd6598;
      99903:data<=16'd7216;
      99904:data<=16'd5761;
      99905:data<=16'd6326;
      99906:data<=16'd4454;
      99907:data<=-16'd5301;
      99908:data<=-16'd12016;
      99909:data<=-16'd10387;
      99910:data<=-16'd9163;
      99911:data<=-16'd9200;
      99912:data<=-16'd8272;
      99913:data<=-16'd8845;
      99914:data<=-16'd8572;
      99915:data<=-16'd6032;
      99916:data<=-16'd4868;
      99917:data<=-16'd5297;
      99918:data<=-16'd5162;
      99919:data<=-16'd4223;
      99920:data<=-16'd3618;
      99921:data<=-16'd3430;
      99922:data<=-16'd2140;
      99923:data<=-16'd775;
      99924:data<=-16'd726;
      99925:data<=-16'd611;
      99926:data<=-16'd661;
      99927:data<=-16'd441;
      99928:data<=16'd1624;
      99929:data<=16'd2761;
      99930:data<=16'd2140;
      99931:data<=16'd2629;
      99932:data<=16'd3062;
      99933:data<=16'd2499;
      99934:data<=16'd3224;
      99935:data<=16'd5034;
      99936:data<=16'd6070;
      99937:data<=16'd5935;
      99938:data<=16'd5815;
      99939:data<=16'd6244;
      99940:data<=16'd5959;
      99941:data<=16'd5984;
      99942:data<=16'd7313;
      99943:data<=16'd7527;
      99944:data<=16'd7194;
      99945:data<=16'd7570;
      99946:data<=16'd6630;
      99947:data<=16'd6293;
      99948:data<=16'd7747;
      99949:data<=16'd7535;
      99950:data<=16'd8975;
      99951:data<=16'd15191;
      99952:data<=16'd18692;
      99953:data<=16'd17261;
      99954:data<=16'd17206;
      99955:data<=16'd18120;
      99956:data<=16'd17200;
      99957:data<=16'd16803;
      99958:data<=16'd17077;
      99959:data<=16'd16010;
      99960:data<=16'd14797;
      99961:data<=16'd14827;
      99962:data<=16'd15628;
      99963:data<=16'd16004;
      99964:data<=16'd14959;
      99965:data<=16'd13664;
      99966:data<=16'd13115;
      99967:data<=16'd12734;
      99968:data<=16'd13433;
      99969:data<=16'd13941;
      99970:data<=16'd12342;
      99971:data<=16'd12483;
      99972:data<=16'd13524;
      99973:data<=16'd11358;
      99974:data<=16'd13232;
      99975:data<=16'd20415;
      99976:data<=16'd21601;
      99977:data<=16'd18862;
      99978:data<=16'd19323;
      99979:data<=16'd18512;
      99980:data<=16'd16345;
      99981:data<=16'd16604;
      99982:data<=16'd16956;
      99983:data<=16'd16352;
      99984:data<=16'd15438;
      99985:data<=16'd14668;
      99986:data<=16'd14677;
      99987:data<=16'd13729;
      99988:data<=16'd12125;
      99989:data<=16'd11430;
      99990:data<=16'd11035;
      99991:data<=16'd11004;
      99992:data<=16'd10433;
      99993:data<=16'd10055;
      99994:data<=16'd10329;
      99995:data<=16'd5234;
      99996:data<=-16'd2927;
      99997:data<=-16'd4927;
      99998:data<=-16'd4226;
      99999:data<=-16'd4810;
      100000:data<=-16'd4106;
      100001:data<=-16'd4611;
      100002:data<=-16'd6269;
      100003:data<=-16'd6307;
      100004:data<=-16'd6837;
      100005:data<=-16'd7339;
      100006:data<=-16'd6434;
      100007:data<=-16'd6388;
      100008:data<=-16'd7621;
      100009:data<=-16'd8573;
      100010:data<=-16'd8111;
      100011:data<=-16'd7423;
      100012:data<=-16'd7970;
      100013:data<=-16'd7891;
      100014:data<=-16'd7794;
      100015:data<=-16'd9570;
      100016:data<=-16'd10436;
      100017:data<=-16'd9629;
      100018:data<=-16'd9323;
      100019:data<=-16'd9169;
      100020:data<=-16'd8921;
      100021:data<=-16'd9259;
      100022:data<=-16'd10049;
      100023:data<=-16'd10477;
      100024:data<=-16'd9721;
      100025:data<=-16'd8589;
      100026:data<=-16'd8473;
      100027:data<=-16'd9386;
      100028:data<=-16'd10207;
      100029:data<=-16'd10217;
      100030:data<=-16'd9988;
      100031:data<=-16'd9515;
      100032:data<=-16'd8813;
      100033:data<=-16'd8634;
      100034:data<=-16'd8974;
      100035:data<=-16'd10249;
      100036:data<=-16'd10725;
      100037:data<=-16'd9389;
      100038:data<=-16'd10534;
      100039:data<=-16'd10246;
      100040:data<=-16'd3283;
      100041:data<=-16'd1556;
      100042:data<=-16'd8313;
      100043:data<=-16'd10213;
      100044:data<=-16'd8363;
      100045:data<=-16'd9163;
      100046:data<=-16'd8880;
      100047:data<=-16'd8534;
      100048:data<=-16'd10161;
      100049:data<=-16'd10302;
      100050:data<=-16'd9268;
      100051:data<=-16'd8696;
      100052:data<=-16'd7964;
      100053:data<=-16'd7539;
      100054:data<=-16'd7806;
      100055:data<=-16'd8210;
      100056:data<=-16'd8617;
      100057:data<=-16'd9168;
      100058:data<=-16'd9166;
      100059:data<=-16'd8194;
      100060:data<=-16'd7717;
      100061:data<=-16'd8325;
      100062:data<=-16'd8614;
      100063:data<=-16'd8128;
      100064:data<=-16'd7677;
      100065:data<=-16'd7318;
      100066:data<=-16'd6511;
      100067:data<=-16'd6522;
      100068:data<=-16'd7818;
      100069:data<=-16'd7849;
      100070:data<=-16'd7178;
      100071:data<=-16'd7514;
      100072:data<=-16'd6658;
      100073:data<=-16'd5221;
      100074:data<=-16'd5770;
      100075:data<=-16'd7122;
      100076:data<=-16'd7612;
      100077:data<=-16'd6796;
      100078:data<=-16'd5953;
      100079:data<=-16'd5544;
      100080:data<=-16'd4487;
      100081:data<=-16'd5523;
      100082:data<=-16'd7110;
      100083:data<=-16'd5218;
      100084:data<=-16'd7556;
      100085:data<=-16'd15168;
      100086:data<=-16'd16847;
      100087:data<=-16'd15158;
      100088:data<=-16'd16392;
      100089:data<=-16'd16245;
      100090:data<=-16'd14600;
      100091:data<=-16'd13844;
      100092:data<=-16'd12925;
      100093:data<=-16'd12123;
      100094:data<=-16'd11544;
      100095:data<=-16'd11505;
      100096:data<=-16'd11388;
      100097:data<=-16'd9803;
      100098:data<=-16'd9007;
      100099:data<=-16'd9133;
      100100:data<=-16'd7884;
      100101:data<=-16'd6214;
      100102:data<=-16'd4949;
      100103:data<=-16'd4813;
      100104:data<=-16'd5042;
      100105:data<=-16'd3483;
      100106:data<=-16'd3127;
      100107:data<=-16'd3371;
      100108:data<=16'd1365;
      100109:data<=16'd7097;
      100110:data<=16'd8493;
      100111:data<=16'd8476;
      100112:data<=16'd8617;
      100113:data<=16'd8486;
      100114:data<=16'd9222;
      100115:data<=16'd10316;
      100116:data<=16'd10198;
      100117:data<=16'd9589;
      100118:data<=16'd9667;
      100119:data<=16'd8840;
      100120:data<=16'd7955;
      100121:data<=16'd9743;
      100122:data<=16'd10725;
      100123:data<=16'd9338;
      100124:data<=16'd9166;
      100125:data<=16'd9215;
      100126:data<=16'd9078;
      100127:data<=16'd9597;
      100128:data<=16'd9506;
      100129:data<=16'd12927;
      100130:data<=16'd19575;
      100131:data<=16'd21196;
      100132:data<=16'd19159;
      100133:data<=16'd18859;
      100134:data<=16'd19255;
      100135:data<=16'd19343;
      100136:data<=16'd18906;
      100137:data<=16'd18647;
      100138:data<=16'd18888;
      100139:data<=16'd17538;
      100140:data<=16'd16557;
      100141:data<=16'd17796;
      100142:data<=16'd17932;
      100143:data<=16'd16760;
      100144:data<=16'd16160;
      100145:data<=16'd15309;
      100146:data<=16'd14383;
      100147:data<=16'd14794;
      100148:data<=16'd16152;
      100149:data<=16'd16190;
      100150:data<=16'd14748;
      100151:data<=16'd14317;
      100152:data<=16'd14390;
      100153:data<=16'd13594;
      100154:data<=16'd13635;
      100155:data<=16'd14242;
      100156:data<=16'd13179;
      100157:data<=16'd11765;
      100158:data<=16'd11958;
      100159:data<=16'd11885;
      100160:data<=16'd11053;
      100161:data<=16'd11775;
      100162:data<=16'd12182;
      100163:data<=16'd10727;
      100164:data<=16'd10624;
      100165:data<=16'd11136;
      100166:data<=16'd10158;
      100167:data<=16'd10031;
      100168:data<=16'd10880;
      100169:data<=16'd10937;
      100170:data<=16'd10426;
      100171:data<=16'd10091;
      100172:data<=16'd9806;
      100173:data<=16'd7277;
      100174:data<=16'd2200;
      100175:data<=-16'd3140;
      100176:data<=-16'd8015;
      100177:data<=-16'd9888;
      100178:data<=-16'd8496;
      100179:data<=-16'd8410;
      100180:data<=-16'd8734;
      100181:data<=-16'd7277;
      100182:data<=-16'd6440;
      100183:data<=-16'd6261;
      100184:data<=-16'd5753;
      100185:data<=-16'd5383;
      100186:data<=-16'd5532;
      100187:data<=-16'd5796;
      100188:data<=-16'd4156;
      100189:data<=-16'd2393;
      100190:data<=-16'd3162;
      100191:data<=-16'd3588;
      100192:data<=-16'd3331;
      100193:data<=-16'd3597;
      100194:data<=-16'd2504;
      100195:data<=-16'd1383;
      100196:data<=-16'd1612;
      100197:data<=-16'd1930;
      100198:data<=-16'd2090;
      100199:data<=-16'd1842;
      100200:data<=-16'd1959;
      100201:data<=-16'd2347;
      100202:data<=-16'd2147;
      100203:data<=-16'd2658;
      100204:data<=-16'd2619;
      100205:data<=-16'd1867;
      100206:data<=-16'd2629;
      100207:data<=-16'd2716;
      100208:data<=-16'd2877;
      100209:data<=-16'd4563;
      100210:data<=-16'd4181;
      100211:data<=-16'd3500;
      100212:data<=-16'd3855;
      100213:data<=-16'd3365;
      100214:data<=-16'd4954;
      100215:data<=-16'd6366;
      100216:data<=-16'd5548;
      100217:data<=-16'd6401;
      100218:data<=-16'd3618;
      100219:data<=16'd3501;
      100220:data<=16'd4516;
      100221:data<=16'd1950;
      100222:data<=16'd2455;
      100223:data<=16'd2617;
      100224:data<=16'd1845;
      100225:data<=16'd1983;
      100226:data<=16'd1462;
      100227:data<=16'd42;
      100228:data<=-16'd1005;
      100229:data<=-16'd1298;
      100230:data<=-16'd978;
      100231:data<=16'd67;
      100232:data<=16'd1011;
      100233:data<=16'd426;
      100234:data<=-16'd795;
      100235:data<=-16'd1131;
      100236:data<=-16'd743;
      100237:data<=-16'd901;
      100238:data<=-16'd1994;
      100239:data<=-16'd2006;
      100240:data<=-16'd1956;
      100241:data<=-16'd3474;
      100242:data<=-16'd1892;
      100243:data<=16'd2168;
      100244:data<=16'd2531;
      100245:data<=16'd1563;
      100246:data<=16'd1741;
      100247:data<=16'd600;
      100248:data<=-16'd614;
      100249:data<=-16'd892;
      100250:data<=-16'd1095;
      100251:data<=-16'd890;
      100252:data<=-16'd931;
      100253:data<=-16'd1500;
      100254:data<=-16'd2473;
      100255:data<=-16'd3513;
      100256:data<=-16'd3494;
      100257:data<=-16'd3383;
      100258:data<=-16'd3433;
      100259:data<=-16'd3068;
      100260:data<=-16'd3750;
      100261:data<=-16'd4476;
      100262:data<=-16'd5520;
      100263:data<=-16'd9838;
      100264:data<=-16'd13342;
      100265:data<=-16'd12381;
      100266:data<=-16'd11873;
      100267:data<=-16'd13470;
      100268:data<=-16'd13652;
      100269:data<=-16'd12786;
      100270:data<=-16'd12951;
      100271:data<=-16'd12956;
      100272:data<=-16'd11919;
      100273:data<=-16'd11879;
      100274:data<=-16'd12756;
      100275:data<=-16'd12539;
      100276:data<=-16'd12202;
      100277:data<=-16'd12290;
      100278:data<=-16'd11509;
      100279:data<=-16'd10618;
      100280:data<=-16'd10772;
      100281:data<=-16'd11685;
      100282:data<=-16'd12070;
      100283:data<=-16'd11122;
      100284:data<=-16'd10292;
      100285:data<=-16'd10070;
      100286:data<=-16'd9749;
      100287:data<=-16'd10287;
      100288:data<=-16'd11209;
      100289:data<=-16'd10830;
      100290:data<=-16'd9737;
      100291:data<=-16'd9083;
      100292:data<=-16'd8887;
      100293:data<=-16'd8467;
      100294:data<=-16'd8334;
      100295:data<=-16'd9333;
      100296:data<=-16'd9873;
      100297:data<=-16'd9412;
      100298:data<=-16'd8768;
      100299:data<=-16'd7896;
      100300:data<=-16'd8531;
      100301:data<=-16'd9809;
      100302:data<=-16'd9041;
      100303:data<=-16'd8661;
      100304:data<=-16'd8502;
      100305:data<=-16'd7163;
      100306:data<=-16'd7564;
      100307:data<=-16'd5278;
      100308:data<=16'd1312;
      100309:data<=16'd1256;
      100310:data<=-16'd4015;
      100311:data<=-16'd4270;
      100312:data<=-16'd2793;
      100313:data<=-16'd2667;
      100314:data<=-16'd1011;
      100315:data<=-16'd232;
      100316:data<=-16'd1046;
      100317:data<=-16'd734;
      100318:data<=-16'd235;
      100319:data<=16'd53;
      100320:data<=16'd1340;
      100321:data<=16'd2390;
      100322:data<=16'd2417;
      100323:data<=16'd2778;
      100324:data<=16'd3172;
      100325:data<=16'd2516;
      100326:data<=16'd2594;
      100327:data<=16'd4385;
      100328:data<=16'd5529;
      100329:data<=16'd5216;
      100330:data<=16'd4710;
      100331:data<=16'd4290;
      100332:data<=16'd4313;
      100333:data<=16'd5432;
      100334:data<=16'd6664;
      100335:data<=16'd6563;
      100336:data<=16'd6176;
      100337:data<=16'd6608;
      100338:data<=16'd6361;
      100339:data<=16'd5949;
      100340:data<=16'd7142;
      100341:data<=16'd8207;
      100342:data<=16'd8296;
      100343:data<=16'd8448;
      100344:data<=16'd8137;
      100345:data<=16'd7686;
      100346:data<=16'd7887;
      100347:data<=16'd8674;
      100348:data<=16'd9429;
      100349:data<=16'd8784;
      100350:data<=16'd8713;
      100351:data<=16'd9470;
      100352:data<=16'd5533;
      100353:data<=16'd287;
      100354:data<=16'd1298;
      100355:data<=16'd3254;
      100356:data<=16'd2103;
      100357:data<=16'd2332;
      100358:data<=16'd3013;
      100359:data<=16'd2637;
      100360:data<=16'd3789;
      100361:data<=16'd5078;
      100362:data<=16'd4884;
      100363:data<=16'd4896;
      100364:data<=16'd5145;
      100365:data<=16'd4840;
      100366:data<=16'd4868;
      100367:data<=16'd5780;
      100368:data<=16'd6279;
      100369:data<=16'd6034;
      100370:data<=16'd6510;
      100371:data<=16'd6811;
      100372:data<=16'd6235;
      100373:data<=16'd6895;
      100374:data<=16'd7890;
      100375:data<=16'd8260;
      100376:data<=16'd10709;
      100377:data<=16'd13624;
      100378:data<=16'd13615;
      100379:data<=16'd13147;
      100380:data<=16'd14108;
      100381:data<=16'd14498;
      100382:data<=16'd13875;
      100383:data<=16'd13550;
      100384:data<=16'd13458;
      100385:data<=16'd12754;
      100386:data<=16'd12499;
      100387:data<=16'd13506;
      100388:data<=16'd13661;
      100389:data<=16'd12654;
      100390:data<=16'd12377;
      100391:data<=16'd11867;
      100392:data<=16'd11015;
      100393:data<=16'd12122;
      100394:data<=16'd13192;
      100395:data<=16'd12066;
      100396:data<=16'd13329;
      100397:data<=16'd18119;
      100398:data<=16'd19920;
      100399:data<=16'd18516;
      100400:data<=16'd18777;
      100401:data<=16'd19067;
      100402:data<=16'd18019;
      100403:data<=16'd17878;
      100404:data<=16'd17324;
      100405:data<=16'd15904;
      100406:data<=16'd15826;
      100407:data<=16'd16213;
      100408:data<=16'd15819;
      100409:data<=16'd15115;
      100410:data<=16'd14284;
      100411:data<=16'd13606;
      100412:data<=16'd13077;
      100413:data<=16'd12505;
      100414:data<=16'd11808;
      100415:data<=16'd10919;
      100416:data<=16'd10329;
      100417:data<=16'd9976;
      100418:data<=16'd9470;
      100419:data<=16'd8472;
      100420:data<=16'd6546;
      100421:data<=16'd5010;
      100422:data<=16'd4799;
      100423:data<=16'd4772;
      100424:data<=16'd4607;
      100425:data<=16'd4181;
      100426:data<=16'd3148;
      100427:data<=16'd1804;
      100428:data<=16'd528;
      100429:data<=16'd111;
      100430:data<=-16'd124;
      100431:data<=-16'd789;
      100432:data<=-16'd796;
      100433:data<=-16'd1809;
      100434:data<=-16'd4026;
      100435:data<=-16'd4223;
      100436:data<=-16'd3529;
      100437:data<=-16'd3650;
      100438:data<=-16'd3880;
      100439:data<=-16'd4531;
      100440:data<=-16'd5325;
      100441:data<=-16'd8313;
      100442:data<=-16'd14372;
      100443:data<=-16'd18336;
      100444:data<=-16'd19306;
      100445:data<=-16'd19764;
      100446:data<=-16'd19560;
      100447:data<=-16'd20107;
      100448:data<=-16'd20615;
      100449:data<=-16'd19585;
      100450:data<=-16'd19233;
      100451:data<=-16'd18753;
      100452:data<=-16'd17834;
      100453:data<=-16'd18638;
      100454:data<=-16'd19244;
      100455:data<=-16'd18835;
      100456:data<=-16'd18633;
      100457:data<=-16'd17893;
      100458:data<=-16'd17291;
      100459:data<=-16'd17417;
      100460:data<=-16'd17421;
      100461:data<=-16'd17103;
      100462:data<=-16'd16480;
      100463:data<=-16'd16334;
      100464:data<=-16'd16261;
      100465:data<=-16'd15315;
      100466:data<=-16'd15194;
      100467:data<=-16'd16117;
      100468:data<=-16'd16116;
      100469:data<=-16'd15256;
      100470:data<=-16'd14763;
      100471:data<=-16'd14684;
      100472:data<=-16'd14258;
      100473:data<=-16'd14311;
      100474:data<=-16'd15127;
      100475:data<=-16'd14669;
      100476:data<=-16'd13587;
      100477:data<=-16'd13079;
      100478:data<=-16'd12260;
      100479:data<=-16'd12357;
      100480:data<=-16'd13280;
      100481:data<=-16'd13077;
      100482:data<=-16'd12383;
      100483:data<=-16'd11943;
      100484:data<=-16'd11571;
      100485:data<=-16'd9250;
      100486:data<=-16'd4375;
      100487:data<=-16'd2238;
      100488:data<=-16'd3275;
      100489:data<=-16'd2684;
      100490:data<=-16'd1912;
      100491:data<=-16'd2314;
      100492:data<=-16'd2370;
      100493:data<=-16'd3054;
      100494:data<=-16'd3912;
      100495:data<=-16'd3800;
      100496:data<=-16'd3341;
      100497:data<=-16'd2776;
      100498:data<=-16'd2440;
      100499:data<=-16'd2602;
      100500:data<=-16'd3454;
      100501:data<=-16'd4255;
      100502:data<=-16'd4088;
      100503:data<=-16'd4190;
      100504:data<=-16'd3777;
      100505:data<=-16'd2490;
      100506:data<=-16'd3394;
      100507:data<=-16'd5131;
      100508:data<=-16'd5300;
      100509:data<=-16'd4193;
      100510:data<=-16'd473;
      100511:data<=16'd2999;
      100512:data<=16'd2426;
      100513:data<=16'd931;
      100514:data<=16'd597;
      100515:data<=16'd605;
      100516:data<=16'd719;
      100517:data<=16'd506;
      100518:data<=16'd550;
      100519:data<=16'd682;
      100520:data<=16'd623;
      100521:data<=16'd860;
      100522:data<=16'd546;
      100523:data<=16'd435;
      100524:data<=16'd611;
      100525:data<=16'd230;
      100526:data<=16'd1563;
      100527:data<=16'd3081;
      100528:data<=16'd2854;
      100529:data<=16'd3418;
      100530:data<=16'd1413;
      100531:data<=-16'd4102;
      100532:data<=-16'd5277;
      100533:data<=-16'd2547;
      100534:data<=-16'd1886;
      100535:data<=-16'd2491;
      100536:data<=-16'd2362;
      100537:data<=-16'd1997;
      100538:data<=-16'd1629;
      100539:data<=-16'd450;
      100540:data<=16'd1090;
      100541:data<=16'd1204;
      100542:data<=16'd917;
      100543:data<=16'd1303;
      100544:data<=16'd1066;
      100545:data<=16'd937;
      100546:data<=16'd2173;
      100547:data<=16'd3867;
      100548:data<=16'd4578;
      100549:data<=16'd4176;
      100550:data<=16'd4065;
      100551:data<=16'd4170;
      100552:data<=16'd4379;
      100553:data<=16'd5603;
      100554:data<=16'd5835;
      100555:data<=16'd4745;
      100556:data<=16'd4789;
      100557:data<=16'd5068;
      100558:data<=16'd5216;
      100559:data<=16'd5970;
      100560:data<=16'd6120;
      100561:data<=16'd6507;
      100562:data<=16'd7395;
      100563:data<=16'd7312;
      100564:data<=16'd7147;
      100565:data<=16'd7250;
      100566:data<=16'd7696;
      100567:data<=16'd8845;
      100568:data<=16'd8969;
      100569:data<=16'd8569;
      100570:data<=16'd8593;
      100571:data<=16'd8049;
      100572:data<=16'd8748;
      100573:data<=16'd9943;
      100574:data<=16'd9864;
      100575:data<=16'd13182;
      100576:data<=16'd17221;
      100577:data<=16'd13759;
      100578:data<=16'd9153;
      100579:data<=16'd10472;
      100580:data<=16'd11899;
      100581:data<=16'd11364;
      100582:data<=16'd11514;
      100583:data<=16'd10937;
      100584:data<=16'd9993;
      100585:data<=16'd10469;
      100586:data<=16'd11550;
      100587:data<=16'd12093;
      100588:data<=16'd11703;
      100589:data<=16'd11235;
      100590:data<=16'd10931;
      100591:data<=16'd10009;
      100592:data<=16'd9906;
      100593:data<=16'd11069;
      100594:data<=16'd11306;
      100595:data<=16'd10504;
      100596:data<=16'd9876;
      100597:data<=16'd9257;
      100598:data<=16'd8395;
      100599:data<=16'd8587;
      100600:data<=16'd10219;
      100601:data<=16'd10473;
      100602:data<=16'd9171;
      100603:data<=16'd8856;
      100604:data<=16'd8249;
      100605:data<=16'd7385;
      100606:data<=16'd8557;
      100607:data<=16'd9351;
      100608:data<=16'd8426;
      100609:data<=16'd8135;
      100610:data<=16'd8061;
      100611:data<=16'd7544;
      100612:data<=16'd7803;
      100613:data<=16'd8111;
      100614:data<=16'd7617;
      100615:data<=16'd7483;
      100616:data<=16'd7244;
      100617:data<=16'd6205;
      100618:data<=16'd6354;
      100619:data<=16'd5756;
      100620:data<=16'd1357;
      100621:data<=-16'd1783;
      100622:data<=-16'd1145;
      100623:data<=-16'd977;
      100624:data<=-16'd1175;
      100625:data<=-16'd1149;
      100626:data<=-16'd1968;
      100627:data<=-16'd2059;
      100628:data<=-16'd2056;
      100629:data<=-16'd2557;
      100630:data<=-16'd2284;
      100631:data<=-16'd2355;
      100632:data<=-16'd3186;
      100633:data<=-16'd4636;
      100634:data<=-16'd5967;
      100635:data<=-16'd5362;
      100636:data<=-16'd4981;
      100637:data<=-16'd5533;
      100638:data<=-16'd5327;
      100639:data<=-16'd6399;
      100640:data<=-16'd7564;
      100641:data<=-16'd7160;
      100642:data<=-16'd7799;
      100643:data<=-16'd6825;
      100644:data<=-16'd2736;
      100645:data<=-16'd1369;
      100646:data<=-16'd3322;
      100647:data<=-16'd3832;
      100648:data<=-16'd2652;
      100649:data<=-16'd2638;
      100650:data<=-16'd3266;
      100651:data<=-16'd2993;
      100652:data<=-16'd3912;
      100653:data<=-16'd5686;
      100654:data<=-16'd5718;
      100655:data<=-16'd5439;
      100656:data<=-16'd5444;
      100657:data<=-16'd5143;
      100658:data<=-16'd5520;
      100659:data<=-16'd6316;
      100660:data<=-16'd7260;
      100661:data<=-16'd7410;
      100662:data<=-16'd7279;
      100663:data<=-16'd8307;
      100664:data<=-16'd5375;
      100665:data<=16'd576;
      100666:data<=16'd632;
      100667:data<=-16'd1372;
      100668:data<=-16'd361;
      100669:data<=-16'd1063;
      100670:data<=-16'd1986;
      100671:data<=-16'd933;
      100672:data<=-16'd1598;
      100673:data<=-16'd3124;
      100674:data<=-16'd3287;
      100675:data<=-16'd3204;
      100676:data<=-16'd3336;
      100677:data<=-16'd2943;
      100678:data<=-16'd2654;
      100679:data<=-16'd4273;
      100680:data<=-16'd6038;
      100681:data<=-16'd5729;
      100682:data<=-16'd5433;
      100683:data<=-16'd5429;
      100684:data<=-16'd5025;
      100685:data<=-16'd5947;
      100686:data<=-16'd7341;
      100687:data<=-16'd7354;
      100688:data<=-16'd6630;
      100689:data<=-16'd6516;
      100690:data<=-16'd6969;
      100691:data<=-16'd6576;
      100692:data<=-16'd6614;
      100693:data<=-16'd8414;
      100694:data<=-16'd9172;
      100695:data<=-16'd8398;
      100696:data<=-16'd8128;
      100697:data<=-16'd7976;
      100698:data<=-16'd7902;
      100699:data<=-16'd8934;
      100700:data<=-16'd10134;
      100701:data<=-16'd9526;
      100702:data<=-16'd8398;
      100703:data<=-16'd8719;
      100704:data<=-16'd8479;
      100705:data<=-16'd8316;
      100706:data<=-16'd9547;
      100707:data<=-16'd8755;
      100708:data<=-16'd8966;
      100709:data<=-16'd14107;
      100710:data<=-16'd18322;
      100711:data<=-16'd20158;
      100712:data<=-16'd22526;
      100713:data<=-16'd23349;
      100714:data<=-16'd22524;
      100715:data<=-16'd21661;
      100716:data<=-16'd20854;
      100717:data<=-16'd20242;
      100718:data<=-16'd19563;
      100719:data<=-16'd19664;
      100720:data<=-16'd19734;
      100721:data<=-16'd18560;
      100722:data<=-16'd18362;
      100723:data<=-16'd18342;
      100724:data<=-16'd17027;
      100725:data<=-16'd16374;
      100726:data<=-16'd16070;
      100727:data<=-16'd15767;
      100728:data<=-16'd15593;
      100729:data<=-16'd14378;
      100730:data<=-16'd13182;
      100731:data<=-16'd12566;
      100732:data<=-16'd12299;
      100733:data<=-16'd12370;
      100734:data<=-16'd11417;
      100735:data<=-16'd10417;
      100736:data<=-16'd9777;
      100737:data<=-16'd8648;
      100738:data<=-16'd8411;
      100739:data<=-16'd7151;
      100740:data<=-16'd4766;
      100741:data<=-16'd4758;
      100742:data<=-16'd4723;
      100743:data<=-16'd3997;
      100744:data<=-16'd4026;
      100745:data<=-16'd2174;
      100746:data<=-16'd393;
      100747:data<=-16'd208;
      100748:data<=16'd585;
      100749:data<=16'd728;
      100750:data<=16'd1248;
      100751:data<=16'd2130;
      100752:data<=16'd1841;
      100753:data<=16'd5685;
      100754:data<=16'd12072;
      100755:data<=16'd13302;
      100756:data<=16'd12179;
      100757:data<=16'd12273;
      100758:data<=16'd12434;
      100759:data<=16'd13359;
      100760:data<=16'd14173;
      100761:data<=16'd13631;
      100762:data<=16'd12975;
      100763:data<=16'd12906;
      100764:data<=16'd12918;
      100765:data<=16'd12951;
      100766:data<=16'd13822;
      100767:data<=16'd14466;
      100768:data<=16'd13952;
      100769:data<=16'd13684;
      100770:data<=16'd12986;
      100771:data<=16'd12396;
      100772:data<=16'd13706;
      100773:data<=16'd14135;
      100774:data<=16'd13565;
      100775:data<=16'd13715;
      100776:data<=16'd12807;
      100777:data<=16'd13697;
      100778:data<=16'd18167;
      100779:data<=16'd20767;
      100780:data<=16'd20395;
      100781:data<=16'd19529;
      100782:data<=16'd18512;
      100783:data<=16'd17920;
      100784:data<=16'd17503;
      100785:data<=16'd17623;
      100786:data<=16'd18656;
      100787:data<=16'd18556;
      100788:data<=16'd17547;
      100789:data<=16'd16844;
      100790:data<=16'd15855;
      100791:data<=16'd15591;
      100792:data<=16'd16512;
      100793:data<=16'd17030;
      100794:data<=16'd16230;
      100795:data<=16'd14844;
      100796:data<=16'd14797;
      100797:data<=16'd14252;
      100798:data<=16'd10147;
      100799:data<=16'd6764;
      100800:data<=16'd7066;
      100801:data<=16'd6910;
      100802:data<=16'd6012;
      100803:data<=16'd6119;
      100804:data<=16'd5598;
      100805:data<=16'd5659;
      100806:data<=16'd7224;
      100807:data<=16'd7423;
      100808:data<=16'd6548;
      100809:data<=16'd6229;
      100810:data<=16'd5683;
      100811:data<=16'd5620;
      100812:data<=16'd6555;
      100813:data<=16'd6956;
      100814:data<=16'd6840;
      100815:data<=16'd6887;
      100816:data<=16'd6546;
      100817:data<=16'd5868;
      100818:data<=16'd5814;
      100819:data<=16'd6716;
      100820:data<=16'd7277;
      100821:data<=16'd6517;
      100822:data<=16'd6024;
      100823:data<=16'd6120;
      100824:data<=16'd5112;
      100825:data<=16'd4924;
      100826:data<=16'd6857;
      100827:data<=16'd7401;
      100828:data<=16'd6664;
      100829:data<=16'd6881;
      100830:data<=16'd6252;
      100831:data<=16'd5739;
      100832:data<=16'd6913;
      100833:data<=16'd7007;
      100834:data<=16'd6763;
      100835:data<=16'd7445;
      100836:data<=16'd7043;
      100837:data<=16'd6566;
      100838:data<=16'd6134;
      100839:data<=16'd5312;
      100840:data<=16'd5636;
      100841:data<=16'd4837;
      100842:data<=16'd5310;
      100843:data<=16'd10941;
      100844:data<=16'd12105;
      100845:data<=16'd5454;
      100846:data<=16'd1767;
      100847:data<=16'd1929;
      100848:data<=16'd1284;
      100849:data<=16'd1227;
      100850:data<=16'd1360;
      100851:data<=16'd481;
      100852:data<=-16'd716;
      100853:data<=-16'd1648;
      100854:data<=-16'd1623;
      100855:data<=-16'd1374;
      100856:data<=-16'd1127;
      100857:data<=-16'd813;
      100858:data<=-16'd2126;
      100859:data<=-16'd3899;
      100860:data<=-16'd4062;
      100861:data<=-16'd4044;
      100862:data<=-16'd4408;
      100863:data<=-16'd4132;
      100864:data<=-16'd3738;
      100865:data<=-16'd4484;
      100866:data<=-16'd5836;
      100867:data<=-16'd6079;
      100868:data<=-16'd5474;
      100869:data<=-16'd4871;
      100870:data<=-16'd4572;
      100871:data<=-16'd5692;
      100872:data<=-16'd7356;
      100873:data<=-16'd7790;
      100874:data<=-16'd7561;
      100875:data<=-16'd7382;
      100876:data<=-16'd7235;
      100877:data<=-16'd6746;
      100878:data<=-16'd6902;
      100879:data<=-16'd8898;
      100880:data<=-16'd9765;
      100881:data<=-16'd8815;
      100882:data<=-16'd8645;
      100883:data<=-16'd7946;
      100884:data<=-16'd7838;
      100885:data<=-16'd9309;
      100886:data<=-16'd8922;
      100887:data<=-16'd10901;
      100888:data<=-16'd16759;
      100889:data<=-16'd17779;
      100890:data<=-16'd15803;
      100891:data<=-16'd16741;
      100892:data<=-16'd17271;
      100893:data<=-16'd17011;
      100894:data<=-16'd17070;
      100895:data<=-16'd16111;
      100896:data<=-16'd15473;
      100897:data<=-16'd15035;
      100898:data<=-16'd15024;
      100899:data<=-16'd16395;
      100900:data<=-16'd16234;
      100901:data<=-16'd15126;
      100902:data<=-16'd15080;
      100903:data<=-16'd13952;
      100904:data<=-16'd13352;
      100905:data<=-16'd14592;
      100906:data<=-16'd14477;
      100907:data<=-16'd13759;
      100908:data<=-16'd13564;
      100909:data<=-16'd12941;
      100910:data<=-16'd13053;
      100911:data<=-16'd11822;
      100912:data<=-16'd8044;
      100913:data<=-16'd6461;
      100914:data<=-16'd6637;
      100915:data<=-16'd5450;
      100916:data<=-16'd4855;
      100917:data<=-16'd4528;
      100918:data<=-16'd4211;
      100919:data<=-16'd5785;
      100920:data<=-16'd6178;
      100921:data<=-16'd4993;
      100922:data<=-16'd5365;
      100923:data<=-16'd5083;
      100924:data<=-16'd4423;
      100925:data<=-16'd5617;
      100926:data<=-16'd6008;
      100927:data<=-16'd5612;
      100928:data<=-16'd5344;
      100929:data<=-16'd4764;
      100930:data<=-16'd5607;
      100931:data<=-16'd4504;
      100932:data<=16'd414;
      100933:data<=16'd2655;
      100934:data<=16'd2018;
      100935:data<=16'd2153;
      100936:data<=16'd2000;
      100937:data<=16'd2303;
      100938:data<=16'd2551;
      100939:data<=16'd1172;
      100940:data<=16'd785;
      100941:data<=16'd1434;
      100942:data<=16'd1468;
      100943:data<=16'd1419;
      100944:data<=16'd955;
      100945:data<=16'd990;
      100946:data<=16'd1898;
      100947:data<=16'd1871;
      100948:data<=16'd1771;
      100949:data<=16'd2093;
      100950:data<=16'd1767;
      100951:data<=16'd2502;
      100952:data<=16'd4490;
      100953:data<=16'd4893;
      100954:data<=16'd4372;
      100955:data<=16'd5090;
      100956:data<=16'd5277;
      100957:data<=16'd4673;
      100958:data<=16'd5883;
      100959:data<=16'd6810;
      100960:data<=16'd5908;
      100961:data<=16'd6231;
      100962:data<=16'd6755;
      100963:data<=16'd6061;
      100964:data<=16'd6470;
      100965:data<=16'd7611;
      100966:data<=16'd8335;
      100967:data<=16'd8025;
      100968:data<=16'd6769;
      100969:data<=16'd6764;
      100970:data<=16'd6742;
      100971:data<=16'd6628;
      100972:data<=16'd8461;
      100973:data<=16'd8376;
      100974:data<=16'd7586;
      100975:data<=16'd9166;
      100976:data<=16'd6299;
      100977:data<=16'd470;
      100978:data<=-16'd1571;
      100979:data<=-16'd3711;
      100980:data<=-16'd5703;
      100981:data<=-16'd4736;
      100982:data<=-16'd4664;
      100983:data<=-16'd4890;
      100984:data<=-16'd3688;
      100985:data<=-16'd2573;
      100986:data<=-16'd1228;
      100987:data<=-16'd796;
      100988:data<=-16'd1280;
      100989:data<=-16'd860;
      100990:data<=-16'd688;
      100991:data<=-16'd349;
      100992:data<=16'd998;
      100993:data<=16'd1415;
      100994:data<=16'd1002;
      100995:data<=16'd854;
      100996:data<=16'd805;
      100997:data<=16'd1518;
      100998:data<=16'd3363;
      100999:data<=16'd4590;
      101000:data<=16'd4112;
      101001:data<=16'd3839;
      101002:data<=16'd4117;
      101003:data<=16'd3733;
      101004:data<=16'd4355;
      101005:data<=16'd5805;
      101006:data<=16'd5947;
      101007:data<=16'd5548;
      101008:data<=16'd5415;
      101009:data<=16'd5905;
      101010:data<=16'd6434;
      101011:data<=16'd6291;
      101012:data<=16'd7464;
      101013:data<=16'd8291;
      101014:data<=16'd7113;
      101015:data<=16'd7154;
      101016:data<=16'd6986;
      101017:data<=16'd6699;
      101018:data<=16'd8887;
      101019:data<=16'd8704;
      101020:data<=16'd8363;
      101021:data<=16'd13373;
      101022:data<=16'd16352;
      101023:data<=16'd15239;
      101024:data<=16'd15505;
      101025:data<=16'd15887;
      101026:data<=16'd15693;
      101027:data<=16'd15277;
      101028:data<=16'd14183;
      101029:data<=16'd13888;
      101030:data<=16'd13217;
      101031:data<=16'd12640;
      101032:data<=16'd13864;
      101033:data<=16'd14005;
      101034:data<=16'd13160;
      101035:data<=16'd13139;
      101036:data<=16'd12590;
      101037:data<=16'd12116;
      101038:data<=16'd12451;
      101039:data<=16'd12687;
      101040:data<=16'd12322;
      101041:data<=16'd11499;
      101042:data<=16'd11392;
      101043:data<=16'd10900;
      101044:data<=16'd9734;
      101045:data<=16'd11861;
      101046:data<=16'd16063;
      101047:data<=16'd17024;
      101048:data<=16'd15402;
      101049:data<=16'd14468;
      101050:data<=16'd14022;
      101051:data<=16'd12807;
      101052:data<=16'd12054;
      101053:data<=16'd11902;
      101054:data<=16'd10543;
      101055:data<=16'd9699;
      101056:data<=16'd9700;
      101057:data<=16'd8067;
      101058:data<=16'd6536;
      101059:data<=16'd5735;
      101060:data<=16'd4769;
      101061:data<=16'd4629;
      101062:data<=16'd3407;
      101063:data<=16'd2488;
      101064:data<=16'd3207;
      101065:data<=-16'd1169;
      101066:data<=-16'd8149;
      101067:data<=-16'd9392;
      101068:data<=-16'd8845;
      101069:data<=-16'd9323;
      101070:data<=-16'd8789;
      101071:data<=-16'd9800;
      101072:data<=-16'd11277;
      101073:data<=-16'd10534;
      101074:data<=-16'd9985;
      101075:data<=-16'd10064;
      101076:data<=-16'd9711;
      101077:data<=-16'd10176;
      101078:data<=-16'd11524;
      101079:data<=-16'd12101;
      101080:data<=-16'd11665;
      101081:data<=-16'd11594;
      101082:data<=-16'd11479;
      101083:data<=-16'd10542;
      101084:data<=-16'd10936;
      101085:data<=-16'd12536;
      101086:data<=-16'd12513;
      101087:data<=-16'd11741;
      101088:data<=-16'd11679;
      101089:data<=-16'd11244;
      101090:data<=-16'd11001;
      101091:data<=-16'd11994;
      101092:data<=-16'd12689;
      101093:data<=-16'd12172;
      101094:data<=-16'd11655;
      101095:data<=-16'd11359;
      101096:data<=-16'd10784;
      101097:data<=-16'd10900;
      101098:data<=-16'd11737;
      101099:data<=-16'd11705;
      101100:data<=-16'd11209;
      101101:data<=-16'd11303;
      101102:data<=-16'd10968;
      101103:data<=-16'd10194;
      101104:data<=-16'd10651;
      101105:data<=-16'd12007;
      101106:data<=-16'd12184;
      101107:data<=-16'd11080;
      101108:data<=-16'd11039;
      101109:data<=-16'd11288;
      101110:data<=-16'd7535;
      101111:data<=-16'd2695;
      101112:data<=-16'd4070;
      101113:data<=-16'd8419;
      101114:data<=-16'd9464;
      101115:data<=-16'd9344;
      101116:data<=-16'd9335;
      101117:data<=-16'd8596;
      101118:data<=-16'd9342;
      101119:data<=-16'd10571;
      101120:data<=-16'd9966;
      101121:data<=-16'd9323;
      101122:data<=-16'd9085;
      101123:data<=-16'd8291;
      101124:data<=-16'd8273;
      101125:data<=-16'd9279;
      101126:data<=-16'd9738;
      101127:data<=-16'd9462;
      101128:data<=-16'd9083;
      101129:data<=-16'd8417;
      101130:data<=-16'd7976;
      101131:data<=-16'd8783;
      101132:data<=-16'd9511;
      101133:data<=-16'd8881;
      101134:data<=-16'd8493;
      101135:data<=-16'd8707;
      101136:data<=-16'd8087;
      101137:data<=-16'd7841;
      101138:data<=-16'd9110;
      101139:data<=-16'd9491;
      101140:data<=-16'd8466;
      101141:data<=-16'd8373;
      101142:data<=-16'd8405;
      101143:data<=-16'd7571;
      101144:data<=-16'd7917;
      101145:data<=-16'd9051;
      101146:data<=-16'd8974;
      101147:data<=-16'd8204;
      101148:data<=-16'd7802;
      101149:data<=-16'd7680;
      101150:data<=-16'd7374;
      101151:data<=-16'd7920;
      101152:data<=-16'd8866;
      101153:data<=-16'd7697;
      101154:data<=-16'd8442;
      101155:data<=-16'd13843;
      101156:data<=-16'd16283;
      101157:data<=-16'd14501;
      101158:data<=-16'd14067;
      101159:data<=-16'd13579;
      101160:data<=-16'd12330;
      101161:data<=-16'd12067;
      101162:data<=-16'd11709;
      101163:data<=-16'd11174;
      101164:data<=-16'd9670;
      101165:data<=-16'd7488;
      101166:data<=-16'd7086;
      101167:data<=-16'd6561;
      101168:data<=-16'd5204;
      101169:data<=-16'd5491;
      101170:data<=-16'd5459;
      101171:data<=-16'd3524;
      101172:data<=-16'd2108;
      101173:data<=-16'd1959;
      101174:data<=-16'd1889;
      101175:data<=-16'd1818;
      101176:data<=-16'd1619;
      101177:data<=-16'd517;
      101178:data<=16'd591;
      101179:data<=16'd2346;
      101180:data<=16'd6304;
      101181:data<=16'd8355;
      101182:data<=16'd7394;
      101183:data<=16'd8079;
      101184:data<=16'd9397;
      101185:data<=16'd9791;
      101186:data<=16'd10050;
      101187:data<=16'd9133;
      101188:data<=16'd8983;
      101189:data<=16'd9638;
      101190:data<=16'd9582;
      101191:data<=16'd10827;
      101192:data<=16'd11068;
      101193:data<=16'd10078;
      101194:data<=16'd11013;
      101195:data<=16'd10671;
      101196:data<=16'd10175;
      101197:data<=16'd11402;
      101198:data<=16'd10766;
      101199:data<=16'd13018;
      101200:data<=16'd19035;
      101201:data<=16'd20334;
      101202:data<=16'd18515;
      101203:data<=16'd18240;
      101204:data<=16'd18813;
      101205:data<=16'd19506;
      101206:data<=16'd18762;
      101207:data<=16'd17602;
      101208:data<=16'd17350;
      101209:data<=16'd16712;
      101210:data<=16'd16845;
      101211:data<=16'd17623;
      101212:data<=16'd17499;
      101213:data<=16'd17176;
      101214:data<=16'd16759;
      101215:data<=16'd16236;
      101216:data<=16'd15209;
      101217:data<=16'd14481;
      101218:data<=16'd15726;
      101219:data<=16'd16111;
      101220:data<=16'd14968;
      101221:data<=16'd14703;
      101222:data<=16'd13952;
      101223:data<=16'd13345;
      101224:data<=16'd14201;
      101225:data<=16'd14647;
      101226:data<=16'd14186;
      101227:data<=16'd12897;
      101228:data<=16'd12222;
      101229:data<=16'd12704;
      101230:data<=16'd12326;
      101231:data<=16'd12730;
      101232:data<=16'd13439;
      101233:data<=16'd11897;
      101234:data<=16'd10748;
      101235:data<=16'd10132;
      101236:data<=16'd9415;
      101237:data<=16'd10199;
      101238:data<=16'd10699;
      101239:data<=16'd10930;
      101240:data<=16'd10437;
      101241:data<=16'd8675;
      101242:data<=16'd9391;
      101243:data<=16'd8392;
      101244:data<=16'd3272;
      101245:data<=16'd1739;
      101246:data<=16'd359;
      101247:data<=-16'd4686;
      101248:data<=-16'd5864;
      101249:data<=-16'd4761;
      101250:data<=-16'd5391;
      101251:data<=-16'd4449;
      101252:data<=-16'd3457;
      101253:data<=-16'd4088;
      101254:data<=-16'd3833;
      101255:data<=-16'd3303;
      101256:data<=-16'd3529;
      101257:data<=-16'd2839;
      101258:data<=-16'd1152;
      101259:data<=-16'd784;
      101260:data<=-16'd1536;
      101261:data<=-16'd1391;
      101262:data<=-16'd910;
      101263:data<=-16'd919;
      101264:data<=-16'd1348;
      101265:data<=-16'd1804;
      101266:data<=-16'd1554;
      101267:data<=-16'd1665;
      101268:data<=-16'd1682;
      101269:data<=-16'd857;
      101270:data<=-16'd2073;
      101271:data<=-16'd4106;
      101272:data<=-16'd4029;
      101273:data<=-16'd4041;
      101274:data<=-16'd4431;
      101275:data<=-16'd4237;
      101276:data<=-16'd4253;
      101277:data<=-16'd4422;
      101278:data<=-16'd5410;
      101279:data<=-16'd5862;
      101280:data<=-16'd4908;
      101281:data<=-16'd5269;
      101282:data<=-16'd5277;
      101283:data<=-16'd4572;
      101284:data<=-16'd6357;
      101285:data<=-16'd6811;
      101286:data<=-16'd5592;
      101287:data<=-16'd7012;
      101288:data<=-16'd5177;
      101289:data<=16'd1375;
      101290:data<=16'd2887;
      101291:data<=-16'd44;
      101292:data<=-16'd191;
      101293:data<=16'd647;
      101294:data<=16'd42;
      101295:data<=16'd42;
      101296:data<=-16'd30;
      101297:data<=-16'd1428;
      101298:data<=-16'd2472;
      101299:data<=-16'd2455;
      101300:data<=-16'd2105;
      101301:data<=-16'd1760;
      101302:data<=-16'd1953;
      101303:data<=-16'd3001;
      101304:data<=-16'd4179;
      101305:data<=-16'd4411;
      101306:data<=-16'd4194;
      101307:data<=-16'd4541;
      101308:data<=-16'd4563;
      101309:data<=-16'd4141;
      101310:data<=-16'd4317;
      101311:data<=-16'd5109;
      101312:data<=-16'd6049;
      101313:data<=-16'd4467;
      101314:data<=-16'd76;
      101315:data<=16'd1715;
      101316:data<=16'd723;
      101317:data<=16'd191;
      101318:data<=-16'd1119;
      101319:data<=-16'd1759;
      101320:data<=-16'd751;
      101321:data<=-16'd1196;
      101322:data<=-16'd1709;
      101323:data<=-16'd1871;
      101324:data<=-16'd3802;
      101325:data<=-16'd4455;
      101326:data<=-16'd3727;
      101327:data<=-16'd4393;
      101328:data<=-16'd3891;
      101329:data<=-16'd2816;
      101330:data<=-16'd4410;
      101331:data<=-16'd5424;
      101332:data<=-16'd5477;
      101333:data<=-16'd9301;
      101334:data<=-16'd13532;
      101335:data<=-16'd13085;
      101336:data<=-16'd12213;
      101337:data<=-16'd13552;
      101338:data<=-16'd13893;
      101339:data<=-16'd13132;
      101340:data<=-16'd12609;
      101341:data<=-16'd12161;
      101342:data<=-16'd11688;
      101343:data<=-16'd11341;
      101344:data<=-16'd12201;
      101345:data<=-16'd12904;
      101346:data<=-16'd11602;
      101347:data<=-16'd11033;
      101348:data<=-16'd11056;
      101349:data<=-16'd9680;
      101350:data<=-16'd9925;
      101351:data<=-16'd11254;
      101352:data<=-16'd10555;
      101353:data<=-16'd9727;
      101354:data<=-16'd9549;
      101355:data<=-16'd9323;
      101356:data<=-16'd9591;
      101357:data<=-16'd9502;
      101358:data<=-16'd9411;
      101359:data<=-16'd9843;
      101360:data<=-16'd9415;
      101361:data<=-16'd8743;
      101362:data<=-16'd8390;
      101363:data<=-16'd7774;
      101364:data<=-16'd8037;
      101365:data<=-16'd8624;
      101366:data<=-16'd7911;
      101367:data<=-16'd7301;
      101368:data<=-16'd7178;
      101369:data<=-16'd6394;
      101370:data<=-16'd5812;
      101371:data<=-16'd5427;
      101372:data<=-16'd4690;
      101373:data<=-16'd4306;
      101374:data<=-16'd3623;
      101375:data<=-16'd3462;
      101376:data<=-16'd4168;
      101377:data<=-16'd701;
      101378:data<=16'd6287;
      101379:data<=16'd8895;
      101380:data<=16'd6282;
      101381:data<=16'd2875;
      101382:data<=16'd1409;
      101383:data<=16'd2502;
      101384:data<=16'd3629;
      101385:data<=16'd3717;
      101386:data<=16'd3789;
      101387:data<=16'd3647;
      101388:data<=16'd3862;
      101389:data<=16'd4196;
      101390:data<=16'd4614;
      101391:data<=16'd6208;
      101392:data<=16'd6819;
      101393:data<=16'd6166;
      101394:data<=16'd6115;
      101395:data<=16'd5533;
      101396:data<=16'd5749;
      101397:data<=16'd7526;
      101398:data<=16'd7900;
      101399:data<=16'd7614;
      101400:data<=16'd7908;
      101401:data<=16'd7903;
      101402:data<=16'd7853;
      101403:data<=16'd7982;
      101404:data<=16'd8887;
      101405:data<=16'd9357;
      101406:data<=16'd8405;
      101407:data<=16'd8554;
      101408:data<=16'd8762;
      101409:data<=16'd8058;
      101410:data<=16'd9012;
      101411:data<=16'd9612;
      101412:data<=16'd8837;
      101413:data<=16'd8769;
      101414:data<=16'd8357;
      101415:data<=16'd7949;
      101416:data<=16'd8445;
      101417:data<=16'd9294;
      101418:data<=16'd9887;
      101419:data<=16'd8425;
      101420:data<=16'd7899;
      101421:data<=16'd9280;
      101422:data<=16'd5460;
      101423:data<=-16'd196;
      101424:data<=16'd564;
      101425:data<=16'd2575;
      101426:data<=16'd1680;
      101427:data<=16'd1295;
      101428:data<=16'd1403;
      101429:data<=16'd1084;
      101430:data<=16'd1777;
      101431:data<=16'd3301;
      101432:data<=16'd3700;
      101433:data<=16'd2875;
      101434:data<=16'd2400;
      101435:data<=16'd2529;
      101436:data<=16'd3290;
      101437:data<=16'd4273;
      101438:data<=16'd4531;
      101439:data<=16'd4661;
      101440:data<=16'd4358;
      101441:data<=16'd3638;
      101442:data<=16'd3736;
      101443:data<=16'd4041;
      101444:data<=16'd5016;
      101445:data<=16'd5671;
      101446:data<=16'd4172;
      101447:data<=16'd5289;
      101448:data<=16'd9459;
      101449:data<=16'd10933;
      101450:data<=16'd11277;
      101451:data<=16'd11843;
      101452:data<=16'd10701;
      101453:data<=16'd10091;
      101454:data<=16'd10288;
      101455:data<=16'd9973;
      101456:data<=16'd10240;
      101457:data<=16'd11086;
      101458:data<=16'd11195;
      101459:data<=16'd9621;
      101460:data<=16'd9047;
      101461:data<=16'd10319;
      101462:data<=16'd9133;
      101463:data<=16'd8775;
      101464:data<=16'd11239;
      101465:data<=16'd9668;
      101466:data<=16'd9238;
      101467:data<=16'd15352;
      101468:data<=16'd18016;
      101469:data<=16'd16172;
      101470:data<=16'd16284;
      101471:data<=16'd16324;
      101472:data<=16'd15734;
      101473:data<=16'd15653;
      101474:data<=16'd14880;
      101475:data<=16'd14163;
      101476:data<=16'd13377;
      101477:data<=16'd12333;
      101478:data<=16'd11973;
      101479:data<=16'd11462;
      101480:data<=16'd10581;
      101481:data<=16'd9871;
      101482:data<=16'd9124;
      101483:data<=16'd7871;
      101484:data<=16'd5903;
      101485:data<=16'd4722;
      101486:data<=16'd4498;
      101487:data<=16'd4140;
      101488:data<=16'd4610;
      101489:data<=16'd4425;
      101490:data<=16'd1988;
      101491:data<=16'd461;
      101492:data<=16'd623;
      101493:data<=16'd347;
      101494:data<=-16'd273;
      101495:data<=-16'd644;
      101496:data<=-16'd984;
      101497:data<=-16'd1908;
      101498:data<=-16'd2605;
      101499:data<=-16'd2461;
      101500:data<=-16'd3338;
      101501:data<=-16'd4008;
      101502:data<=-16'd3548;
      101503:data<=-16'd5037;
      101504:data<=-16'd6434;
      101505:data<=-16'd6100;
      101506:data<=-16'd6742;
      101507:data<=-16'd6378;
      101508:data<=-16'd5956;
      101509:data<=-16'd7592;
      101510:data<=-16'd7339;
      101511:data<=-16'd9409;
      101512:data<=-16'd15850;
      101513:data<=-16'd16851;
      101514:data<=-16'd16137;
      101515:data<=-16'd20956;
      101516:data<=-16'd23041;
      101517:data<=-16'd21646;
      101518:data<=-16'd22527;
      101519:data<=-16'd22230;
      101520:data<=-16'd20372;
      101521:data<=-16'd19664;
      101522:data<=-16'd19299;
      101523:data<=-16'd20178;
      101524:data<=-16'd21147;
      101525:data<=-16'd19851;
      101526:data<=-16'd18494;
      101527:data<=-16'd17987;
      101528:data<=-16'd17353;
      101529:data<=-16'd17708;
      101530:data<=-16'd18662;
      101531:data<=-16'd18265;
      101532:data<=-16'd17214;
      101533:data<=-16'd17136;
      101534:data<=-16'd16985;
      101535:data<=-16'd15749;
      101536:data<=-16'd15233;
      101537:data<=-16'd16084;
      101538:data<=-16'd16301;
      101539:data<=-16'd15280;
      101540:data<=-16'd14311;
      101541:data<=-16'd13890;
      101542:data<=-16'd13788;
      101543:data<=-16'd14293;
      101544:data<=-16'd14647;
      101545:data<=-16'd13538;
      101546:data<=-16'd12205;
      101547:data<=-16'd11723;
      101548:data<=-16'd11479;
      101549:data<=-16'd11913;
      101550:data<=-16'd12430;
      101551:data<=-16'd12054;
      101552:data<=-16'd11546;
      101553:data<=-16'd10860;
      101554:data<=-16'd10442;
      101555:data<=-16'd9289;
      101556:data<=-16'd4896;
      101557:data<=-16'd1548;
      101558:data<=-16'd2206;
      101559:data<=-16'd1847;
      101560:data<=-16'd561;
      101561:data<=-16'd1068;
      101562:data<=-16'd1639;
      101563:data<=-16'd2537;
      101564:data<=-16'd3268;
      101565:data<=-16'd2760;
      101566:data<=-16'd3122;
      101567:data<=-16'd3066;
      101568:data<=-16'd1710;
      101569:data<=-16'd2012;
      101570:data<=-16'd3259;
      101571:data<=-16'd3911;
      101572:data<=-16'd4094;
      101573:data<=-16'd3548;
      101574:data<=-16'd3324;
      101575:data<=-16'd2907;
      101576:data<=-16'd2505;
      101577:data<=-16'd4085;
      101578:data<=-16'd4360;
      101579:data<=-16'd2908;
      101580:data<=-16'd3930;
      101581:data<=-16'd3112;
      101582:data<=16'd1842;
      101583:data<=16'd4055;
      101584:data<=16'd3541;
      101585:data<=16'd3905;
      101586:data<=16'd3513;
      101587:data<=16'd3011;
      101588:data<=16'd3475;
      101589:data<=16'd3703;
      101590:data<=16'd4616;
      101591:data<=16'd5327;
      101592:data<=16'd4643;
      101593:data<=16'd4878;
      101594:data<=16'd5169;
      101595:data<=16'd4619;
      101596:data<=16'd5749;
      101597:data<=16'd6416;
      101598:data<=16'd5830;
      101599:data<=16'd7009;
      101600:data<=16'd4910;
      101601:data<=-16'd1959;
      101602:data<=-16'd3701;
      101603:data<=-16'd411;
      101604:data<=-16'd164;
      101605:data<=-16'd1172;
      101606:data<=-16'd490;
      101607:data<=-16'd385;
      101608:data<=-16'd508;
      101609:data<=16'd640;
      101610:data<=16'd1997;
      101611:data<=16'd2306;
      101612:data<=16'd2088;
      101613:data<=16'd2191;
      101614:data<=16'd1926;
      101615:data<=16'd1803;
      101616:data<=16'd3338;
      101617:data<=16'd4654;
      101618:data<=16'd4173;
      101619:data<=16'd3988;
      101620:data<=16'd4372;
      101621:data<=16'd3842;
      101622:data<=16'd3982;
      101623:data<=16'd5479;
      101624:data<=16'd5764;
      101625:data<=16'd5245;
      101626:data<=16'd5623;
      101627:data<=16'd5275;
      101628:data<=16'd4773;
      101629:data<=16'd5944;
      101630:data<=16'd6909;
      101631:data<=16'd7265;
      101632:data<=16'd7711;
      101633:data<=16'd6896;
      101634:data<=16'd5900;
      101635:data<=16'd6578;
      101636:data<=16'd8337;
      101637:data<=16'd9521;
      101638:data<=16'd8845;
      101639:data<=16'd8128;
      101640:data<=16'd8404;
      101641:data<=16'd8046;
      101642:data<=16'd8514;
      101643:data<=16'd9495;
      101644:data<=16'd9101;
      101645:data<=16'd11455;
      101646:data<=16'd16713;
      101647:data<=16'd18028;
      101648:data<=16'd14257;
      101649:data<=16'd10540;
      101650:data<=16'd10261;
      101651:data<=16'd10813;
      101652:data<=16'd9605;
      101653:data<=16'd9219;
      101654:data<=16'd9356;
      101655:data<=16'd8728;
      101656:data<=16'd9624;
      101657:data<=16'd10207;
      101658:data<=16'd9188;
      101659:data<=16'd9092;
      101660:data<=16'd8883;
      101661:data<=16'd8208;
      101662:data<=16'd8451;
      101663:data<=16'd9145;
      101664:data<=16'd9840;
      101665:data<=16'd9210;
      101666:data<=16'd8416;
      101667:data<=16'd8971;
      101668:data<=16'd8062;
      101669:data<=16'd7571;
      101670:data<=16'd9652;
      101671:data<=16'd9781;
      101672:data<=16'd8423;
      101673:data<=16'd8381;
      101674:data<=16'd8156;
      101675:data<=16'd8140;
      101676:data<=16'd8607;
      101677:data<=16'd8413;
      101678:data<=16'd8085;
      101679:data<=16'd7979;
      101680:data<=16'd7639;
      101681:data<=16'd6781;
      101682:data<=16'd6805;
      101683:data<=16'd7598;
      101684:data<=16'd6948;
      101685:data<=16'd6534;
      101686:data<=16'd6419;
      101687:data<=16'd5371;
      101688:data<=16'd6140;
      101689:data<=16'd4567;
      101690:data<=-16'd1788;
      101691:data<=-16'd4322;
      101692:data<=-16'd3474;
      101693:data<=-16'd4131;
      101694:data<=-16'd3582;
      101695:data<=-16'd3492;
      101696:data<=-16'd5389;
      101697:data<=-16'd6164;
      101698:data<=-16'd6273;
      101699:data<=-16'd6338;
      101700:data<=-16'd6123;
      101701:data<=-16'd5927;
      101702:data<=-16'd6166;
      101703:data<=-16'd7600;
      101704:data<=-16'd7755;
      101705:data<=-16'd6849;
      101706:data<=-16'd7661;
      101707:data<=-16'd7394;
      101708:data<=-16'd6507;
      101709:data<=-16'd7486;
      101710:data<=-16'd7953;
      101711:data<=-16'd8449;
      101712:data<=-16'd8769;
      101713:data<=-16'd7829;
      101714:data<=-16'd7793;
      101715:data<=-16'd6131;
      101716:data<=-16'd3168;
      101717:data<=-16'd3195;
      101718:data<=-16'd3344;
      101719:data<=-16'd3033;
      101720:data<=-16'd3479;
      101721:data<=-16'd2473;
      101722:data<=-16'd2773;
      101723:data<=-16'd4508;
      101724:data<=-16'd4220;
      101725:data<=-16'd3888;
      101726:data<=-16'd3855;
      101727:data<=-16'd3269;
      101728:data<=-16'd3336;
      101729:data<=-16'd4062;
      101730:data<=-16'd5442;
      101731:data<=-16'd5266;
      101732:data<=-16'd4382;
      101733:data<=-16'd5523;
      101734:data<=-16'd2541;
      101735:data<=16'd3459;
      101736:data<=16'd2996;
      101737:data<=16'd813;
      101738:data<=16'd2000;
      101739:data<=16'd1968;
      101740:data<=16'd1589;
      101741:data<=16'd1806;
      101742:data<=16'd359;
      101743:data<=-16'd1014;
      101744:data<=-16'd1327;
      101745:data<=-16'd1394;
      101746:data<=-16'd1055;
      101747:data<=-16'd450;
      101748:data<=-16'd644;
      101749:data<=-16'd2406;
      101750:data<=-16'd3277;
      101751:data<=-16'd2055;
      101752:data<=-16'd1757;
      101753:data<=-16'd2346;
      101754:data<=-16'd2362;
      101755:data<=-16'd2889;
      101756:data<=-16'd3556;
      101757:data<=-16'd3612;
      101758:data<=-16'd3626;
      101759:data<=-16'd4111;
      101760:data<=-16'd4557;
      101761:data<=-16'd3788;
      101762:data<=-16'd3604;
      101763:data<=-16'd5083;
      101764:data<=-16'd5365;
      101765:data<=-16'd4739;
      101766:data<=-16'd4614;
      101767:data<=-16'd3999;
      101768:data<=-16'd4162;
      101769:data<=-16'd5557;
      101770:data<=-16'd6347;
      101771:data<=-16'd6200;
      101772:data<=-16'd5671;
      101773:data<=-16'd5752;
      101774:data<=-16'd5841;
      101775:data<=-16'd5705;
      101776:data<=-16'd7130;
      101777:data<=-16'd7291;
      101778:data<=-16'd6622;
      101779:data<=-16'd11251;
      101780:data<=-16'd15074;
      101781:data<=-16'd12678;
      101782:data<=-16'd14530;
      101783:data<=-16'd21017;
      101784:data<=-16'd21598;
      101785:data<=-16'd19077;
      101786:data<=-16'd18751;
      101787:data<=-16'd17887;
      101788:data<=-16'd17236;
      101789:data<=-16'd18157;
      101790:data<=-16'd17729;
      101791:data<=-16'd16762;
      101792:data<=-16'd17220;
      101793:data<=-16'd16512;
      101794:data<=-16'd14727;
      101795:data<=-16'd14427;
      101796:data<=-16'd13856;
      101797:data<=-16'd12228;
      101798:data<=-16'd11295;
      101799:data<=-16'd10383;
      101800:data<=-16'd9812;
      101801:data<=-16'd10064;
      101802:data<=-16'd8751;
      101803:data<=-16'd6490;
      101804:data<=-16'd5501;
      101805:data<=-16'd4810;
      101806:data<=-16'd4234;
      101807:data<=-16'd4432;
      101808:data<=-16'd3665;
      101809:data<=-16'd1177;
      101810:data<=16'd390;
      101811:data<=-16'd126;
      101812:data<=-16'd241;
      101813:data<=16'd405;
      101814:data<=16'd567;
      101815:data<=16'd1689;
      101816:data<=16'd3469;
      101817:data<=16'd3943;
      101818:data<=16'd3636;
      101819:data<=16'd3418;
      101820:data<=16'd3971;
      101821:data<=16'd4272;
      101822:data<=16'd3858;
      101823:data<=16'd7486;
      101824:data<=16'd13744;
      101825:data<=16'd15203;
      101826:data<=16'd14202;
      101827:data<=16'd14472;
      101828:data<=16'd14408;
      101829:data<=16'd15265;
      101830:data<=16'd15963;
      101831:data<=16'd14718;
      101832:data<=16'd14434;
      101833:data<=16'd14433;
      101834:data<=16'd13838;
      101835:data<=16'd14897;
      101836:data<=16'd15790;
      101837:data<=16'd15235;
      101838:data<=16'd14784;
      101839:data<=16'd14111;
      101840:data<=16'd13405;
      101841:data<=16'd13388;
      101842:data<=16'd13878;
      101843:data<=16'd14546;
      101844:data<=16'd14296;
      101845:data<=16'd13544;
      101846:data<=16'd13456;
      101847:data<=16'd12706;
      101848:data<=16'd12016;
      101849:data<=16'd15238;
      101850:data<=16'd20110;
      101851:data<=16'd20333;
      101852:data<=16'd18468;
      101853:data<=16'd18726;
      101854:data<=16'd17525;
      101855:data<=16'd16295;
      101856:data<=16'd18371;
      101857:data<=16'd18539;
      101858:data<=16'd16712;
      101859:data<=16'd16365;
      101860:data<=16'd14957;
      101861:data<=16'd13910;
      101862:data<=16'd15001;
      101863:data<=16'd15177;
      101864:data<=16'd14216;
      101865:data<=16'd12845;
      101866:data<=16'd12625;
      101867:data<=16'd13047;
      101868:data<=16'd9185;
      101869:data<=16'd4708;
      101870:data<=16'd4689;
      101871:data<=16'd4467;
      101872:data<=16'd3453;
      101873:data<=16'd3413;
      101874:data<=16'd2319;
      101875:data<=16'd2337;
      101876:data<=16'd4190;
      101877:data<=16'd4399;
      101878:data<=16'd3300;
      101879:data<=16'd2784;
      101880:data<=16'd2567;
      101881:data<=16'd2340;
      101882:data<=16'd3391;
      101883:data<=16'd4761;
      101884:data<=16'd3739;
      101885:data<=16'd3036;
      101886:data<=16'd3826;
      101887:data<=16'd2925;
      101888:data<=16'd2889;
      101889:data<=16'd4473;
      101890:data<=16'd3982;
      101891:data<=16'd3262;
      101892:data<=16'd3224;
      101893:data<=16'd2341;
      101894:data<=16'd2341;
      101895:data<=16'd3441;
      101896:data<=16'd4394;
      101897:data<=16'd4545;
      101898:data<=16'd3777;
      101899:data<=16'd3536;
      101900:data<=16'd3755;
      101901:data<=16'd3460;
      101902:data<=16'd2648;
      101903:data<=16'd2061;
      101904:data<=16'd2487;
      101905:data<=16'd2162;
      101906:data<=16'd1797;
      101907:data<=16'd2661;
      101908:data<=16'd1139;
      101909:data<=-16'd485;
      101910:data<=-16'd350;
      101911:data<=-16'd2667;
      101912:data<=-16'd1512;
      101913:data<=16'd4816;
      101914:data<=16'd6792;
      101915:data<=16'd5504;
      101916:data<=16'd2458;
      101917:data<=-16'd3104;
      101918:data<=-16'd4131;
      101919:data<=-16'd2631;
      101920:data<=-16'd3378;
      101921:data<=-16'd3498;
      101922:data<=-16'd4679;
      101923:data<=-16'd5955;
      101924:data<=-16'd4857;
      101925:data<=-16'd5021;
      101926:data<=-16'd5242;
      101927:data<=-16'd4673;
      101928:data<=-16'd5548;
      101929:data<=-16'd6132;
      101930:data<=-16'd6822;
      101931:data<=-16'd7238;
      101932:data<=-16'd6293;
      101933:data<=-16'd6449;
      101934:data<=-16'd6387;
      101935:data<=-16'd6432;
      101936:data<=-16'd8325;
      101937:data<=-16'd8284;
      101938:data<=-16'd7491;
      101939:data<=-16'd8043;
      101940:data<=-16'd7409;
      101941:data<=-16'd7548;
      101942:data<=-16'd8868;
      101943:data<=-16'd9138;
      101944:data<=-16'd9182;
      101945:data<=-16'd8760;
      101946:data<=-16'd8451;
      101947:data<=-16'd8434;
      101948:data<=-16'd8498;
      101949:data<=-16'd10378;
      101950:data<=-16'd10847;
      101951:data<=-16'd9547;
      101952:data<=-16'd10187;
      101953:data<=-16'd9368;
      101954:data<=-16'd8728;
      101955:data<=-16'd10928;
      101956:data<=-16'd10351;
      101957:data<=-16'd11646;
      101958:data<=-16'd17697;
      101959:data<=-16'd18545;
      101960:data<=-16'd16292;
      101961:data<=-16'd17428;
      101962:data<=-16'd18330;
      101963:data<=-16'd17979;
      101964:data<=-16'd17330;
      101965:data<=-16'd16594;
      101966:data<=-16'd16452;
      101967:data<=-16'd15509;
      101968:data<=-16'd14960;
      101969:data<=-16'd15694;
      101970:data<=-16'd15825;
      101971:data<=-16'd15673;
      101972:data<=-16'd14853;
      101973:data<=-16'd13834;
      101974:data<=-16'd14093;
      101975:data<=-16'd14028;
      101976:data<=-16'd14037;
      101977:data<=-16'd13978;
      101978:data<=-16'd12689;
      101979:data<=-16'd12750;
      101980:data<=-16'd12481;
      101981:data<=-16'd11301;
      101982:data<=-16'd12739;
      101983:data<=-16'd10974;
      101984:data<=-16'd5189;
      101985:data<=-16'd4423;
      101986:data<=-16'd5101;
      101987:data<=-16'd2934;
      101988:data<=-16'd3630;
      101989:data<=-16'd5559;
      101990:data<=-16'd5069;
      101991:data<=-16'd4619;
      101992:data<=-16'd4308;
      101993:data<=-16'd3657;
      101994:data<=-16'd4046;
      101995:data<=-16'd5177;
      101996:data<=-16'd5410;
      101997:data<=-16'd4266;
      101998:data<=-16'd3595;
      101999:data<=-16'd3970;
      102000:data<=-16'd4250;
      102001:data<=-16'd3797;
      102002:data<=-16'd867;
      102003:data<=16'd2886;
      102004:data<=16'd3475;
      102005:data<=16'd3119;
      102006:data<=16'd3674;
      102007:data<=16'd3233;
      102008:data<=16'd2939;
      102009:data<=16'd3277;
      102010:data<=16'd3333;
      102011:data<=16'd3930;
      102012:data<=16'd4059;
      102013:data<=16'd3321;
      102014:data<=16'd3814;
      102015:data<=16'd5392;
      102016:data<=16'd6143;
      102017:data<=16'd5755;
      102018:data<=16'd5607;
      102019:data<=16'd5715;
      102020:data<=16'd5332;
      102021:data<=16'd5979;
      102022:data<=16'd7200;
      102023:data<=16'd7319;
      102024:data<=16'd7788;
      102025:data<=16'd7890;
      102026:data<=16'd6542;
      102027:data<=16'd6300;
      102028:data<=16'd7200;
      102029:data<=16'd7934;
      102030:data<=16'd8511;
      102031:data<=16'd8061;
      102032:data<=16'd7145;
      102033:data<=16'd6799;
      102034:data<=16'd7150;
      102035:data<=16'd8275;
      102036:data<=16'd8634;
      102037:data<=16'd8046;
      102038:data<=16'd7947;
      102039:data<=16'd7852;
      102040:data<=16'd7568;
      102041:data<=16'd7741;
      102042:data<=16'd8605;
      102043:data<=16'd8954;
      102044:data<=16'd7999;
      102045:data<=16'd8331;
      102046:data<=16'd7153;
      102047:data<=16'd867;
      102048:data<=-16'd1577;
      102049:data<=16'd1158;
      102050:data<=-16'd1750;
      102051:data<=-16'd6713;
      102052:data<=-16'd6566;
      102053:data<=-16'd5896;
      102054:data<=-16'd5456;
      102055:data<=-16'd3419;
      102056:data<=-16'd2858;
      102057:data<=-16'd3509;
      102058:data<=-16'd2960;
      102059:data<=-16'd2698;
      102060:data<=-16'd3328;
      102061:data<=-16'd1983;
      102062:data<=16'd435;
      102063:data<=16'd466;
      102064:data<=16'd42;
      102065:data<=16'd382;
      102066:data<=-16'd372;
      102067:data<=-16'd353;
      102068:data<=16'd1007;
      102069:data<=16'd1635;
      102070:data<=16'd1789;
      102071:data<=16'd1905;
      102072:data<=16'd2268;
      102073:data<=16'd2472;
      102074:data<=16'd2455;
      102075:data<=16'd3764;
      102076:data<=16'd4299;
      102077:data<=16'd3424;
      102078:data<=16'd4126;
      102079:data<=16'd4234;
      102080:data<=16'd3007;
      102081:data<=16'd3747;
      102082:data<=16'd5319;
      102083:data<=16'd5921;
      102084:data<=16'd5600;
      102085:data<=16'd5045;
      102086:data<=16'd4987;
      102087:data<=16'd4842;
      102088:data<=16'd6241;
      102089:data<=16'd7298;
      102090:data<=16'd4899;
      102091:data<=16'd6821;
      102092:data<=16'd13524;
      102093:data<=16'd14515;
      102094:data<=16'd13220;
      102095:data<=16'd14924;
      102096:data<=16'd14754;
      102097:data<=16'd13694;
      102098:data<=16'd13941;
      102099:data<=16'd12695;
      102100:data<=16'd11145;
      102101:data<=16'd12088;
      102102:data<=16'd13913;
      102103:data<=16'd13494;
      102104:data<=16'd11831;
      102105:data<=16'd11300;
      102106:data<=16'd10912;
      102107:data<=16'd11116;
      102108:data<=16'd12207;
      102109:data<=16'd11705;
      102110:data<=16'd10800;
      102111:data<=16'd10881;
      102112:data<=16'd10627;
      102113:data<=16'd10569;
      102114:data<=16'd10246;
      102115:data<=16'd8922;
      102116:data<=16'd8734;
      102117:data<=16'd10806;
      102118:data<=16'd13359;
      102119:data<=16'd13805;
      102120:data<=16'd12689;
      102121:data<=16'd11611;
      102122:data<=16'd9544;
      102123:data<=16'd7847;
      102124:data<=16'd7761;
      102125:data<=16'd7501;
      102126:data<=16'd7799;
      102127:data<=16'd7239;
      102128:data<=16'd4137;
      102129:data<=16'd2922;
      102130:data<=16'd3568;
      102131:data<=16'd3107;
      102132:data<=16'd2995;
      102133:data<=16'd2281;
      102134:data<=16'd1230;
      102135:data<=16'd1095;
      102136:data<=-16'd2660;
      102137:data<=-16'd8561;
      102138:data<=-16'd10082;
      102139:data<=-16'd9365;
      102140:data<=-16'd9633;
      102141:data<=-16'd10120;
      102142:data<=-16'd11159;
      102143:data<=-16'd11609;
      102144:data<=-16'd10665;
      102145:data<=-16'd10185;
      102146:data<=-16'd10116;
      102147:data<=-16'd10313;
      102148:data<=-16'd11561;
      102149:data<=-16'd11782;
      102150:data<=-16'd10445;
      102151:data<=-16'd10386;
      102152:data<=-16'd11009;
      102153:data<=-16'd10255;
      102154:data<=-16'd9868;
      102155:data<=-16'd10971;
      102156:data<=-16'd11617;
      102157:data<=-16'd11154;
      102158:data<=-16'd10810;
      102159:data<=-16'd10649;
      102160:data<=-16'd10387;
      102161:data<=-16'd11069;
      102162:data<=-16'd12129;
      102163:data<=-16'd11677;
      102164:data<=-16'd10874;
      102165:data<=-16'd10763;
      102166:data<=-16'd9926;
      102167:data<=-16'd9512;
      102168:data<=-16'd10815;
      102169:data<=-16'd11458;
      102170:data<=-16'd11050;
      102171:data<=-16'd11065;
      102172:data<=-16'd10210;
      102173:data<=-16'd8666;
      102174:data<=-16'd9095;
      102175:data<=-16'd10610;
      102176:data<=-16'd10602;
      102177:data<=-16'd9451;
      102178:data<=-16'd8936;
      102179:data<=-16'd9368;
      102180:data<=-16'd8348;
      102181:data<=-16'd4613;
      102182:data<=-16'd1424;
      102183:data<=-16'd1146;
      102184:data<=-16'd3477;
      102185:data<=-16'd6799;
      102186:data<=-16'd7245;
      102187:data<=-16'd6008;
      102188:data<=-16'd7374;
      102189:data<=-16'd8125;
      102190:data<=-16'd6739;
      102191:data<=-16'd6868;
      102192:data<=-16'd6860;
      102193:data<=-16'd5799;
      102194:data<=-16'd6584;
      102195:data<=-16'd7941;
      102196:data<=-16'd7409;
      102197:data<=-16'd6147;
      102198:data<=-16'd6369;
      102199:data<=-16'd6663;
      102200:data<=-16'd5515;
      102201:data<=-16'd6228;
      102202:data<=-16'd7418;
      102203:data<=-16'd5653;
      102204:data<=-16'd5285;
      102205:data<=-16'd5979;
      102206:data<=-16'd4358;
      102207:data<=-16'd4675;
      102208:data<=-16'd6501;
      102209:data<=-16'd6049;
      102210:data<=-16'd5553;
      102211:data<=-16'd5767;
      102212:data<=-16'd5468;
      102213:data<=-16'd5031;
      102214:data<=-16'd5468;
      102215:data<=-16'd6625;
      102216:data<=-16'd6129;
      102217:data<=-16'd5338;
      102218:data<=-16'd5882;
      102219:data<=-16'd5277;
      102220:data<=-16'd4799;
      102221:data<=-16'd4805;
      102222:data<=-16'd3670;
      102223:data<=-16'd3425;
      102224:data<=-16'd2781;
      102225:data<=-16'd3541;
      102226:data<=-16'd9086;
      102227:data<=-16'd11177;
      102228:data<=-16'd8128;
      102229:data<=-16'd7480;
      102230:data<=-16'd7436;
      102231:data<=-16'd6625;
      102232:data<=-16'd6825;
      102233:data<=-16'd6302;
      102234:data<=-16'd5338;
      102235:data<=-16'd3850;
      102236:data<=-16'd2426;
      102237:data<=-16'd2654;
      102238:data<=-16'd2423;
      102239:data<=-16'd2129;
      102240:data<=-16'd1679;
      102241:data<=16'd681;
      102242:data<=16'd1333;
      102243:data<=16'd629;
      102244:data<=16'd1530;
      102245:data<=16'd1589;
      102246:data<=16'd1337;
      102247:data<=16'd2393;
      102248:data<=16'd3527;
      102249:data<=16'd4188;
      102250:data<=16'd4590;
      102251:data<=16'd7417;
      102252:data<=16'd10907;
      102253:data<=16'd10460;
      102254:data<=16'd10558;
      102255:data<=16'd12652;
      102256:data<=16'd12232;
      102257:data<=16'd11637;
      102258:data<=16'd11749;
      102259:data<=16'd10819;
      102260:data<=16'd11135;
      102261:data<=16'd12609;
      102262:data<=16'd13259;
      102263:data<=16'd12511;
      102264:data<=16'd11681;
      102265:data<=16'd12081;
      102266:data<=16'd11579;
      102267:data<=16'd11600;
      102268:data<=16'd13179;
      102269:data<=16'd12166;
      102270:data<=16'd13297;
      102271:data<=16'd19185;
      102272:data<=16'd20295;
      102273:data<=16'd18122;
      102274:data<=16'd19682;
      102275:data<=16'd20730;
      102276:data<=16'd19588;
      102277:data<=16'd19035;
      102278:data<=16'd18221;
      102279:data<=16'd17286;
      102280:data<=16'd17473;
      102281:data<=16'd18130;
      102282:data<=16'd17854;
      102283:data<=16'd16841;
      102284:data<=16'd16381;
      102285:data<=16'd15605;
      102286:data<=16'd14310;
      102287:data<=16'd14475;
      102288:data<=16'd15638;
      102289:data<=16'd15682;
      102290:data<=16'd14545;
      102291:data<=16'd13894;
      102292:data<=16'd13626;
      102293:data<=16'd12787;
      102294:data<=16'd13397;
      102295:data<=16'd14615;
      102296:data<=16'd13130;
      102297:data<=16'd11796;
      102298:data<=16'd12120;
      102299:data<=16'd11235;
      102300:data<=16'd10743;
      102301:data<=16'd11700;
      102302:data<=16'd11508;
      102303:data<=16'd10199;
      102304:data<=16'd9477;
      102305:data<=16'd9482;
      102306:data<=16'd8642;
      102307:data<=16'd7934;
      102308:data<=16'd9545;
      102309:data<=16'd9777;
      102310:data<=16'd7830;
      102311:data<=16'd7864;
      102312:data<=16'd7368;
      102313:data<=16'd6542;
      102314:data<=16'd8401;
      102315:data<=16'd5920;
      102316:data<=-16'd796;
      102317:data<=-16'd2629;
      102318:data<=-16'd3215;
      102319:data<=-16'd6405;
      102320:data<=-16'd6473;
      102321:data<=-16'd4529;
      102322:data<=-16'd4511;
      102323:data<=-16'd4522;
      102324:data<=-16'd4225;
      102325:data<=-16'd4523;
      102326:data<=-16'd4525;
      102327:data<=-16'd4428;
      102328:data<=-16'd4667;
      102329:data<=-16'd4796;
      102330:data<=-16'd4795;
      102331:data<=-16'd4754;
      102332:data<=-16'd4696;
      102333:data<=-16'd5304;
      102334:data<=-16'd6702;
      102335:data<=-16'd7430;
      102336:data<=-16'd6874;
      102337:data<=-16'd6338;
      102338:data<=-16'd6498;
      102339:data<=-16'd6774;
      102340:data<=-16'd7034;
      102341:data<=-16'd7759;
      102342:data<=-16'd8437;
      102343:data<=-16'd8178;
      102344:data<=-16'd7979;
      102345:data<=-16'd8163;
      102346:data<=-16'd7688;
      102347:data<=-16'd7818;
      102348:data<=-16'd8769;
      102349:data<=-16'd8831;
      102350:data<=-16'd8828;
      102351:data<=-16'd8634;
      102352:data<=-16'd7647;
      102353:data<=-16'd8088;
      102354:data<=-16'd9324;
      102355:data<=-16'd9489;
      102356:data<=-16'd9274;
      102357:data<=-16'd8868;
      102358:data<=-16'd9241;
      102359:data<=-16'd8757;
      102360:data<=-16'd4350;
      102361:data<=-16'd1392;
      102362:data<=-16'd2692;
      102363:data<=-16'd2511;
      102364:data<=-16'd1632;
      102365:data<=-16'd2282;
      102366:data<=-16'd1712;
      102367:data<=-16'd1956;
      102368:data<=-16'd3841;
      102369:data<=-16'd3782;
      102370:data<=-16'd3275;
      102371:data<=-16'd3723;
      102372:data<=-16'd3230;
      102373:data<=-16'd3453;
      102374:data<=-16'd5432;
      102375:data<=-16'd6061;
      102376:data<=-16'd5200;
      102377:data<=-16'd5447;
      102378:data<=-16'd5568;
      102379:data<=-16'd4387;
      102380:data<=-16'd4811;
      102381:data<=-16'd6733;
      102382:data<=-16'd7069;
      102383:data<=-16'd6451;
      102384:data<=-16'd5588;
      102385:data<=-16'd3347;
      102386:data<=-16'd1636;
      102387:data<=-16'd2619;
      102388:data<=-16'd3868;
      102389:data<=-16'd3281;
      102390:data<=-16'd3087;
      102391:data<=-16'd3688;
      102392:data<=-16'd3303;
      102393:data<=-16'd3865;
      102394:data<=-16'd5380;
      102395:data<=-16'd5074;
      102396:data<=-16'd4921;
      102397:data<=-16'd5591;
      102398:data<=-16'd4951;
      102399:data<=-16'd4599;
      102400:data<=-16'd5339;
      102401:data<=-16'd6499;
      102402:data<=-16'd7106;
      102403:data<=-16'd5686;
      102404:data<=-16'd6862;
      102405:data<=-16'd12424;
      102406:data<=-16'd15153;
      102407:data<=-16'd14868;
      102408:data<=-16'd15303;
      102409:data<=-16'd14727;
      102410:data<=-16'd14166;
      102411:data<=-16'd14325;
      102412:data<=-16'd13546;
      102413:data<=-16'd13729;
      102414:data<=-16'd14540;
      102415:data<=-16'd14001;
      102416:data<=-16'd13320;
      102417:data<=-16'd12753;
      102418:data<=-16'd12046;
      102419:data<=-16'd11617;
      102420:data<=-16'd11708;
      102421:data<=-16'd12486;
      102422:data<=-16'd12413;
      102423:data<=-16'd11494;
      102424:data<=-16'd11215;
      102425:data<=-16'd10684;
      102426:data<=-16'd10525;
      102427:data<=-16'd11470;
      102428:data<=-16'd11461;
      102429:data<=-16'd10821;
      102430:data<=-16'd10549;
      102431:data<=-16'd9741;
      102432:data<=-16'd8869;
      102433:data<=-16'd8725;
      102434:data<=-16'd8655;
      102435:data<=-16'd7764;
      102436:data<=-16'd6696;
      102437:data<=-16'd6243;
      102438:data<=-16'd5524;
      102439:data<=-16'd5219;
      102440:data<=-16'd5072;
      102441:data<=-16'd3209;
      102442:data<=-16'd2391;
      102443:data<=-16'd2875;
      102444:data<=-16'd1739;
      102445:data<=-16'd1536;
      102446:data<=-16'd1304;
      102447:data<=16'd557;
      102448:data<=-16'd141;
      102449:data<=16'd1497;
      102450:data<=16'd8483;
      102451:data<=16'd10144;
      102452:data<=16'd6267;
      102453:data<=16'd5419;
      102454:data<=16'd6458;
      102455:data<=16'd6940;
      102456:data<=16'd7360;
      102457:data<=16'd7456;
      102458:data<=16'd7370;
      102459:data<=16'd6731;
      102460:data<=16'd6810;
      102461:data<=16'd8235;
      102462:data<=16'd8363;
      102463:data<=16'd7746;
      102464:data<=16'd8026;
      102465:data<=16'd7764;
      102466:data<=16'd7456;
      102467:data<=16'd8526;
      102468:data<=16'd9497;
      102469:data<=16'd9053;
      102470:data<=16'd8507;
      102471:data<=16'd8530;
      102472:data<=16'd7882;
      102473:data<=16'd7884;
      102474:data<=16'd9758;
      102475:data<=16'd10461;
      102476:data<=16'd9288;
      102477:data<=16'd8548;
      102478:data<=16'd8420;
      102479:data<=16'd8801;
      102480:data<=16'd9561;
      102481:data<=16'd9746;
      102482:data<=16'd9109;
      102483:data<=16'd8334;
      102484:data<=16'd8267;
      102485:data<=16'd7971;
      102486:data<=16'd8000;
      102487:data<=16'd10160;
      102488:data<=16'd10604;
      102489:data<=16'd8661;
      102490:data<=16'd9256;
      102491:data<=16'd9367;
      102492:data<=16'd7682;
      102493:data<=16'd8939;
      102494:data<=16'd8064;
      102495:data<=16'd2115;
      102496:data<=-16'd694;
      102497:data<=16'd329;
      102498:data<=16'd262;
      102499:data<=16'd293;
      102500:data<=16'd1704;
      102501:data<=16'd2631;
      102502:data<=16'd2130;
      102503:data<=16'd1636;
      102504:data<=16'd1952;
      102505:data<=16'd1817;
      102506:data<=16'd1950;
      102507:data<=16'd3189;
      102508:data<=16'd3535;
      102509:data<=16'd3133;
      102510:data<=16'd3466;
      102511:data<=16'd3369;
      102512:data<=16'd2690;
      102513:data<=16'd3339;
      102514:data<=16'd4990;
      102515:data<=16'd5518;
      102516:data<=16'd4916;
      102517:data<=16'd4429;
      102518:data<=16'd4690;
      102519:data<=16'd6724;
      102520:data<=16'd9379;
      102521:data<=16'd9844;
      102522:data<=16'd9209;
      102523:data<=16'd9238;
      102524:data<=16'd8845;
      102525:data<=16'd8281;
      102526:data<=16'd8831;
      102527:data<=16'd9991;
      102528:data<=16'd10119;
      102529:data<=16'd9198;
      102530:data<=16'd9195;
      102531:data<=16'd9062;
      102532:data<=16'd7661;
      102533:data<=16'd8232;
      102534:data<=16'd9911;
      102535:data<=16'd9411;
      102536:data<=16'd8737;
      102537:data<=16'd8084;
      102538:data<=16'd7635;
      102539:data<=16'd11392;
      102540:data<=16'd15775;
      102541:data<=16'd15399;
      102542:data<=16'd14267;
      102543:data<=16'd14246;
      102544:data<=16'd12837;
      102545:data<=16'd11656;
      102546:data<=16'd11124;
      102547:data<=16'd9606;
      102548:data<=16'd8630;
      102549:data<=16'd8551;
      102550:data<=16'd7783;
      102551:data<=16'd7133;
      102552:data<=16'd7021;
      102553:data<=16'd5839;
      102554:data<=16'd4000;
      102555:data<=16'd3263;
      102556:data<=16'd2933;
      102557:data<=16'd2273;
      102558:data<=16'd2419;
      102559:data<=16'd2361;
      102560:data<=16'd761;
      102561:data<=-16'd211;
      102562:data<=16'd91;
      102563:data<=-16'd85;
      102564:data<=-16'd209;
      102565:data<=-16'd6;
      102566:data<=-16'd755;
      102567:data<=-16'd1964;
      102568:data<=-16'd2555;
      102569:data<=-16'd2684;
      102570:data<=-16'd2861;
      102571:data<=-16'd3022;
      102572:data<=-16'd2872;
      102573:data<=-16'd3463;
      102574:data<=-16'd5074;
      102575:data<=-16'd5530;
      102576:data<=-16'd4860;
      102577:data<=-16'd5040;
      102578:data<=-16'd5022;
      102579:data<=-16'd4578;
      102580:data<=-16'd6264;
      102581:data<=-16'd7735;
      102582:data<=-16'd6143;
      102583:data<=-16'd7121;
      102584:data<=-16'd12481;
      102585:data<=-16'd15744;
      102586:data<=-16'd17511;
      102587:data<=-16'd20380;
      102588:data<=-16'd20324;
      102589:data<=-16'd18404;
      102590:data<=-16'd18155;
      102591:data<=-16'd17655;
      102592:data<=-16'd17229;
      102593:data<=-16'd18127;
      102594:data<=-16'd18431;
      102595:data<=-16'd17787;
      102596:data<=-16'd16939;
      102597:data<=-16'd16126;
      102598:data<=-16'd15434;
      102599:data<=-16'd15135;
      102600:data<=-16'd15855;
      102601:data<=-16'd15869;
      102602:data<=-16'd14477;
      102603:data<=-16'd13943;
      102604:data<=-16'd13520;
      102605:data<=-16'd12649;
      102606:data<=-16'd13212;
      102607:data<=-16'd13957;
      102608:data<=-16'd13653;
      102609:data<=-16'd13330;
      102610:data<=-16'd12787;
      102611:data<=-16'd11903;
      102612:data<=-16'd11681;
      102613:data<=-16'd12264;
      102614:data<=-16'd12138;
      102615:data<=-16'd11154;
      102616:data<=-16'd10892;
      102617:data<=-16'd10378;
      102618:data<=-16'd9379;
      102619:data<=-16'd9600;
      102620:data<=-16'd9931;
      102621:data<=-16'd9917;
      102622:data<=-16'd9697;
      102623:data<=-16'd8542;
      102624:data<=-16'd7991;
      102625:data<=-16'd7520;
      102626:data<=-16'd7614;
      102627:data<=-16'd9949;
      102628:data<=-16'd7694;
      102629:data<=-16'd458;
      102630:data<=16'd1726;
      102631:data<=16'd588;
      102632:data<=16'd831;
      102633:data<=-16'd399;
      102634:data<=-16'd1202;
      102635:data<=-16'd243;
      102636:data<=-16'd390;
      102637:data<=-16'd553;
      102638:data<=-16'd18;
      102639:data<=-16'd635;
      102640:data<=-16'd2199;
      102641:data<=-16'd2673;
      102642:data<=-16'd1575;
      102643:data<=-16'd755;
      102644:data<=-16'd552;
      102645:data<=-16'd657;
      102646:data<=-16'd1199;
      102647:data<=-16'd796;
      102648:data<=-16'd256;
      102649:data<=-16'd250;
      102650:data<=16'd591;
      102651:data<=16'd584;
      102652:data<=16'd1196;
      102653:data<=16'd5407;
      102654:data<=16'd8334;
      102655:data<=16'd7635;
      102656:data<=16'd7260;
      102657:data<=16'd7732;
      102658:data<=16'd7739;
      102659:data<=16'd7732;
      102660:data<=16'd8526;
      102661:data<=16'd9063;
      102662:data<=16'd8493;
      102663:data<=16'd8851;
      102664:data<=16'd8799;
      102665:data<=16'd7104;
      102666:data<=16'd7844;
      102667:data<=16'd9591;
      102668:data<=16'd9230;
      102669:data<=16'd9089;
      102670:data<=16'd8525;
      102671:data<=16'd8094;
      102672:data<=16'd9271;
      102673:data<=16'd6975;
      102674:data<=16'd1835;
      102675:data<=16'd118;
      102676:data<=16'd757;
      102677:data<=16'd1131;
      102678:data<=16'd1389;
      102679:data<=16'd1485;
      102680:data<=16'd2347;
      102681:data<=16'd3563;
      102682:data<=16'd3471;
      102683:data<=16'd2917;
      102684:data<=16'd3045;
      102685:data<=16'd3243;
      102686:data<=16'd3941;
      102687:data<=16'd5474;
      102688:data<=16'd5447;
      102689:data<=16'd4156;
      102690:data<=16'd4540;
      102691:data<=16'd5112;
      102692:data<=16'd5200;
      102693:data<=16'd6664;
      102694:data<=16'd6989;
      102695:data<=16'd5708;
      102696:data<=16'd5994;
      102697:data<=16'd6328;
      102698:data<=16'd5409;
      102699:data<=16'd5762;
      102700:data<=16'd7453;
      102701:data<=16'd7871;
      102702:data<=16'd6746;
      102703:data<=16'd6510;
      102704:data<=16'd6872;
      102705:data<=16'd6529;
      102706:data<=16'd7580;
      102707:data<=16'd8810;
      102708:data<=16'd7674;
      102709:data<=16'd7198;
      102710:data<=16'd7553;
      102711:data<=16'd6693;
      102712:data<=16'd7013;
      102713:data<=16'd8260;
      102714:data<=16'd8593;
      102715:data<=16'd8718;
      102716:data<=16'd7761;
      102717:data<=16'd7824;
      102718:data<=16'd12014;
      102719:data<=16'd15100;
      102720:data<=16'd13420;
      102721:data<=16'd11653;
      102722:data<=16'd11568;
      102723:data<=16'd10991;
      102724:data<=16'd10302;
      102725:data<=16'd10442;
      102726:data<=16'd10985;
      102727:data<=16'd11185;
      102728:data<=16'd10774;
      102729:data<=16'd10396;
      102730:data<=16'd9868;
      102731:data<=16'd8831;
      102732:data<=16'd8636;
      102733:data<=16'd9447;
      102734:data<=16'd9715;
      102735:data<=16'd9367;
      102736:data<=16'd8863;
      102737:data<=16'd7888;
      102738:data<=16'd7260;
      102739:data<=16'd8322;
      102740:data<=16'd9685;
      102741:data<=16'd9260;
      102742:data<=16'd8445;
      102743:data<=16'd8281;
      102744:data<=16'd7524;
      102745:data<=16'd7456;
      102746:data<=16'd8849;
      102747:data<=16'd9086;
      102748:data<=16'd8220;
      102749:data<=16'd7941;
      102750:data<=16'd7201;
      102751:data<=16'd6047;
      102752:data<=16'd6141;
      102753:data<=16'd6331;
      102754:data<=16'd5344;
      102755:data<=16'd4807;
      102756:data<=16'd4640;
      102757:data<=16'd3982;
      102758:data<=16'd3932;
      102759:data<=16'd2734;
      102760:data<=16'd749;
      102761:data<=16'd1334;
      102762:data<=-16'd879;
      102763:data<=-16'd7515;
      102764:data<=-16'd9462;
      102765:data<=-16'd8393;
      102766:data<=-16'd10099;
      102767:data<=-16'd10928;
      102768:data<=-16'd10652;
      102769:data<=-16'd10710;
      102770:data<=-16'd10006;
      102771:data<=-16'd10131;
      102772:data<=-16'd10411;
      102773:data<=-16'd10605;
      102774:data<=-16'd11558;
      102775:data<=-16'd10836;
      102776:data<=-16'd10146;
      102777:data<=-16'd10696;
      102778:data<=-16'd9890;
      102779:data<=-16'd10232;
      102780:data<=-16'd11712;
      102781:data<=-16'd11217;
      102782:data<=-16'd10828;
      102783:data<=-16'd10633;
      102784:data<=-16'd10037;
      102785:data<=-16'd10783;
      102786:data<=-16'd10643;
      102787:data<=-16'd8393;
      102788:data<=-16'd6672;
      102789:data<=-16'd6536;
      102790:data<=-16'd6868;
      102791:data<=-16'd6579;
      102792:data<=-16'd6936;
      102793:data<=-16'd8282;
      102794:data<=-16'd8345;
      102795:data<=-16'd7694;
      102796:data<=-16'd7918;
      102797:data<=-16'd8019;
      102798:data<=-16'd7468;
      102799:data<=-16'd7924;
      102800:data<=-16'd9555;
      102801:data<=-16'd9010;
      102802:data<=-16'd7395;
      102803:data<=-16'd7975;
      102804:data<=-16'd7614;
      102805:data<=-16'd7953;
      102806:data<=-16'd10813;
      102807:data<=-16'd7512;
      102808:data<=-16'd851;
      102809:data<=-16'd607;
      102810:data<=-16'd1228;
      102811:data<=16'd274;
      102812:data<=-16'd931;
      102813:data<=-16'd2705;
      102814:data<=-16'd2761;
      102815:data<=-16'd2276;
      102816:data<=-16'd2077;
      102817:data<=-16'd2384;
      102818:data<=-16'd2400;
      102819:data<=-16'd3363;
      102820:data<=-16'd4896;
      102821:data<=-16'd4481;
      102822:data<=-16'd4023;
      102823:data<=-16'd4350;
      102824:data<=-16'd3973;
      102825:data<=-16'd4219;
      102826:data<=-16'd5239;
      102827:data<=-16'd5820;
      102828:data<=-16'd5791;
      102829:data<=-16'd5621;
      102830:data<=-16'd5673;
      102831:data<=-16'd4908;
      102832:data<=-16'd4825;
      102833:data<=-16'd6771;
      102834:data<=-16'd7097;
      102835:data<=-16'd5826;
      102836:data<=-16'd5680;
      102837:data<=-16'd5180;
      102838:data<=-16'd4660;
      102839:data<=-16'd5846;
      102840:data<=-16'd6907;
      102841:data<=-16'd6343;
      102842:data<=-16'd5882;
      102843:data<=-16'd6473;
      102844:data<=-16'd5937;
      102845:data<=-16'd5579;
      102846:data<=-16'd7574;
      102847:data<=-16'd8058;
      102848:data<=-16'd7285;
      102849:data<=-16'd7409;
      102850:data<=-16'd5662;
      102851:data<=-16'd6730;
      102852:data<=-16'd13591;
      102853:data<=-16'd18039;
      102854:data<=-16'd19124;
      102855:data<=-16'd20118;
      102856:data<=-16'd19338;
      102857:data<=-16'd18221;
      102858:data<=-16'd17606;
      102859:data<=-16'd16537;
      102860:data<=-16'd15910;
      102861:data<=-16'd14944;
      102862:data<=-16'd13973;
      102863:data<=-16'd13617;
      102864:data<=-16'd12652;
      102865:data<=-16'd11649;
      102866:data<=-16'd10193;
      102867:data<=-16'd8486;
      102868:data<=-16'd8263;
      102869:data<=-16'd7765;
      102870:data<=-16'd7097;
      102871:data<=-16'd7319;
      102872:data<=-16'd5562;
      102873:data<=-16'd2922;
      102874:data<=-16'd2378;
      102875:data<=-16'd2373;
      102876:data<=-16'd2314;
      102877:data<=-16'd2663;
      102878:data<=-16'd2015;
      102879:data<=-16'd147;
      102880:data<=16'd1071;
      102881:data<=16'd837;
      102882:data<=16'd737;
      102883:data<=16'd1140;
      102884:data<=16'd1372;
      102885:data<=16'd2325;
      102886:data<=16'd3571;
      102887:data<=16'd4105;
      102888:data<=16'd4275;
      102889:data<=16'd4219;
      102890:data<=16'd4684;
      102891:data<=16'd5028;
      102892:data<=16'd4998;
      102893:data<=16'd6821;
      102894:data<=16'd7262;
      102895:data<=16'd5131;
      102896:data<=16'd8308;
      102897:data<=16'd14700;
      102898:data<=16'd15825;
      102899:data<=16'd15397;
      102900:data<=16'd16493;
      102901:data<=16'd15802;
      102902:data<=16'd14819;
      102903:data<=16'd14713;
      102904:data<=16'd14040;
      102905:data<=16'd13944;
      102906:data<=16'd14647;
      102907:data<=16'd14838;
      102908:data<=16'd14407;
      102909:data<=16'd13840;
      102910:data<=16'd13439;
      102911:data<=16'd13179;
      102912:data<=16'd13737;
      102913:data<=16'd14662;
      102914:data<=16'd14014;
      102915:data<=16'd12910;
      102916:data<=16'd12774;
      102917:data<=16'd12487;
      102918:data<=16'd12495;
      102919:data<=16'd13235;
      102920:data<=16'd14270;
      102921:data<=16'd16076;
      102922:data<=16'd17111;
      102923:data<=16'd16114;
      102924:data<=16'd15027;
      102925:data<=16'd15311;
      102926:data<=16'd16472;
      102927:data<=16'd16551;
      102928:data<=16'd14998;
      102929:data<=16'd13881;
      102930:data<=16'd13382;
      102931:data<=16'd13235;
      102932:data<=16'd14040;
      102933:data<=16'd14189;
      102934:data<=16'd13259;
      102935:data<=16'd12584;
      102936:data<=16'd11982;
      102937:data<=16'd11206;
      102938:data<=16'd10915;
      102939:data<=16'd11964;
      102940:data<=16'd11262;
      102941:data<=16'd5648;
      102942:data<=16'd1383;
      102943:data<=16'd1591;
      102944:data<=16'd952;
      102945:data<=16'd1180;
      102946:data<=16'd3448;
      102947:data<=16'd3169;
      102948:data<=16'd2394;
      102949:data<=16'd2499;
      102950:data<=16'd1656;
      102951:data<=16'd2228;
      102952:data<=16'd3532;
      102953:data<=16'd3477;
      102954:data<=16'd3294;
      102955:data<=16'd2943;
      102956:data<=16'd2651;
      102957:data<=16'd2614;
      102958:data<=16'd2896;
      102959:data<=16'd4205;
      102960:data<=16'd4261;
      102961:data<=16'd3213;
      102962:data<=16'd3359;
      102963:data<=16'd2842;
      102964:data<=16'd2243;
      102965:data<=16'd2863;
      102966:data<=16'd2376;
      102967:data<=16'd1516;
      102968:data<=16'd1290;
      102969:data<=16'd1030;
      102970:data<=16'd1321;
      102971:data<=16'd561;
      102972:data<=-16'd1657;
      102973:data<=-16'd2402;
      102974:data<=-16'd1575;
      102975:data<=-16'd1457;
      102976:data<=-16'd2224;
      102977:data<=-16'd2217;
      102978:data<=-16'd2519;
      102979:data<=-16'd4429;
      102980:data<=-16'd4934;
      102981:data<=-16'd4397;
      102982:data<=-16'd4795;
      102983:data<=-16'd4393;
      102984:data<=-16'd4780;
      102985:data<=-16'd4128;
      102986:data<=16'd793;
      102987:data<=16'd1582;
      102988:data<=-16'd2881;
      102989:data<=-16'd3369;
      102990:data<=-16'd2519;
      102991:data<=-16'd4249;
      102992:data<=-16'd5403;
      102993:data<=-16'd5824;
      102994:data<=-16'd5509;
      102995:data<=-16'd5095;
      102996:data<=-16'd5697;
      102997:data<=-16'd5474;
      102998:data<=-16'd5697;
      102999:data<=-16'd7104;
      103000:data<=-16'd6995;
      103001:data<=-16'd6529;
      103002:data<=-16'd7027;
      103003:data<=-16'd6974;
      103004:data<=-16'd6475;
      103005:data<=-16'd6839;
      103006:data<=-16'd8069;
      103007:data<=-16'd8317;
      103008:data<=-16'd7739;
      103009:data<=-16'd8014;
      103010:data<=-16'd7870;
      103011:data<=-16'd7749;
      103012:data<=-16'd9109;
      103013:data<=-16'd9420;
      103014:data<=-16'd8457;
      103015:data<=-16'd8325;
      103016:data<=-16'd8058;
      103017:data<=-16'd7374;
      103018:data<=-16'd8102;
      103019:data<=-16'd9981;
      103020:data<=-16'd10272;
      103021:data<=-16'd9059;
      103022:data<=-16'd8772;
      103023:data<=-16'd8378;
      103024:data<=-16'd7993;
      103025:data<=-16'd9492;
      103026:data<=-16'd10223;
      103027:data<=-16'd9426;
      103028:data<=-16'd8810;
      103029:data<=-16'd8257;
      103030:data<=-16'd10652;
      103031:data<=-16'd15306;
      103032:data<=-16'd16460;
      103033:data<=-16'd15396;
      103034:data<=-16'd15112;
      103035:data<=-16'd14468;
      103036:data<=-16'd13391;
      103037:data<=-16'd12372;
      103038:data<=-16'd12719;
      103039:data<=-16'd14158;
      103040:data<=-16'd13597;
      103041:data<=-16'd12173;
      103042:data<=-16'd11627;
      103043:data<=-16'd10604;
      103044:data<=-16'd10498;
      103045:data<=-16'd11679;
      103046:data<=-16'd11574;
      103047:data<=-16'd10625;
      103048:data<=-16'd10223;
      103049:data<=-16'd9940;
      103050:data<=-16'd9379;
      103051:data<=-16'd8915;
      103052:data<=-16'd9394;
      103053:data<=-16'd9858;
      103054:data<=-16'd8026;
      103055:data<=-16'd4840;
      103056:data<=-16'd3115;
      103057:data<=-16'd2919;
      103058:data<=-16'd3463;
      103059:data<=-16'd4563;
      103060:data<=-16'd4661;
      103061:data<=-16'd3862;
      103062:data<=-16'd3641;
      103063:data<=-16'd2971;
      103064:data<=-16'd2713;
      103065:data<=-16'd4082;
      103066:data<=-16'd4258;
      103067:data<=-16'd3624;
      103068:data<=-16'd3847;
      103069:data<=-16'd3240;
      103070:data<=-16'd2792;
      103071:data<=-16'd2786;
      103072:data<=-16'd2256;
      103073:data<=-16'd2919;
      103074:data<=-16'd1401;
      103075:data<=16'd4131;
      103076:data<=16'd6561;
      103077:data<=16'd5462;
      103078:data<=16'd6423;
      103079:data<=16'd8076;
      103080:data<=16'd7931;
      103081:data<=16'd7412;
      103082:data<=16'd7580;
      103083:data<=16'd7741;
      103084:data<=16'd7794;
      103085:data<=16'd8739;
      103086:data<=16'd9427;
      103087:data<=16'd8948;
      103088:data<=16'd9044;
      103089:data<=16'd9353;
      103090:data<=16'd8963;
      103091:data<=16'd9227;
      103092:data<=16'd10188;
      103093:data<=16'd10627;
      103094:data<=16'd10425;
      103095:data<=16'd10384;
      103096:data<=16'd10025;
      103097:data<=16'd9016;
      103098:data<=16'd9788;
      103099:data<=16'd11330;
      103100:data<=16'd10677;
      103101:data<=16'd10390;
      103102:data<=16'd10710;
      103103:data<=16'd9580;
      103104:data<=16'd9937;
      103105:data<=16'd11512;
      103106:data<=16'd11374;
      103107:data<=16'd10675;
      103108:data<=16'd10295;
      103109:data<=16'd10254;
      103110:data<=16'd10013;
      103111:data<=16'd9588;
      103112:data<=16'd10843;
      103113:data<=16'd11461;
      103114:data<=16'd10342;
      103115:data<=16'd10586;
      103116:data<=16'd10091;
      103117:data<=16'd9215;
      103118:data<=16'd11153;
      103119:data<=16'd10379;
      103120:data<=16'd5424;
      103121:data<=16'd2237;
      103122:data<=16'd303;
      103123:data<=-16'd1424;
      103124:data<=-16'd593;
      103125:data<=16'd1424;
      103126:data<=16'd1959;
      103127:data<=16'd1377;
      103128:data<=16'd1745;
      103129:data<=16'd2355;
      103130:data<=16'd1572;
      103131:data<=16'd1965;
      103132:data<=16'd3688;
      103133:data<=16'd3691;
      103134:data<=16'd3307;
      103135:data<=16'd3406;
      103136:data<=16'd2769;
      103137:data<=16'd2878;
      103138:data<=16'd4079;
      103139:data<=16'd4831;
      103140:data<=16'd4854;
      103141:data<=16'd4576;
      103142:data<=16'd4437;
      103143:data<=16'd4262;
      103144:data<=16'd4684;
      103145:data<=16'd5990;
      103146:data<=16'd6026;
      103147:data<=16'd5382;
      103148:data<=16'd5800;
      103149:data<=16'd5056;
      103150:data<=16'd3573;
      103151:data<=16'd4632;
      103152:data<=16'd6711;
      103153:data<=16'd6842;
      103154:data<=16'd5846;
      103155:data<=16'd5429;
      103156:data<=16'd5285;
      103157:data<=16'd5438;
      103158:data<=16'd6646;
      103159:data<=16'd7154;
      103160:data<=16'd6476;
      103161:data<=16'd6402;
      103162:data<=16'd5595;
      103163:data<=16'd5529;
      103164:data<=16'd9911;
      103165:data<=16'd13800;
      103166:data<=16'd13232;
      103167:data<=16'd12507;
      103168:data<=16'd12410;
      103169:data<=16'd11048;
      103170:data<=16'd10128;
      103171:data<=16'd10775;
      103172:data<=16'd11800;
      103173:data<=16'd11512;
      103174:data<=16'd10313;
      103175:data<=16'd9931;
      103176:data<=16'd9759;
      103177:data<=16'd9371;
      103178:data<=16'd9025;
      103179:data<=16'd8108;
      103180:data<=16'd7454;
      103181:data<=16'd7124;
      103182:data<=16'd6669;
      103183:data<=16'd6768;
      103184:data<=16'd5554;
      103185:data<=16'd3262;
      103186:data<=16'd2728;
      103187:data<=16'd2382;
      103188:data<=16'd2561;
      103189:data<=16'd5366;
      103190:data<=16'd6871;
      103191:data<=16'd5142;
      103192:data<=16'd3178;
      103193:data<=16'd2174;
      103194:data<=16'd1950;
      103195:data<=16'd1835;
      103196:data<=16'd1551;
      103197:data<=16'd1027;
      103198:data<=-16'd631;
      103199:data<=-16'd1760;
      103200:data<=-16'd1366;
      103201:data<=-16'd1770;
      103202:data<=-16'd2601;
      103203:data<=-16'd2397;
      103204:data<=-16'd2632;
      103205:data<=-16'd4244;
      103206:data<=-16'd5083;
      103207:data<=-16'd4140;
      103208:data<=-16'd5859;
      103209:data<=-16'd10522;
      103210:data<=-16'd11721;
      103211:data<=-16'd11402;
      103212:data<=-16'd13405;
      103213:data<=-16'd13464;
      103214:data<=-16'd12155;
      103215:data<=-16'd12320;
      103216:data<=-16'd11781;
      103217:data<=-16'd11749;
      103218:data<=-16'd13156;
      103219:data<=-16'd13480;
      103220:data<=-16'd13016;
      103221:data<=-16'd12659;
      103222:data<=-16'd12458;
      103223:data<=-16'd12210;
      103224:data<=-16'd11941;
      103225:data<=-16'd13054;
      103226:data<=-16'd13867;
      103227:data<=-16'd12792;
      103228:data<=-16'd12231;
      103229:data<=-16'd11787;
      103230:data<=-16'd11186;
      103231:data<=-16'd12492;
      103232:data<=-16'd13376;
      103233:data<=-16'd12283;
      103234:data<=-16'd11737;
      103235:data<=-16'd11826;
      103236:data<=-16'd11411;
      103237:data<=-16'd11421;
      103238:data<=-16'd12345;
      103239:data<=-16'd12578;
      103240:data<=-16'd11847;
      103241:data<=-16'd11908;
      103242:data<=-16'd11676;
      103243:data<=-16'd10361;
      103244:data<=-16'd10693;
      103245:data<=-16'd12161;
      103246:data<=-16'd12005;
      103247:data<=-16'd10831;
      103248:data<=-16'd10137;
      103249:data<=-16'd9908;
      103250:data<=-16'd9841;
      103251:data<=-16'd10980;
      103252:data<=-16'd11873;
      103253:data<=-16'd8056;
      103254:data<=-16'd3115;
      103255:data<=-16'd4034;
      103256:data<=-16'd7241;
      103257:data<=-16'd8141;
      103258:data<=-16'd8725;
      103259:data<=-16'd9222;
      103260:data<=-16'd8763;
      103261:data<=-16'd8264;
      103262:data<=-16'd7430;
      103263:data<=-16'd6311;
      103264:data<=-16'd6772;
      103265:data<=-16'd8473;
      103266:data<=-16'd8551;
      103267:data<=-16'd7397;
      103268:data<=-16'd7241;
      103269:data<=-16'd7244;
      103270:data<=-16'd7283;
      103271:data<=-16'd8225;
      103272:data<=-16'd8490;
      103273:data<=-16'd7733;
      103274:data<=-16'd7230;
      103275:data<=-16'd7078;
      103276:data<=-16'd6978;
      103277:data<=-16'd6899;
      103278:data<=-16'd7301;
      103279:data<=-16'd7559;
      103280:data<=-16'd6963;
      103281:data<=-16'd6768;
      103282:data<=-16'd6507;
      103283:data<=-16'd5708;
      103284:data<=-16'd5785;
      103285:data<=-16'd5527;
      103286:data<=-16'd4499;
      103287:data<=-16'd3996;
      103288:data<=-16'd3527;
      103289:data<=-16'd3660;
      103290:data<=-16'd3432;
      103291:data<=-16'd1362;
      103292:data<=-16'd217;
      103293:data<=-16'd294;
      103294:data<=-16'd173;
      103295:data<=-16'd199;
      103296:data<=16'd713;
      103297:data<=16'd325;
      103298:data<=-16'd2614;
      103299:data<=-16'd3404;
      103300:data<=-16'd2638;
      103301:data<=-16'd2864;
      103302:data<=-16'd2362;
      103303:data<=-16'd2017;
      103304:data<=-16'd1600;
      103305:data<=16'd261;
      103306:data<=16'd920;
      103307:data<=16'd597;
      103308:data<=16'd1115;
      103309:data<=16'd1193;
      103310:data<=16'd1695;
      103311:data<=16'd3563;
      103312:data<=16'd4410;
      103313:data<=16'd4011;
      103314:data<=16'd4416;
      103315:data<=16'd4714;
      103316:data<=16'd3962;
      103317:data<=16'd4585;
      103318:data<=16'd6441;
      103319:data<=16'd6939;
      103320:data<=16'd6569;
      103321:data<=16'd6275;
      103322:data<=16'd7282;
      103323:data<=16'd10410;
      103324:data<=16'd12463;
      103325:data<=16'd12674;
      103326:data<=16'd12847;
      103327:data<=16'd12125;
      103328:data<=16'd11314;
      103329:data<=16'd11100;
      103330:data<=16'd11041;
      103331:data<=16'd12419;
      103332:data<=16'd12977;
      103333:data<=16'd11737;
      103334:data<=16'd12007;
      103335:data<=16'd12216;
      103336:data<=16'd11285;
      103337:data<=16'd11702;
      103338:data<=16'd12731;
      103339:data<=16'd13524;
      103340:data<=16'd12891;
      103341:data<=16'd11032;
      103342:data<=16'd12921;
      103343:data<=16'd17414;
      103344:data<=16'd19015;
      103345:data<=16'd18635;
      103346:data<=16'd17987;
      103347:data<=16'd17118;
      103348:data<=16'd16577;
      103349:data<=16'd15838;
      103350:data<=16'd15620;
      103351:data<=16'd16299;
      103352:data<=16'd16075;
      103353:data<=16'd15024;
      103354:data<=16'd14590;
      103355:data<=16'd14407;
      103356:data<=16'd13353;
      103357:data<=16'd12891;
      103358:data<=16'd14143;
      103359:data<=16'd14025;
      103360:data<=16'd12437;
      103361:data<=16'd12002;
      103362:data<=16'd11091;
      103363:data<=16'd10194;
      103364:data<=16'd11215;
      103365:data<=16'd11491;
      103366:data<=16'd10675;
      103367:data<=16'd10235;
      103368:data<=16'd9482;
      103369:data<=16'd8950;
      103370:data<=16'd8942;
      103371:data<=16'd9418;
      103372:data<=16'd10075;
      103373:data<=16'd9385;
      103374:data<=16'd8614;
      103375:data<=16'd8361;
      103376:data<=16'd7300;
      103377:data<=16'd7447;
      103378:data<=16'd8561;
      103379:data<=16'd8147;
      103380:data<=16'd7303;
      103381:data<=16'd6586;
      103382:data<=16'd6117;
      103383:data<=16'd6287;
      103384:data<=16'd6526;
      103385:data<=16'd7248;
      103386:data<=16'd5629;
      103387:data<=16'd816;
      103388:data<=-16'd1284;
      103389:data<=-16'd2076;
      103390:data<=-16'd5318;
      103391:data<=-16'd6376;
      103392:data<=-16'd5600;
      103393:data<=-16'd6481;
      103394:data<=-16'd6704;
      103395:data<=-16'd6202;
      103396:data<=-16'd6115;
      103397:data<=-16'd6370;
      103398:data<=-16'd7891;
      103399:data<=-16'd8570;
      103400:data<=-16'd7823;
      103401:data<=-16'd7956;
      103402:data<=-16'd7705;
      103403:data<=-16'd7556;
      103404:data<=-16'd9438;
      103405:data<=-16'd10675;
      103406:data<=-16'd10151;
      103407:data<=-16'd9498;
      103408:data<=-16'd8994;
      103409:data<=-16'd8963;
      103410:data<=-16'd9488;
      103411:data<=-16'd10381;
      103412:data<=-16'd11151;
      103413:data<=-16'd10727;
      103414:data<=-16'd10220;
      103415:data<=-16'd10251;
      103416:data<=-16'd9714;
      103417:data<=-16'd10211;
      103418:data<=-16'd11835;
      103419:data<=-16'd11637;
      103420:data<=-16'd10598;
      103421:data<=-16'd10392;
      103422:data<=-16'd9878;
      103423:data<=-16'd10179;
      103424:data<=-16'd11756;
      103425:data<=-16'd11520;
      103426:data<=-16'd10151;
      103427:data<=-16'd10501;
      103428:data<=-16'd10492;
      103429:data<=-16'd9514;
      103430:data<=-16'd10152;
      103431:data<=-16'd9461;
      103432:data<=-16'd5612;
      103433:data<=-16'd3789;
      103434:data<=-16'd4381;
      103435:data<=-16'd3838;
      103436:data<=-16'd3607;
      103437:data<=-16'd4731;
      103438:data<=-16'd5679;
      103439:data<=-16'd5850;
      103440:data<=-16'd5245;
      103441:data<=-16'd4886;
      103442:data<=-16'd4833;
      103443:data<=-16'd4872;
      103444:data<=-16'd6305;
      103445:data<=-16'd7185;
      103446:data<=-16'd6273;
      103447:data<=-16'd6536;
      103448:data<=-16'd6760;
      103449:data<=-16'd5416;
      103450:data<=-16'd5821;
      103451:data<=-16'd7635;
      103452:data<=-16'd7984;
      103453:data<=-16'd7054;
      103454:data<=-16'd6161;
      103455:data<=-16'd6061;
      103456:data<=-16'd5124;
      103457:data<=-16'd3054;
      103458:data<=-16'd2934;
      103459:data<=-16'd3524;
      103460:data<=-16'd2435;
      103461:data<=-16'd1868;
      103462:data<=-16'd1939;
      103463:data<=-16'd2085;
      103464:data<=-16'd3803;
      103465:data<=-16'd4619;
      103466:data<=-16'd3224;
      103467:data<=-16'd3131;
      103468:data<=-16'd3523;
      103469:data<=-16'd2453;
      103470:data<=-16'd3116;
      103471:data<=-16'd5106;
      103472:data<=-16'd4937;
      103473:data<=-16'd4114;
      103474:data<=-16'd3762;
      103475:data<=-16'd3768;
      103476:data<=-16'd6849;
      103477:data<=-16'd11095;
      103478:data<=-16'd11790;
      103479:data<=-16'd10860;
      103480:data<=-16'd10681;
      103481:data<=-16'd10006;
      103482:data<=-16'd9365;
      103483:data<=-16'd9749;
      103484:data<=-16'd10434;
      103485:data<=-16'd10505;
      103486:data<=-16'd9818;
      103487:data<=-16'd9338;
      103488:data<=-16'd9107;
      103489:data<=-16'd8467;
      103490:data<=-16'd8407;
      103491:data<=-16'd9091;
      103492:data<=-16'd8969;
      103493:data<=-16'd8117;
      103494:data<=-16'd7674;
      103495:data<=-16'd7504;
      103496:data<=-16'd7077;
      103497:data<=-16'd6323;
      103498:data<=-16'd5395;
      103499:data<=-16'd4890;
      103500:data<=-16'd4792;
      103501:data<=-16'd4437;
      103502:data<=-16'd3985;
      103503:data<=-16'd2975;
      103504:data<=-16'd1251;
      103505:data<=-16'd617;
      103506:data<=-16'd679;
      103507:data<=16'd27;
      103508:data<=16'd356;
      103509:data<=16'd338;
      103510:data<=16'd1268;
      103511:data<=16'd2795;
      103512:data<=16'd3626;
      103513:data<=16'd3128;
      103514:data<=16'd3072;
      103515:data<=16'd3711;
      103516:data<=16'd3773;
      103517:data<=16'd5383;
      103518:data<=16'd6840;
      103519:data<=16'd5345;
      103520:data<=16'd6599;
      103521:data<=16'd11162;
      103522:data<=16'd12533;
      103523:data<=16'd11291;
      103524:data<=16'd9806;
      103525:data<=16'd8757;
      103526:data<=16'd9274;
      103527:data<=16'd9336;
      103528:data<=16'd8404;
      103529:data<=16'd8346;
      103530:data<=16'd9344;
      103531:data<=16'd10727;
      103532:data<=16'd10569;
      103533:data<=16'd9544;
      103534:data<=16'd9626;
      103535:data<=16'd9071;
      103536:data<=16'd8872;
      103537:data<=16'd10352;
      103538:data<=16'd10687;
      103539:data<=16'd10182;
      103540:data<=16'd9976;
      103541:data<=16'd9732;
      103542:data<=16'd9753;
      103543:data<=16'd9332;
      103544:data<=16'd10131;
      103545:data<=16'd11806;
      103546:data<=16'd10733;
      103547:data<=16'd9611;
      103548:data<=16'd9752;
      103549:data<=16'd9209;
      103550:data<=16'd10857;
      103551:data<=16'd12875;
      103552:data<=16'd11696;
      103553:data<=16'd10580;
      103554:data<=16'd10363;
      103555:data<=16'd10194;
      103556:data<=16'd10783;
      103557:data<=16'd11394;
      103558:data<=16'd11808;
      103559:data<=16'd11142;
      103560:data<=16'd10248;
      103561:data<=16'd10555;
      103562:data<=16'd9467;
      103563:data<=16'd9313;
      103564:data<=16'd11600;
      103565:data<=16'd9209;
      103566:data<=16'd3943;
      103567:data<=16'd2910;
      103568:data<=16'd3243;
      103569:data<=16'd2867;
      103570:data<=16'd3761;
      103571:data<=16'd4578;
      103572:data<=16'd4205;
      103573:data<=16'd4043;
      103574:data<=16'd4441;
      103575:data<=16'd3809;
      103576:data<=16'd3283;
      103577:data<=16'd4772;
      103578:data<=16'd5298;
      103579:data<=16'd4490;
      103580:data<=16'd5046;
      103581:data<=16'd5009;
      103582:data<=16'd4155;
      103583:data<=16'd4790;
      103584:data<=16'd5827;
      103585:data<=16'd6150;
      103586:data<=16'd5759;
      103587:data<=16'd5506;
      103588:data<=16'd5623;
      103589:data<=16'd5150;
      103590:data<=16'd6777;
      103591:data<=16'd10383;
      103592:data<=16'd11103;
      103593:data<=16'd10323;
      103594:data<=16'd9953;
      103595:data<=16'd8560;
      103596:data<=16'd8508;
      103597:data<=16'd9784;
      103598:data<=16'd9568;
      103599:data<=16'd8875;
      103600:data<=16'd8454;
      103601:data<=16'd7999;
      103602:data<=16'd7736;
      103603:data<=16'd7501;
      103604:data<=16'd7239;
      103605:data<=16'd6361;
      103606:data<=16'd5814;
      103607:data<=16'd6100;
      103608:data<=16'd5236;
      103609:data<=16'd5407;
      103610:data<=16'd7949;
      103611:data<=16'd8733;
      103612:data<=16'd8191;
      103613:data<=16'd8043;
      103614:data<=16'd6848;
      103615:data<=16'd6241;
      103616:data<=16'd5914;
      103617:data<=16'd3604;
      103618:data<=16'd2026;
      103619:data<=16'd2256;
      103620:data<=16'd2050;
      103621:data<=16'd1747;
      103622:data<=16'd1756;
      103623:data<=16'd657;
      103624:data<=-16'd1547;
      103625:data<=-16'd2541;
      103626:data<=-16'd1947;
      103627:data<=-16'd1970;
      103628:data<=-16'd2243;
      103629:data<=-16'd2579;
      103630:data<=-16'd4329;
      103631:data<=-16'd5034;
      103632:data<=-16'd4212;
      103633:data<=-16'd4780;
      103634:data<=-16'd5160;
      103635:data<=-16'd4701;
      103636:data<=-16'd5714;
      103637:data<=-16'd6921;
      103638:data<=-16'd7118;
      103639:data<=-16'd6998;
      103640:data<=-16'd6611;
      103641:data<=-16'd6472;
      103642:data<=-16'd6842;
      103643:data<=-16'd7785;
      103644:data<=-16'd8634;
      103645:data<=-16'd8244;
      103646:data<=-16'd8053;
      103647:data<=-16'd8440;
      103648:data<=-16'd8381;
      103649:data<=-16'd9016;
      103650:data<=-16'd9817;
      103651:data<=-16'd10011;
      103652:data<=-16'd9781;
      103653:data<=-16'd8836;
      103654:data<=-16'd10913;
      103655:data<=-16'd15282;
      103656:data<=-16'd15981;
      103657:data<=-16'd17344;
      103658:data<=-16'd21488;
      103659:data<=-16'd21372;
      103660:data<=-16'd19426;
      103661:data<=-16'd19456;
      103662:data<=-16'd18753;
      103663:data<=-16'd18980;
      103664:data<=-16'd19758;
      103665:data<=-16'd18531;
      103666:data<=-16'd17987;
      103667:data<=-16'd18019;
      103668:data<=-16'd16839;
      103669:data<=-16'd16230;
      103670:data<=-16'd16739;
      103671:data<=-16'd17108;
      103672:data<=-16'd16431;
      103673:data<=-16'd15637;
      103674:data<=-16'd15341;
      103675:data<=-16'd14164;
      103676:data<=-16'd13987;
      103677:data<=-16'd15531;
      103678:data<=-16'd14951;
      103679:data<=-16'd13436;
      103680:data<=-16'd13388;
      103681:data<=-16'd12674;
      103682:data<=-16'd12093;
      103683:data<=-16'd12871;
      103684:data<=-16'd12816;
      103685:data<=-16'd11949;
      103686:data<=-16'd11586;
      103687:data<=-16'd11201;
      103688:data<=-16'd10583;
      103689:data<=-16'd10640;
      103690:data<=-16'd11441;
      103691:data<=-16'd11635;
      103692:data<=-16'd10819;
      103693:data<=-16'd10164;
      103694:data<=-16'd9955;
      103695:data<=-16'd9371;
      103696:data<=-16'd9276;
      103697:data<=-16'd10640;
      103698:data<=-16'd9949;
      103699:data<=-16'd5374;
      103700:data<=-16'd2055;
      103701:data<=-16'd1820;
      103702:data<=-16'd2011;
      103703:data<=-16'd2884;
      103704:data<=-16'd3485;
      103705:data<=-16'd2843;
      103706:data<=-16'd3118;
      103707:data<=-16'd3319;
      103708:data<=-16'd2332;
      103709:data<=-16'd2097;
      103710:data<=-16'd2079;
      103711:data<=-16'd1512;
      103712:data<=-16'd1243;
      103713:data<=-16'd963;
      103714:data<=-16'd975;
      103715:data<=-16'd1093;
      103716:data<=16'd372;
      103717:data<=16'd2259;
      103718:data<=16'd2434;
      103719:data<=16'd2224;
      103720:data<=16'd2689;
      103721:data<=16'd2778;
      103722:data<=16'd2925;
      103723:data<=16'd3977;
      103724:data<=16'd6014;
      103725:data<=16'd8669;
      103726:data<=16'd9541;
      103727:data<=16'd8705;
      103728:data<=16'd9069;
      103729:data<=16'd9847;
      103730:data<=16'd10390;
      103731:data<=16'd10951;
      103732:data<=16'd10100;
      103733:data<=16'd10013;
      103734:data<=16'd10790;
      103735:data<=16'd9693;
      103736:data<=16'd10076;
      103737:data<=16'd11797;
      103738:data<=16'd11264;
      103739:data<=16'd11036;
      103740:data<=16'd10780;
      103741:data<=16'd9881;
      103742:data<=16'd10981;
      103743:data<=16'd9896;
      103744:data<=16'd5642;
      103745:data<=16'd4059;
      103746:data<=16'd4488;
      103747:data<=16'd4585;
      103748:data<=16'd4849;
      103749:data<=16'd4951;
      103750:data<=16'd5303;
      103751:data<=16'd5776;
      103752:data<=16'd6028;
      103753:data<=16'd6075;
      103754:data<=16'd5404;
      103755:data<=16'd5454;
      103756:data<=16'd6570;
      103757:data<=16'd7074;
      103758:data<=16'd7069;
      103759:data<=16'd6857;
      103760:data<=16'd6775;
      103761:data<=16'd6751;
      103762:data<=16'd6660;
      103763:data<=16'd7990;
      103764:data<=16'd8825;
      103765:data<=16'd7559;
      103766:data<=16'd7432;
      103767:data<=16'd7847;
      103768:data<=16'd7166;
      103769:data<=16'd7644;
      103770:data<=16'd8827;
      103771:data<=16'd8992;
      103772:data<=16'd8326;
      103773:data<=16'd7658;
      103774:data<=16'd7445;
      103775:data<=16'd7171;
      103776:data<=16'd8100;
      103777:data<=16'd9207;
      103778:data<=16'd7649;
      103779:data<=16'd7003;
      103780:data<=16'd7720;
      103781:data<=16'd6464;
      103782:data<=16'd6799;
      103783:data<=16'd8325;
      103784:data<=16'd7636;
      103785:data<=16'd7588;
      103786:data<=16'd7511;
      103787:data<=16'd6796;
      103788:data<=16'd9077;
      103789:data<=16'd12860;
      103790:data<=16'd14819;
      103791:data<=16'd12965;
      103792:data<=16'd8704;
      103793:data<=16'd7503;
      103794:data<=16'd8003;
      103795:data<=16'd7394;
      103796:data<=16'd8211;
      103797:data<=16'd8760;
      103798:data<=16'd7978;
      103799:data<=16'd8170;
      103800:data<=16'd7806;
      103801:data<=16'd7013;
      103802:data<=16'd7467;
      103803:data<=16'd8109;
      103804:data<=16'd8322;
      103805:data<=16'd7724;
      103806:data<=16'd7071;
      103807:data<=16'd6865;
      103808:data<=16'd6112;
      103809:data<=16'd6520;
      103810:data<=16'd7777;
      103811:data<=16'd7162;
      103812:data<=16'd6214;
      103813:data<=16'd5917;
      103814:data<=16'd5551;
      103815:data<=16'd5374;
      103816:data<=16'd4695;
      103817:data<=16'd4494;
      103818:data<=16'd5053;
      103819:data<=16'd4498;
      103820:data<=16'd3970;
      103821:data<=16'd3635;
      103822:data<=16'd2009;
      103823:data<=16'd438;
      103824:data<=-16'd126;
      103825:data<=-16'd174;
      103826:data<=-16'd769;
      103827:data<=-16'd1504;
      103828:data<=-16'd870;
      103829:data<=-16'd1889;
      103830:data<=-16'd4272;
      103831:data<=-16'd3479;
      103832:data<=-16'd4293;
      103833:data<=-16'd9051;
      103834:data<=-16'd10859;
      103835:data<=-16'd10710;
      103836:data<=-16'd11834;
      103837:data<=-16'd11822;
      103838:data<=-16'd11532;
      103839:data<=-16'd11806;
      103840:data<=-16'd11373;
      103841:data<=-16'd11063;
      103842:data<=-16'd11480;
      103843:data<=-16'd12375;
      103844:data<=-16'd12452;
      103845:data<=-16'd11620;
      103846:data<=-16'd11808;
      103847:data<=-16'd11564;
      103848:data<=-16'd10640;
      103849:data<=-16'd11523;
      103850:data<=-16'd12231;
      103851:data<=-16'd11721;
      103852:data<=-16'd11550;
      103853:data<=-16'd11183;
      103854:data<=-16'd11115;
      103855:data<=-16'd11323;
      103856:data<=-16'd11520;
      103857:data<=-16'd12257;
      103858:data<=-16'd10662;
      103859:data<=-16'd7498;
      103860:data<=-16'd6893;
      103861:data<=-16'd6848;
      103862:data<=-16'd6710;
      103863:data<=-16'd8066;
      103864:data<=-16'd8523;
      103865:data<=-16'd7993;
      103866:data<=-16'd7680;
      103867:data<=-16'd6995;
      103868:data<=-16'd6912;
      103869:data<=-16'd7962;
      103870:data<=-16'd9251;
      103871:data<=-16'd9021;
      103872:data<=-16'd7662;
      103873:data<=-16'd8009;
      103874:data<=-16'd7918;
      103875:data<=-16'd7174;
      103876:data<=-16'd9135;
      103877:data<=-16'd7920;
      103878:data<=-16'd2334;
      103879:data<=-16'd1139;
      103880:data<=-16'd2185;
      103881:data<=-16'd1166;
      103882:data<=-16'd1859;
      103883:data<=-16'd3463;
      103884:data<=-16'd3695;
      103885:data<=-16'd3707;
      103886:data<=-16'd3482;
      103887:data<=-16'd3036;
      103888:data<=-16'd2945;
      103889:data<=-16'd3744;
      103890:data<=-16'd4410;
      103891:data<=-16'd3758;
      103892:data<=-16'd3959;
      103893:data<=-16'd4369;
      103894:data<=-16'd3069;
      103895:data<=-16'd3204;
      103896:data<=-16'd4840;
      103897:data<=-16'd5128;
      103898:data<=-16'd4851;
      103899:data<=-16'd4602;
      103900:data<=-16'd4185;
      103901:data<=-16'd3762;
      103902:data<=-16'd3983;
      103903:data<=-16'd5351;
      103904:data<=-16'd5523;
      103905:data<=-16'd4679;
      103906:data<=-16'd5049;
      103907:data<=-16'd4634;
      103908:data<=-16'd4006;
      103909:data<=-16'd5207;
      103910:data<=-16'd5659;
      103911:data<=-16'd5269;
      103912:data<=-16'd5433;
      103913:data<=-16'd4822;
      103914:data<=-16'd3959;
      103915:data<=-16'd4317;
      103916:data<=-16'd5486;
      103917:data<=-16'd6008;
      103918:data<=-16'd5677;
      103919:data<=-16'd5422;
      103920:data<=-16'd4569;
      103921:data<=-16'd4948;
      103922:data<=-16'd8575;
      103923:data<=-16'd10642;
      103924:data<=-16'd9940;
      103925:data<=-16'd10969;
      103926:data<=-16'd12615;
      103927:data<=-16'd12712;
      103928:data<=-16'd11614;
      103929:data<=-16'd9110;
      103930:data<=-16'd7518;
      103931:data<=-16'd7830;
      103932:data<=-16'd7303;
      103933:data<=-16'd6258;
      103934:data<=-16'd6243;
      103935:data<=-16'd5377;
      103936:data<=-16'd3090;
      103937:data<=-16'd2100;
      103938:data<=-16'd2319;
      103939:data<=-16'd1478;
      103940:data<=-16'd926;
      103941:data<=-16'd1209;
      103942:data<=-16'd30;
      103943:data<=16'd1612;
      103944:data<=16'd2043;
      103945:data<=16'd2162;
      103946:data<=16'd2303;
      103947:data<=16'd2464;
      103948:data<=16'd3083;
      103949:data<=16'd4417;
      103950:data<=16'd5632;
      103951:data<=16'd5723;
      103952:data<=16'd5888;
      103953:data<=16'd5956;
      103954:data<=16'd5215;
      103955:data<=16'd6108;
      103956:data<=16'd7567;
      103957:data<=16'd7071;
      103958:data<=16'd6980;
      103959:data<=16'd7574;
      103960:data<=16'd7441;
      103961:data<=16'd7582;
      103962:data<=16'd8199;
      103963:data<=16'd9470;
      103964:data<=16'd9946;
      103965:data<=16'd8772;
      103966:data<=16'd10426;
      103967:data<=16'd14366;
      103968:data<=16'd15499;
      103969:data<=16'd15760;
      103970:data<=16'd16606;
      103971:data<=16'd15885;
      103972:data<=16'd15227;
      103973:data<=16'd15065;
      103974:data<=16'd13916;
      103975:data<=16'd13976;
      103976:data<=16'd15670;
      103977:data<=16'd15820;
      103978:data<=16'd14794;
      103979:data<=16'd14710;
      103980:data<=16'd14440;
      103981:data<=16'd13855;
      103982:data<=16'd14501;
      103983:data<=16'd14998;
      103984:data<=16'd14336;
      103985:data<=16'd13896;
      103986:data<=16'd13702;
      103987:data<=16'd13229;
      103988:data<=16'd13007;
      103989:data<=16'd13541;
      103990:data<=16'd13867;
      103991:data<=16'd13106;
      103992:data<=16'd13784;
      103993:data<=16'd15894;
      103994:data<=16'd15670;
      103995:data<=16'd15242;
      103996:data<=16'd16530;
      103997:data<=16'd15957;
      103998:data<=16'd14621;
      103999:data<=16'd14393;
      104000:data<=16'd13573;
      104001:data<=16'd13514;
      104002:data<=16'd14305;
      104003:data<=16'd13975;
      104004:data<=16'd13441;
      104005:data<=16'd12771;
      104006:data<=16'd11771;
      104007:data<=16'd11147;
      104008:data<=16'd11056;
      104009:data<=16'd12351;
      104010:data<=16'd12287;
      104011:data<=16'd8155;
      104012:data<=16'd4652;
      104013:data<=16'd3929;
      104014:data<=16'd3251;
      104015:data<=16'd3571;
      104016:data<=16'd4849;
      104017:data<=16'd4598;
      104018:data<=16'd3845;
      104019:data<=16'd3859;
      104020:data<=16'd3621;
      104021:data<=16'd3457;
      104022:data<=16'd4375;
      104023:data<=16'd5059;
      104024:data<=16'd4679;
      104025:data<=16'd4636;
      104026:data<=16'd4463;
      104027:data<=16'd3654;
      104028:data<=16'd3688;
      104029:data<=16'd3539;
      104030:data<=16'd2696;
      104031:data<=16'd2645;
      104032:data<=16'd2161;
      104033:data<=16'd1474;
      104034:data<=16'd1807;
      104035:data<=16'd784;
      104036:data<=-16'd1124;
      104037:data<=-16'd1343;
      104038:data<=-16'd1224;
      104039:data<=-16'd1597;
      104040:data<=-16'd1612;
      104041:data<=-16'd1939;
      104042:data<=-16'd3237;
      104043:data<=-16'd4316;
      104044:data<=-16'd4105;
      104045:data<=-16'd4079;
      104046:data<=-16'd4532;
      104047:data<=-16'd4153;
      104048:data<=-16'd4711;
      104049:data<=-16'd6094;
      104050:data<=-16'd6038;
      104051:data<=-16'd5971;
      104052:data<=-16'd5906;
      104053:data<=-16'd5544;
      104054:data<=-16'd6543;
      104055:data<=-16'd5877;
      104056:data<=-16'd2705;
      104057:data<=-16'd1143;
      104058:data<=-16'd1348;
      104059:data<=-16'd3057;
      104060:data<=-16'd5521;
      104061:data<=-16'd6097;
      104062:data<=-16'd6804;
      104063:data<=-16'd8019;
      104064:data<=-16'd7460;
      104065:data<=-16'd7330;
      104066:data<=-16'd7515;
      104067:data<=-16'd6711;
      104068:data<=-16'd7363;
      104069:data<=-16'd8669;
      104070:data<=-16'd8621;
      104071:data<=-16'd8185;
      104072:data<=-16'd7990;
      104073:data<=-16'd7856;
      104074:data<=-16'd7618;
      104075:data<=-16'd8478;
      104076:data<=-16'd9931;
      104077:data<=-16'd9150;
      104078:data<=-16'd8258;
      104079:data<=-16'd8690;
      104080:data<=-16'd7885;
      104081:data<=-16'd8047;
      104082:data<=-16'd9829;
      104083:data<=-16'd9914;
      104084:data<=-16'd9415;
      104085:data<=-16'd9216;
      104086:data<=-16'd8636;
      104087:data<=-16'd8621;
      104088:data<=-16'd9317;
      104089:data<=-16'd10571;
      104090:data<=-16'd10680;
      104091:data<=-16'd9394;
      104092:data<=-16'd9417;
      104093:data<=-16'd9259;
      104094:data<=-16'd8931;
      104095:data<=-16'd10622;
      104096:data<=-16'd10895;
      104097:data<=-16'd9938;
      104098:data<=-16'd9903;
      104099:data<=-16'd8866;
      104100:data<=-16'd10255;
      104101:data<=-16'd14806;
      104102:data<=-16'd16569;
      104103:data<=-16'd16105;
      104104:data<=-16'd15547;
      104105:data<=-16'd14739;
      104106:data<=-16'd14389;
      104107:data<=-16'd13261;
      104108:data<=-16'd12842;
      104109:data<=-16'd14302;
      104110:data<=-16'd14007;
      104111:data<=-16'd12739;
      104112:data<=-16'd12552;
      104113:data<=-16'd11882;
      104114:data<=-16'd11527;
      104115:data<=-16'd12232;
      104116:data<=-16'd12700;
      104117:data<=-16'd12339;
      104118:data<=-16'd11430;
      104119:data<=-16'd10859;
      104120:data<=-16'd10345;
      104121:data<=-16'd10249;
      104122:data<=-16'd11192;
      104123:data<=-16'd11059;
      104124:data<=-16'd10343;
      104125:data<=-16'd10070;
      104126:data<=-16'd7482;
      104127:data<=-16'd4252;
      104128:data<=-16'd4126;
      104129:data<=-16'd5168;
      104130:data<=-16'd5080;
      104131:data<=-16'd4555;
      104132:data<=-16'd4555;
      104133:data<=-16'd4525;
      104134:data<=-16'd3783;
      104135:data<=-16'd3316;
      104136:data<=-16'd3310;
      104137:data<=-16'd3216;
      104138:data<=-16'd2814;
      104139:data<=-16'd2111;
      104140:data<=-16'd2224;
      104141:data<=-16'd1425;
      104142:data<=16'd1105;
      104143:data<=16'd1356;
      104144:data<=16'd2064;
      104145:data<=16'd6631;
      104146:data<=16'd8601;
      104147:data<=16'd7497;
      104148:data<=16'd8466;
      104149:data<=16'd9643;
      104150:data<=16'd9691;
      104151:data<=16'd9636;
      104152:data<=16'd9072;
      104153:data<=16'd8780;
      104154:data<=16'd9144;
      104155:data<=16'd10056;
      104156:data<=16'd10684;
      104157:data<=16'd9988;
      104158:data<=16'd9856;
      104159:data<=16'd10210;
      104160:data<=16'd9517;
      104161:data<=16'd9726;
      104162:data<=16'd10875;
      104163:data<=16'd11227;
      104164:data<=16'd11024;
      104165:data<=16'd10455;
      104166:data<=16'd9961;
      104167:data<=16'd9729;
      104168:data<=16'd10146;
      104169:data<=16'd11449;
      104170:data<=16'd11356;
      104171:data<=16'd10440;
      104172:data<=16'd10568;
      104173:data<=16'd9884;
      104174:data<=16'd9511;
      104175:data<=16'd10615;
      104176:data<=16'd10511;
      104177:data<=16'd9932;
      104178:data<=16'd9849;
      104179:data<=16'd9280;
      104180:data<=16'd8969;
      104181:data<=16'd9077;
      104182:data<=16'd9950;
      104183:data<=16'd10351;
      104184:data<=16'd8907;
      104185:data<=16'd8869;
      104186:data<=16'd8942;
      104187:data<=16'd7659;
      104188:data<=16'd9646;
      104189:data<=16'd9561;
      104190:data<=16'd3714;
      104191:data<=16'd2115;
      104192:data<=16'd3192;
      104193:data<=-16'd94;
      104194:data<=-16'd1735;
      104195:data<=-16'd123;
      104196:data<=16'd293;
      104197:data<=16'd168;
      104198:data<=16'd49;
      104199:data<=-16'd18;
      104200:data<=16'd132;
      104201:data<=16'd265;
      104202:data<=16'd1421;
      104203:data<=16'd1979;
      104204:data<=16'd1081;
      104205:data<=16'd1152;
      104206:data<=16'd1442;
      104207:data<=16'd1456;
      104208:data<=16'd2567;
      104209:data<=16'd3130;
      104210:data<=16'd2692;
      104211:data<=16'd2678;
      104212:data<=16'd2366;
      104213:data<=16'd1733;
      104214:data<=16'd2152;
      104215:data<=16'd3462;
      104216:data<=16'd4252;
      104217:data<=16'd4055;
      104218:data<=16'd3774;
      104219:data<=16'd3579;
      104220:data<=16'd3253;
      104221:data<=16'd3858;
      104222:data<=16'd5288;
      104223:data<=16'd5450;
      104224:data<=16'd4423;
      104225:data<=16'd4134;
      104226:data<=16'd4020;
      104227:data<=16'd3689;
      104228:data<=16'd4684;
      104229:data<=16'd5523;
      104230:data<=16'd5057;
      104231:data<=16'd5190;
      104232:data<=16'd4808;
      104233:data<=16'd4541;
      104234:data<=16'd8208;
      104235:data<=16'd12261;
      104236:data<=16'd12373;
      104237:data<=16'd11377;
      104238:data<=16'd10671;
      104239:data<=16'd9875;
      104240:data<=16'd9720;
      104241:data<=16'd9062;
      104242:data<=16'd7950;
      104243:data<=16'd7626;
      104244:data<=16'd7210;
      104245:data<=16'd6757;
      104246:data<=16'd6813;
      104247:data<=16'd5985;
      104248:data<=16'd4188;
      104249:data<=16'd3153;
      104250:data<=16'd2889;
      104251:data<=16'd2278;
      104252:data<=16'd1812;
      104253:data<=16'd2082;
      104254:data<=16'd1671;
      104255:data<=16'd14;
      104256:data<=-16'd901;
      104257:data<=-16'd678;
      104258:data<=-16'd1104;
      104259:data<=-16'd952;
      104260:data<=16'd1227;
      104261:data<=16'd1858;
      104262:data<=16'd18;
      104263:data<=-16'd422;
      104264:data<=-16'd161;
      104265:data<=-16'd839;
      104266:data<=-16'd754;
      104267:data<=-16'd1239;
      104268:data<=-16'd3069;
      104269:data<=-16'd3559;
      104270:data<=-16'd3048;
      104271:data<=-16'd3274;
      104272:data<=-16'd3930;
      104273:data<=-16'd4168;
      104274:data<=-16'd4414;
      104275:data<=-16'd6266;
      104276:data<=-16'd7269;
      104277:data<=-16'd5638;
      104278:data<=-16'd7016;
      104279:data<=-16'd11430;
      104280:data<=-16'd12834;
      104281:data<=-16'd13145;
      104282:data<=-16'd14272;
      104283:data<=-16'd13759;
      104284:data<=-16'd13314;
      104285:data<=-16'd13511;
      104286:data<=-16'd12794;
      104287:data<=-16'd12775;
      104288:data<=-16'd13473;
      104289:data<=-16'd13414;
      104290:data<=-16'd13147;
      104291:data<=-16'd13066;
      104292:data<=-16'd12784;
      104293:data<=-16'd12057;
      104294:data<=-16'd12158;
      104295:data<=-16'd13659;
      104296:data<=-16'd13747;
      104297:data<=-16'd12372;
      104298:data<=-16'd12367;
      104299:data<=-16'd12571;
      104300:data<=-16'd11975;
      104301:data<=-16'd12610;
      104302:data<=-16'd13629;
      104303:data<=-16'd12766;
      104304:data<=-16'd11535;
      104305:data<=-16'd11544;
      104306:data<=-16'd11028;
      104307:data<=-16'd10292;
      104308:data<=-16'd11294;
      104309:data<=-16'd11626;
      104310:data<=-16'd10246;
      104311:data<=-16'd9908;
      104312:data<=-16'd9864;
      104313:data<=-16'd9030;
      104314:data<=-16'd9194;
      104315:data<=-16'd10275;
      104316:data<=-16'd10631;
      104317:data<=-16'd9529;
      104318:data<=-16'd8505;
      104319:data<=-16'd8563;
      104320:data<=-16'd7926;
      104321:data<=-16'd8017;
      104322:data<=-16'd9194;
      104323:data<=-16'd6633;
      104324:data<=-16'd2359;
      104325:data<=-16'd1292;
      104326:data<=-16'd1835;
      104327:data<=-16'd3944;
      104328:data<=-16'd6983;
      104329:data<=-16'd7215;
      104330:data<=-16'd6232;
      104331:data<=-16'd6187;
      104332:data<=-16'd5799;
      104333:data<=-16'd5450;
      104334:data<=-16'd5805;
      104335:data<=-16'd6370;
      104336:data<=-16'd6223;
      104337:data<=-16'd5456;
      104338:data<=-16'd5510;
      104339:data<=-16'd5412;
      104340:data<=-16'd4717;
      104341:data<=-16'd5275;
      104342:data<=-16'd5870;
      104343:data<=-16'd5386;
      104344:data<=-16'd4945;
      104345:data<=-16'd4400;
      104346:data<=-16'd4065;
      104347:data<=-16'd3891;
      104348:data<=-16'd3204;
      104349:data<=-16'd3110;
      104350:data<=-16'd3153;
      104351:data<=-16'd2352;
      104352:data<=-16'd2138;
      104353:data<=-16'd2344;
      104354:data<=-16'd1350;
      104355:data<=16'd299;
      104356:data<=16'd923;
      104357:data<=16'd661;
      104358:data<=16'd837;
      104359:data<=16'd1052;
      104360:data<=16'd1353;
      104361:data<=16'd2784;
      104362:data<=16'd3814;
      104363:data<=16'd3519;
      104364:data<=16'd3213;
      104365:data<=16'd3868;
      104366:data<=16'd5559;
      104367:data<=16'd5262;
      104368:data<=16'd2285;
      104369:data<=16'd1293;
      104370:data<=16'd1955;
      104371:data<=16'd1638;
      104372:data<=16'd1572;
      104373:data<=16'd1400;
      104374:data<=16'd2073;
      104375:data<=16'd4299;
      104376:data<=16'd4579;
      104377:data<=16'd4079;
      104378:data<=16'd4678;
      104379:data<=16'd4285;
      104380:data<=16'd4642;
      104381:data<=16'd6169;
      104382:data<=16'd6334;
      104383:data<=16'd6128;
      104384:data<=16'd6072;
      104385:data<=16'd6003;
      104386:data<=16'd6184;
      104387:data<=16'd6267;
      104388:data<=16'd7359;
      104389:data<=16'd8025;
      104390:data<=16'd7177;
      104391:data<=16'd7423;
      104392:data<=16'd7518;
      104393:data<=16'd7507;
      104394:data<=16'd10084;
      104395:data<=16'd11677;
      104396:data<=16'd10847;
      104397:data<=16'd10769;
      104398:data<=16'd10944;
      104399:data<=16'd10778;
      104400:data<=16'd11148;
      104401:data<=16'd12051;
      104402:data<=16'd12524;
      104403:data<=16'd11800;
      104404:data<=16'd11527;
      104405:data<=16'd11388;
      104406:data<=16'd10530;
      104407:data<=16'd11257;
      104408:data<=16'd12372;
      104409:data<=16'd12443;
      104410:data<=16'd12067;
      104411:data<=16'd10517;
      104412:data<=16'd11973;
      104413:data<=16'd16756;
      104414:data<=16'd17899;
      104415:data<=16'd17182;
      104416:data<=16'd17399;
      104417:data<=16'd16465;
      104418:data<=16'd16184;
      104419:data<=16'd15685;
      104420:data<=16'd14425;
      104421:data<=16'd15396;
      104422:data<=16'd15791;
      104423:data<=16'd14598;
      104424:data<=16'd14402;
      104425:data<=16'd13668;
      104426:data<=16'd12636;
      104427:data<=16'd13077;
      104428:data<=16'd14152;
      104429:data<=16'd14251;
      104430:data<=16'd12760;
      104431:data<=16'd11953;
      104432:data<=16'd12187;
      104433:data<=16'd11897;
      104434:data<=16'd12369;
      104435:data<=16'd12648;
      104436:data<=16'd11691;
      104437:data<=16'd11297;
      104438:data<=16'd10580;
      104439:data<=16'd9456;
      104440:data<=16'd9512;
      104441:data<=16'd10369;
      104442:data<=16'd10906;
      104443:data<=16'd9679;
      104444:data<=16'd8340;
      104445:data<=16'd8361;
      104446:data<=16'd7592;
      104447:data<=16'd7823;
      104448:data<=16'd9442;
      104449:data<=16'd8789;
      104450:data<=16'd7674;
      104451:data<=16'd7594;
      104452:data<=16'd7259;
      104453:data<=16'd6792;
      104454:data<=16'd5573;
      104455:data<=16'd5277;
      104456:data<=16'd4902;
      104457:data<=16'd607;
      104458:data<=-16'd2649;
      104459:data<=-16'd2147;
      104460:data<=-16'd3378;
      104461:data<=-16'd6208;
      104462:data<=-16'd7644;
      104463:data<=-16'd7624;
      104464:data<=-16'd7050;
      104465:data<=-16'd6948;
      104466:data<=-16'd6646;
      104467:data<=-16'd7194;
      104468:data<=-16'd9086;
      104469:data<=-16'd9213;
      104470:data<=-16'd8589;
      104471:data<=-16'd8725;
      104472:data<=-16'd8188;
      104473:data<=-16'd8722;
      104474:data<=-16'd10316;
      104475:data<=-16'd10610;
      104476:data<=-16'd10273;
      104477:data<=-16'd9888;
      104478:data<=-16'd9667;
      104479:data<=-16'd9683;
      104480:data<=-16'd9755;
      104481:data<=-16'd10520;
      104482:data<=-16'd10716;
      104483:data<=-16'd10113;
      104484:data<=-16'd10108;
      104485:data<=-16'd9615;
      104486:data<=-16'd9468;
      104487:data<=-16'd10798;
      104488:data<=-16'd11210;
      104489:data<=-16'd10525;
      104490:data<=-16'd10100;
      104491:data<=-16'd9879;
      104492:data<=-16'd9694;
      104493:data<=-16'd9782;
      104494:data<=-16'd11088;
      104495:data<=-16'd11793;
      104496:data<=-16'd10530;
      104497:data<=-16'd10386;
      104498:data<=-16'd10390;
      104499:data<=-16'd9323;
      104500:data<=-16'd10305;
      104501:data<=-16'd9606;
      104502:data<=-16'd4902;
      104503:data<=-16'd3022;
      104504:data<=-16'd4081;
      104505:data<=-16'd3759;
      104506:data<=-16'd3859;
      104507:data<=-16'd5145;
      104508:data<=-16'd5762;
      104509:data<=-16'd5670;
      104510:data<=-16'd5653;
      104511:data<=-16'd5865;
      104512:data<=-16'd5468;
      104513:data<=-16'd5195;
      104514:data<=-16'd6355;
      104515:data<=-16'd7066;
      104516:data<=-16'd6440;
      104517:data<=-16'd6053;
      104518:data<=-16'd5648;
      104519:data<=-16'd5181;
      104520:data<=-16'd5981;
      104521:data<=-16'd7200;
      104522:data<=-16'd7285;
      104523:data<=-16'd6721;
      104524:data<=-16'd6166;
      104525:data<=-16'd5698;
      104526:data<=-16'd6029;
      104527:data<=-16'd6620;
      104528:data<=-16'd5852;
      104529:data<=-16'd4836;
      104530:data<=-16'd5007;
      104531:data<=-16'd4871;
      104532:data<=-16'd4068;
      104533:data<=-16'd4461;
      104534:data<=-16'd6120;
      104535:data<=-16'd6918;
      104536:data<=-16'd6058;
      104537:data<=-16'd5298;
      104538:data<=-16'd4989;
      104539:data<=-16'd4387;
      104540:data<=-16'd5195;
      104541:data<=-16'd6807;
      104542:data<=-16'd6634;
      104543:data<=-16'd6290;
      104544:data<=-16'd6247;
      104545:data<=-16'd5836;
      104546:data<=-16'd8622;
      104547:data<=-16'd13126;
      104548:data<=-16'd13675;
      104549:data<=-16'd12424;
      104550:data<=-16'd12455;
      104551:data<=-16'd11905;
      104552:data<=-16'd11025;
      104553:data<=-16'd11289;
      104554:data<=-16'd12098;
      104555:data<=-16'd12167;
      104556:data<=-16'd11044;
      104557:data<=-16'd10290;
      104558:data<=-16'd10426;
      104559:data<=-16'd9981;
      104560:data<=-16'd9094;
      104561:data<=-16'd8294;
      104562:data<=-16'd7608;
      104563:data<=-16'd7548;
      104564:data<=-16'd7524;
      104565:data<=-16'd6953;
      104566:data<=-16'd5993;
      104567:data<=-16'd4414;
      104568:data<=-16'd3206;
      104569:data<=-16'd3313;
      104570:data<=-16'd3491;
      104571:data<=-16'd3040;
      104572:data<=-16'd2537;
      104573:data<=-16'd1519;
      104574:data<=16'd82;
      104575:data<=16'd672;
      104576:data<=16'd588;
      104577:data<=16'd1368;
      104578:data<=16'd1636;
      104579:data<=16'd1336;
      104580:data<=16'd2585;
      104581:data<=16'd3915;
      104582:data<=16'd3792;
      104583:data<=16'd3600;
      104584:data<=16'd3785;
      104585:data<=16'd4009;
      104586:data<=16'd4470;
      104587:data<=16'd5865;
      104588:data<=16'd6755;
      104589:data<=16'd5577;
      104590:data<=16'd7156;
      104591:data<=16'd11916;
      104592:data<=16'd12787;
      104593:data<=16'd12179;
      104594:data<=16'd13314;
      104595:data<=16'd11947;
      104596:data<=16'd10709;
      104597:data<=16'd11439;
      104598:data<=16'd10422;
      104599:data<=16'd9993;
      104600:data<=16'd11229;
      104601:data<=16'd11691;
      104602:data<=16'd11552;
      104603:data<=16'd10687;
      104604:data<=16'd10466;
      104605:data<=16'd10831;
      104606:data<=16'd10137;
      104607:data<=16'd10945;
      104608:data<=16'd12000;
      104609:data<=16'd10845;
      104610:data<=16'd10836;
      104611:data<=16'd11201;
      104612:data<=16'd10252;
      104613:data<=16'd10753;
      104614:data<=16'd12051;
      104615:data<=16'd12176;
      104616:data<=16'd11441;
      104617:data<=16'd10677;
      104618:data<=16'd10198;
      104619:data<=16'd9717;
      104620:data<=16'd10596;
      104621:data<=16'd11565;
      104622:data<=16'd10102;
      104623:data<=16'd9339;
      104624:data<=16'd9734;
      104625:data<=16'd8945;
      104626:data<=16'd8969;
      104627:data<=16'd9756;
      104628:data<=16'd10025;
      104629:data<=16'd9823;
      104630:data<=16'd8809;
      104631:data<=16'd8396;
      104632:data<=16'd7703;
      104633:data<=16'd7306;
      104634:data<=16'd9514;
      104635:data<=16'd7961;
      104636:data<=16'd2284;
      104637:data<=16'd1177;
      104638:data<=16'd1968;
      104639:data<=16'd1259;
      104640:data<=16'd2306;
      104641:data<=16'd3049;
      104642:data<=16'd2570;
      104643:data<=16'd2736;
      104644:data<=16'd2573;
      104645:data<=16'd2244;
      104646:data<=16'd2388;
      104647:data<=16'd3369;
      104648:data<=16'd4328;
      104649:data<=16'd3381;
      104650:data<=16'd2626;
      104651:data<=16'd2796;
      104652:data<=16'd2165;
      104653:data<=16'd2763;
      104654:data<=16'd4356;
      104655:data<=16'd4200;
      104656:data<=16'd3351;
      104657:data<=16'd3204;
      104658:data<=16'd3469;
      104659:data<=16'd3651;
      104660:data<=16'd3982;
      104661:data<=16'd5112;
      104662:data<=16'd6191;
      104663:data<=16'd6602;
      104664:data<=16'd6278;
      104665:data<=16'd5325;
      104666:data<=16'd5159;
      104667:data<=16'd5253;
      104668:data<=16'd4610;
      104669:data<=16'd4205;
      104670:data<=16'd3718;
      104671:data<=16'd3377;
      104672:data<=16'd3378;
      104673:data<=16'd2085;
      104674:data<=16'd543;
      104675:data<=16'd49;
      104676:data<=16'd85;
      104677:data<=16'd415;
      104678:data<=-16'd174;
      104679:data<=-16'd144;
      104680:data<=16'd2282;
      104681:data<=16'd3556;
      104682:data<=16'd3027;
      104683:data<=16'd2874;
      104684:data<=16'd2457;
      104685:data<=16'd2194;
      104686:data<=16'd1568;
      104687:data<=-16'd224;
      104688:data<=-16'd907;
      104689:data<=-16'd1074;
      104690:data<=-16'd1668;
      104691:data<=-16'd1061;
      104692:data<=-16'd1048;
      104693:data<=-16'd2798;
      104694:data<=-16'd3880;
      104695:data<=-16'd3742;
      104696:data<=-16'd3560;
      104697:data<=-16'd3918;
      104698:data<=-16'd4355;
      104699:data<=-16'd4730;
      104700:data<=-16'd5639;
      104701:data<=-16'd5965;
      104702:data<=-16'd5767;
      104703:data<=-16'd6473;
      104704:data<=-16'd6537;
      104705:data<=-16'd5815;
      104706:data<=-16'd6492;
      104707:data<=-16'd7952;
      104708:data<=-16'd8740;
      104709:data<=-16'd8446;
      104710:data<=-16'd7771;
      104711:data<=-16'd7827;
      104712:data<=-16'd8169;
      104713:data<=-16'd9127;
      104714:data<=-16'd10337;
      104715:data<=-16'd9794;
      104716:data<=-16'd9053;
      104717:data<=-16'd9414;
      104718:data<=-16'd9385;
      104719:data<=-16'd9679;
      104720:data<=-16'd10710;
      104721:data<=-16'd11579;
      104722:data<=-16'd11603;
      104723:data<=-16'd10525;
      104724:data<=-16'd11690;
      104725:data<=-16'd15555;
      104726:data<=-16'd17130;
      104727:data<=-16'd16941;
      104728:data<=-16'd17656;
      104729:data<=-16'd17928;
      104730:data<=-16'd17716;
      104731:data<=-16'd17217;
      104732:data<=-16'd16540;
      104733:data<=-16'd16920;
      104734:data<=-16'd17071;
      104735:data<=-16'd16217;
      104736:data<=-16'd15711;
      104737:data<=-16'd15455;
      104738:data<=-16'd14977;
      104739:data<=-16'd14663;
      104740:data<=-16'd15164;
      104741:data<=-16'd15594;
      104742:data<=-16'd14299;
      104743:data<=-16'd12863;
      104744:data<=-16'd12401;
      104745:data<=-16'd11779;
      104746:data<=-16'd12091;
      104747:data<=-16'd13098;
      104748:data<=-16'd12657;
      104749:data<=-16'd11697;
      104750:data<=-16'd11159;
      104751:data<=-16'd10379;
      104752:data<=-16'd9919;
      104753:data<=-16'd10386;
      104754:data<=-16'd10768;
      104755:data<=-16'd10229;
      104756:data<=-16'd9635;
      104757:data<=-16'd9127;
      104758:data<=-16'd8187;
      104759:data<=-16'd8103;
      104760:data<=-16'd8983;
      104761:data<=-16'd9307;
      104762:data<=-16'd8771;
      104763:data<=-16'd7718;
      104764:data<=-16'd7039;
      104765:data<=-16'd6680;
      104766:data<=-16'd6593;
      104767:data<=-16'd7777;
      104768:data<=-16'd6996;
      104769:data<=-16'd2441;
      104770:data<=16'd625;
      104771:data<=16'd901;
      104772:data<=16'd1233;
      104773:data<=16'd1378;
      104774:data<=16'd1345;
      104775:data<=16'd1533;
      104776:data<=16'd1949;
      104777:data<=16'd2590;
      104778:data<=16'd2596;
      104779:data<=16'd3218;
      104780:data<=16'd4851;
      104781:data<=16'd5257;
      104782:data<=16'd5197;
      104783:data<=16'd5639;
      104784:data<=16'd5503;
      104785:data<=16'd5409;
      104786:data<=16'd6363;
      104787:data<=16'd7586;
      104788:data<=16'd7624;
      104789:data<=16'd7544;
      104790:data<=16'd8476;
      104791:data<=16'd8237;
      104792:data<=16'd8254;
      104793:data<=16'd10111;
      104794:data<=16'd10081;
      104795:data<=16'd9815;
      104796:data<=16'd11671;
      104797:data<=16'd11802;
      104798:data<=16'd11113;
      104799:data<=16'd11876;
      104800:data<=16'd12666;
      104801:data<=16'd13333;
      104802:data<=16'd12982;
      104803:data<=16'd12243;
      104804:data<=16'd12269;
      104805:data<=16'd11674;
      104806:data<=16'd12407;
      104807:data<=16'd13891;
      104808:data<=16'd13062;
      104809:data<=16'd12807;
      104810:data<=16'd12698;
      104811:data<=16'd11464;
      104812:data<=16'd12417;
      104813:data<=16'd11850;
      104814:data<=16'd7829;
      104815:data<=16'd6225;
      104816:data<=16'd6549;
      104817:data<=16'd6288;
      104818:data<=16'd6279;
      104819:data<=16'd6366;
      104820:data<=16'd7350;
      104821:data<=16'd8125;
      104822:data<=16'd7421;
      104823:data<=16'd7457;
      104824:data<=16'd7485;
      104825:data<=16'd7138;
      104826:data<=16'd8619;
      104827:data<=16'd9744;
      104828:data<=16'd9086;
      104829:data<=16'd8846;
      104830:data<=16'd8931;
      104831:data<=16'd8584;
      104832:data<=16'd8645;
      104833:data<=16'd9620;
      104834:data<=16'd10172;
      104835:data<=16'd9210;
      104836:data<=16'd8657;
      104837:data<=16'd8692;
      104838:data<=16'd7702;
      104839:data<=16'd7920;
      104840:data<=16'd9787;
      104841:data<=16'd10126;
      104842:data<=16'd9289;
      104843:data<=16'd8742;
      104844:data<=16'd8281;
      104845:data<=16'd8484;
      104846:data<=16'd9360;
      104847:data<=16'd9794;
      104848:data<=16'd9265;
      104849:data<=16'd8760;
      104850:data<=16'd8880;
      104851:data<=16'd8260;
      104852:data<=16'd7864;
      104853:data<=16'd9271;
      104854:data<=16'd9975;
      104855:data<=16'd9450;
      104856:data<=16'd8792;
      104857:data<=16'd7511;
      104858:data<=16'd9039;
      104859:data<=16'd13773;
      104860:data<=16'd15666;
      104861:data<=16'd14803;
      104862:data<=16'd13790;
      104863:data<=16'd11762;
      104864:data<=16'd10507;
      104865:data<=16'd10777;
      104866:data<=16'd11001;
      104867:data<=16'd11264;
      104868:data<=16'd10801;
      104869:data<=16'd10097;
      104870:data<=16'd9903;
      104871:data<=16'd8863;
      104872:data<=16'd8853;
      104873:data<=16'd10446;
      104874:data<=16'd10364;
      104875:data<=16'd9312;
      104876:data<=16'd8633;
      104877:data<=16'd7655;
      104878:data<=16'd7423;
      104879:data<=16'd7629;
      104880:data<=16'd7133;
      104881:data<=16'd6416;
      104882:data<=16'd5777;
      104883:data<=16'd5524;
      104884:data<=16'd5148;
      104885:data<=16'd3873;
      104886:data<=16'd2614;
      104887:data<=16'd1980;
      104888:data<=16'd1635;
      104889:data<=16'd1022;
      104890:data<=16'd177;
      104891:data<=-16'd73;
      104892:data<=-16'd632;
      104893:data<=-16'd2135;
      104894:data<=-16'd2860;
      104895:data<=-16'd2867;
      104896:data<=-16'd3357;
      104897:data<=-16'd3527;
      104898:data<=-16'd3404;
      104899:data<=-16'd4854;
      104900:data<=-16'd6598;
      104901:data<=-16'd6114;
      104902:data<=-16'd7051;
      104903:data<=-16'd11159;
      104904:data<=-16'd12891;
      104905:data<=-16'd12841;
      104906:data<=-16'd14242;
      104907:data<=-16'd13929;
      104908:data<=-16'd13051;
      104909:data<=-16'd13916;
      104910:data<=-16'd13379;
      104911:data<=-16'd12296;
      104912:data<=-16'd12753;
      104913:data<=-16'd13544;
      104914:data<=-16'd14178;
      104915:data<=-16'd13863;
      104916:data<=-16'd13153;
      104917:data<=-16'd12865;
      104918:data<=-16'd12349;
      104919:data<=-16'd13086;
      104920:data<=-16'd14230;
      104921:data<=-16'd13532;
      104922:data<=-16'd12916;
      104923:data<=-16'd12754;
      104924:data<=-16'd12417;
      104925:data<=-16'd12863;
      104926:data<=-16'd13288;
      104927:data<=-16'd13540;
      104928:data<=-16'd13494;
      104929:data<=-16'd12210;
      104930:data<=-16'd10628;
      104931:data<=-16'd9497;
      104932:data<=-16'd9949;
      104933:data<=-16'd11696;
      104934:data<=-16'd11509;
      104935:data<=-16'd10141;
      104936:data<=-16'd9709;
      104937:data<=-16'd9297;
      104938:data<=-16'd9295;
      104939:data<=-16'd10066;
      104940:data<=-16'd10658;
      104941:data<=-16'd10272;
      104942:data<=-16'd9235;
      104943:data<=-16'd9229;
      104944:data<=-16'd8965;
      104945:data<=-16'd8505;
      104946:data<=-16'd10190;
      104947:data<=-16'd9056;
      104948:data<=-16'd4006;
      104949:data<=-16'd2587;
      104950:data<=-16'd3301;
      104951:data<=-16'd2202;
      104952:data<=-16'd2692;
      104953:data<=-16'd4402;
      104954:data<=-16'd4605;
      104955:data<=-16'd4219;
      104956:data<=-16'd3991;
      104957:data<=-16'd3673;
      104958:data<=-16'd3512;
      104959:data<=-16'd4402;
      104960:data<=-16'd5427;
      104961:data<=-16'd5002;
      104962:data<=-16'd4786;
      104963:data<=-16'd4948;
      104964:data<=-16'd3961;
      104965:data<=-16'd3967;
      104966:data<=-16'd5560;
      104967:data<=-16'd6002;
      104968:data<=-16'd5300;
      104969:data<=-16'd4942;
      104970:data<=-16'd4522;
      104971:data<=-16'd3894;
      104972:data<=-16'd4566;
      104973:data<=-16'd6122;
      104974:data<=-16'd6220;
      104975:data<=-16'd5448;
      104976:data<=-16'd5244;
      104977:data<=-16'd4934;
      104978:data<=-16'd4863;
      104979:data<=-16'd5947;
      104980:data<=-16'd7059;
      104981:data<=-16'd6616;
      104982:data<=-16'd5588;
      104983:data<=-16'd5480;
      104984:data<=-16'd5033;
      104985:data<=-16'd4364;
      104986:data<=-16'd4796;
      104987:data<=-16'd4651;
      104988:data<=-16'd4040;
      104989:data<=-16'd3849;
      104990:data<=-16'd2939;
      104991:data<=-16'd3657;
      104992:data<=-16'd6587;
      104993:data<=-16'd7633;
      104994:data<=-16'd6855;
      104995:data<=-16'd6355;
      104996:data<=-16'd6605;
      104997:data<=-16'd7620;
      104998:data<=-16'd7347;
      104999:data<=-16'd5491;
      105000:data<=-16'd4441;
      105001:data<=-16'd4334;
      105002:data<=-16'd4014;
      105003:data<=-16'd3359;
      105004:data<=-16'd3137;
      105005:data<=-16'd2714;
      105006:data<=-16'd960;
      105007:data<=16'd168;
      105008:data<=16'd318;
      105009:data<=16'd879;
      105010:data<=16'd496;
      105011:data<=16'd432;
      105012:data<=16'd2291;
      105013:data<=16'd3389;
      105014:data<=16'd3453;
      105015:data<=16'd3530;
      105016:data<=16'd3263;
      105017:data<=16'd3468;
      105018:data<=16'd4037;
      105019:data<=16'd4924;
      105020:data<=16'd6032;
      105021:data<=16'd5985;
      105022:data<=16'd5999;
      105023:data<=16'd6291;
      105024:data<=16'd5591;
      105025:data<=16'd6209;
      105026:data<=16'd7990;
      105027:data<=16'd8264;
      105028:data<=16'd7835;
      105029:data<=16'd7353;
      105030:data<=16'd6998;
      105031:data<=16'd7450;
      105032:data<=16'd8266;
      105033:data<=16'd9394;
      105034:data<=16'd9365;
      105035:data<=16'd8069;
      105036:data<=16'd9812;
      105037:data<=16'd13866;
      105038:data<=16'd15579;
      105039:data<=16'd15978;
      105040:data<=16'd16409;
      105041:data<=16'd15732;
      105042:data<=16'd15111;
      105043:data<=16'd14915;
      105044:data<=16'd14149;
      105045:data<=16'd14120;
      105046:data<=16'd15127;
      105047:data<=16'd15120;
      105048:data<=16'd14090;
      105049:data<=16'd13449;
      105050:data<=16'd13000;
      105051:data<=16'd12701;
      105052:data<=16'd13258;
      105053:data<=16'd13747;
      105054:data<=16'd13220;
      105055:data<=16'd12686;
      105056:data<=16'd12384;
      105057:data<=16'd11734;
      105058:data<=16'd11685;
      105059:data<=16'd12422;
      105060:data<=16'd12636;
      105061:data<=16'd12243;
      105062:data<=16'd11756;
      105063:data<=16'd11449;
      105064:data<=16'd11759;
      105065:data<=16'd12466;
      105066:data<=16'd13059;
      105067:data<=16'd12983;
      105068:data<=16'd12158;
      105069:data<=16'd11483;
      105070:data<=16'd10898;
      105071:data<=16'd10445;
      105072:data<=16'd11041;
      105073:data<=16'd11661;
      105074:data<=16'd11315;
      105075:data<=16'd10443;
      105076:data<=16'd9182;
      105077:data<=16'd8298;
      105078:data<=16'd8264;
      105079:data<=16'd9206;
      105080:data<=16'd9852;
      105081:data<=16'd6499;
      105082:data<=16'd1659;
      105083:data<=16'd785;
      105084:data<=16'd1137;
      105085:data<=16'd1292;
      105086:data<=16'd2863;
      105087:data<=16'd2528;
      105088:data<=16'd1049;
      105089:data<=16'd1530;
      105090:data<=16'd1387;
      105091:data<=16'd505;
      105092:data<=16'd581;
      105093:data<=16'd425;
      105094:data<=16'd11;
      105095:data<=-16'd364;
      105096:data<=-16'd676;
      105097:data<=-16'd707;
      105098:data<=-16'd1366;
      105099:data<=-16'd2684;
      105100:data<=-16'd3773;
      105101:data<=-16'd4015;
      105102:data<=-16'd3748;
      105103:data<=-16'd3927;
      105104:data<=-16'd3911;
      105105:data<=-16'd4378;
      105106:data<=-16'd6310;
      105107:data<=-16'd7084;
      105108:data<=-16'd6537;
      105109:data<=-16'd6434;
      105110:data<=-16'd6152;
      105111:data<=-16'd6805;
      105112:data<=-16'd8376;
      105113:data<=-16'd8469;
      105114:data<=-16'd8076;
      105115:data<=-16'd8437;
      105116:data<=-16'd8404;
      105117:data<=-16'd7758;
      105118:data<=-16'd8117;
      105119:data<=-16'd9826;
      105120:data<=-16'd10255;
      105121:data<=-16'd9483;
      105122:data<=-16'd9313;
      105123:data<=-16'd8793;
      105124:data<=-16'd8998;
      105125:data<=-16'd9097;
      105126:data<=-16'd6021;
      105127:data<=-16'd3889;
      105128:data<=-16'd4296;
      105129:data<=-16'd3627;
      105130:data<=-16'd4255;
      105131:data<=-16'd6737;
      105132:data<=-16'd7793;
      105133:data<=-16'd7990;
      105134:data<=-16'd7832;
      105135:data<=-16'd7847;
      105136:data<=-16'd8317;
      105137:data<=-16'd7749;
      105138:data<=-16'd7877;
      105139:data<=-16'd9332;
      105140:data<=-16'd9506;
      105141:data<=-16'd9027;
      105142:data<=-16'd8907;
      105143:data<=-16'd8607;
      105144:data<=-16'd8821;
      105145:data<=-16'd9721;
      105146:data<=-16'd10179;
      105147:data<=-16'd9697;
      105148:data<=-16'd9468;
      105149:data<=-16'd9682;
      105150:data<=-16'd9144;
      105151:data<=-16'd9097;
      105152:data<=-16'd10076;
      105153:data<=-16'd10237;
      105154:data<=-16'd9840;
      105155:data<=-16'd9676;
      105156:data<=-16'd9294;
      105157:data<=-16'd8678;
      105158:data<=-16'd8916;
      105159:data<=-16'd10373;
      105160:data<=-16'd10422;
      105161:data<=-16'd9309;
      105162:data<=-16'd9544;
      105163:data<=-16'd8837;
      105164:data<=-16'd8081;
      105165:data<=-16'd9826;
      105166:data<=-16'd10134;
      105167:data<=-16'd9561;
      105168:data<=-16'd10208;
      105169:data<=-16'd9047;
      105170:data<=-16'd9697;
      105171:data<=-16'd14342;
      105172:data<=-16'd16427;
      105173:data<=-16'd15750;
      105174:data<=-16'd15655;
      105175:data<=-16'd14945;
      105176:data<=-16'd13635;
      105177:data<=-16'd12754;
      105178:data<=-16'd12753;
      105179:data<=-16'd13649;
      105180:data<=-16'd13652;
      105181:data<=-16'd12346;
      105182:data<=-16'd11429;
      105183:data<=-16'd11235;
      105184:data<=-16'd11176;
      105185:data<=-16'd11561;
      105186:data<=-16'd12005;
      105187:data<=-16'd11345;
      105188:data<=-16'd10457;
      105189:data<=-16'd9940;
      105190:data<=-16'd9044;
      105191:data<=-16'd9172;
      105192:data<=-16'd10404;
      105193:data<=-16'd10364;
      105194:data<=-16'd9236;
      105195:data<=-16'd8348;
      105196:data<=-16'd7990;
      105197:data<=-16'd7185;
      105198:data<=-16'd5175;
      105199:data<=-16'd3985;
      105200:data<=-16'd3776;
      105201:data<=-16'd3078;
      105202:data<=-16'd2925;
      105203:data<=-16'd2628;
      105204:data<=-16'd1416;
      105205:data<=-16'd340;
      105206:data<=16'd1027;
      105207:data<=16'd1510;
      105208:data<=16'd1037;
      105209:data<=16'd1639;
      105210:data<=16'd1921;
      105211:data<=16'd2563;
      105212:data<=16'd4564;
      105213:data<=16'd4875;
      105214:data<=16'd5805;
      105215:data<=16'd9730;
      105216:data<=16'd11984;
      105217:data<=16'd11806;
      105218:data<=16'd12378;
      105219:data<=16'd13503;
      105220:data<=16'd13591;
      105221:data<=16'd12700;
      105222:data<=16'd12298;
      105223:data<=16'd12343;
      105224:data<=16'd12552;
      105225:data<=16'd13679;
      105226:data<=16'd14013;
      105227:data<=16'd13141;
      105228:data<=16'd13254;
      105229:data<=16'd13462;
      105230:data<=16'd12698;
      105231:data<=16'd12601;
      105232:data<=16'd13846;
      105233:data<=16'd14687;
      105234:data<=16'd13837;
      105235:data<=16'd13206;
      105236:data<=16'd13264;
      105237:data<=16'd12652;
      105238:data<=16'd13289;
      105239:data<=16'd14510;
      105240:data<=16'd13664;
      105241:data<=16'd13044;
      105242:data<=16'd13021;
      105243:data<=16'd12116;
      105244:data<=16'd12395;
      105245:data<=16'd13396;
      105246:data<=16'd13174;
      105247:data<=16'd12756;
      105248:data<=16'd12771;
      105249:data<=16'd12675;
      105250:data<=16'd12037;
      105251:data<=16'd12128;
      105252:data<=16'd13881;
      105253:data<=16'd14307;
      105254:data<=16'd13063;
      105255:data<=16'd12777;
      105256:data<=16'd11888;
      105257:data<=16'd10966;
      105258:data<=16'd12316;
      105259:data<=16'd11271;
      105260:data<=16'd6673;
      105261:data<=16'd4898;
      105262:data<=16'd5629;
      105263:data<=16'd4817;
      105264:data<=16'd3983;
      105265:data<=16'd4243;
      105266:data<=16'd4469;
      105267:data<=16'd4592;
      105268:data<=16'd4356;
      105269:data<=16'd3773;
      105270:data<=16'd3250;
      105271:data<=16'd3686;
      105272:data<=16'd5559;
      105273:data<=16'd6119;
      105274:data<=16'd4846;
      105275:data<=16'd4560;
      105276:data<=16'd4396;
      105277:data<=16'd4152;
      105278:data<=16'd5388;
      105279:data<=16'd5958;
      105280:data<=16'd5544;
      105281:data<=16'd5673;
      105282:data<=16'd5259;
      105283:data<=16'd4642;
      105284:data<=16'd5107;
      105285:data<=16'd6364;
      105286:data<=16'd7015;
      105287:data<=16'd6117;
      105288:data<=16'd5691;
      105289:data<=16'd5873;
      105290:data<=16'd5104;
      105291:data<=16'd5729;
      105292:data<=16'd7274;
      105293:data<=16'd6842;
      105294:data<=16'd6134;
      105295:data<=16'd5938;
      105296:data<=16'd5453;
      105297:data<=16'd5691;
      105298:data<=16'd6428;
      105299:data<=16'd6554;
      105300:data<=16'd6134;
      105301:data<=16'd6070;
      105302:data<=16'd5876;
      105303:data<=16'd5507;
      105304:data<=16'd8137;
      105305:data<=16'd11715;
      105306:data<=16'd11264;
      105307:data<=16'd9937;
      105308:data<=16'd10031;
      105309:data<=16'd9511;
      105310:data<=16'd9039;
      105311:data<=16'd7964;
      105312:data<=16'd6091;
      105313:data<=16'd5300;
      105314:data<=16'd4930;
      105315:data<=16'd4902;
      105316:data<=16'd4851;
      105317:data<=16'd3363;
      105318:data<=16'd1582;
      105319:data<=16'd446;
      105320:data<=16'd516;
      105321:data<=16'd1183;
      105322:data<=16'd588;
      105323:data<=16'd138;
      105324:data<=-16'd373;
      105325:data<=-16'd2294;
      105326:data<=-16'd3004;
      105327:data<=-16'd2676;
      105328:data<=-16'd2776;
      105329:data<=-16'd2496;
      105330:data<=-16'd2928;
      105331:data<=-16'd3653;
      105332:data<=-16'd3456;
      105333:data<=-16'd3295;
      105334:data<=-16'd3157;
      105335:data<=-16'd3456;
      105336:data<=-16'd4170;
      105337:data<=-16'd4545;
      105338:data<=-16'd5395;
      105339:data<=-16'd5949;
      105340:data<=-16'd5692;
      105341:data<=-16'd5673;
      105342:data<=-16'd5568;
      105343:data<=-16'd5521;
      105344:data<=-16'd5779;
      105345:data<=-16'd6959;
      105346:data<=-16'd8366;
      105347:data<=-16'd7447;
      105348:data<=-16'd8205;
      105349:data<=-16'd12609;
      105350:data<=-16'd14198;
      105351:data<=-16'd14070;
      105352:data<=-16'd15218;
      105353:data<=-16'd14730;
      105354:data<=-16'd14609;
      105355:data<=-16'd15192;
      105356:data<=-16'd13838;
      105357:data<=-16'd13418;
      105358:data<=-16'd14381;
      105359:data<=-16'd14668;
      105360:data<=-16'd14560;
      105361:data<=-16'd14081;
      105362:data<=-16'd13617;
      105363:data<=-16'd12756;
      105364:data<=-16'd12502;
      105365:data<=-16'd14287;
      105366:data<=-16'd14572;
      105367:data<=-16'd13242;
      105368:data<=-16'd13042;
      105369:data<=-16'd12117;
      105370:data<=-16'd11535;
      105371:data<=-16'd12841;
      105372:data<=-16'd13164;
      105373:data<=-16'd12475;
      105374:data<=-16'd12054;
      105375:data<=-16'd11693;
      105376:data<=-16'd11227;
      105377:data<=-16'd10558;
      105378:data<=-16'd11054;
      105379:data<=-16'd11885;
      105380:data<=-16'd11094;
      105381:data<=-16'd10552;
      105382:data<=-16'd10502;
      105383:data<=-16'd9693;
      105384:data<=-16'd9624;
      105385:data<=-16'd10504;
      105386:data<=-16'd10815;
      105387:data<=-16'd9937;
      105388:data<=-16'd8978;
      105389:data<=-16'd9051;
      105390:data<=-16'd8856;
      105391:data<=-16'd9036;
      105392:data<=-16'd10044;
      105393:data<=-16'd7538;
      105394:data<=-16'd2749;
      105395:data<=-16'd1556;
      105396:data<=-16'd1748;
      105397:data<=-16'd861;
      105398:data<=-16'd2570;
      105399:data<=-16'd5386;
      105400:data<=-16'd5018;
      105401:data<=-16'd4062;
      105402:data<=-16'd4325;
      105403:data<=-16'd3682;
      105404:data<=-16'd3685;
      105405:data<=-16'd4937;
      105406:data<=-16'd4962;
      105407:data<=-16'd4760;
      105408:data<=-16'd4805;
      105409:data<=-16'd3924;
      105410:data<=-16'd3365;
      105411:data<=-16'd2977;
      105412:data<=-16'd2382;
      105413:data<=-16'd2619;
      105414:data<=-16'd2601;
      105415:data<=-16'd1996;
      105416:data<=-16'd1632;
      105417:data<=-16'd939;
      105418:data<=16'd76;
      105419:data<=16'd949;
      105420:data<=16'd1441;
      105421:data<=16'd1779;
      105422:data<=16'd1949;
      105423:data<=16'd1441;
      105424:data<=16'd2382;
      105425:data<=16'd4523;
      105426:data<=16'd4132;
      105427:data<=16'd3356;
      105428:data<=16'd4068;
      105429:data<=16'd3883;
      105430:data<=16'd4601;
      105431:data<=16'd6328;
      105432:data<=16'd6325;
      105433:data<=16'd6175;
      105434:data<=16'd6282;
      105435:data<=16'd6188;
      105436:data<=16'd6763;
      105437:data<=16'd5747;
      105438:data<=16'd3031;
      105439:data<=16'd1595;
      105440:data<=16'd1427;
      105441:data<=16'd1600;
      105442:data<=16'd1597;
      105443:data<=16'd1536;
      105444:data<=16'd2500;
      105445:data<=16'd3560;
      105446:data<=16'd3767;
      105447:data<=16'd3883;
      105448:data<=16'd3820;
      105449:data<=16'd3495;
      105450:data<=16'd3704;
      105451:data<=16'd4799;
      105452:data<=16'd5947;
      105453:data<=16'd6161;
      105454:data<=16'd5959;
      105455:data<=16'd5636;
      105456:data<=16'd5049;
      105457:data<=16'd5538;
      105458:data<=16'd6921;
      105459:data<=16'd7313;
      105460:data<=16'd7056;
      105461:data<=16'd7033;
      105462:data<=16'd6739;
      105463:data<=16'd6381;
      105464:data<=16'd7059;
      105465:data<=16'd8763;
      105466:data<=16'd10055;
      105467:data<=16'd10261;
      105468:data<=16'd10020;
      105469:data<=16'd9559;
      105470:data<=16'd9527;
      105471:data<=16'd10643;
      105472:data<=16'd11285;
      105473:data<=16'd10646;
      105474:data<=16'd10310;
      105475:data<=16'd9976;
      105476:data<=16'd9256;
      105477:data<=16'd9650;
      105478:data<=16'd10584;
      105479:data<=16'd10792;
      105480:data<=16'd10091;
      105481:data<=16'd8916;
      105482:data<=16'd10340;
      105483:data<=16'd14428;
      105484:data<=16'd16419;
      105485:data<=16'd16236;
      105486:data<=16'd16043;
      105487:data<=16'd15249;
      105488:data<=16'd14427;
      105489:data<=16'd13624;
      105490:data<=16'd13092;
      105491:data<=16'd14154;
      105492:data<=16'd14460;
      105493:data<=16'd13233;
      105494:data<=16'd12783;
      105495:data<=16'd12058;
      105496:data<=16'd10954;
      105497:data<=16'd11307;
      105498:data<=16'd12003;
      105499:data<=16'd11746;
      105500:data<=16'd10927;
      105501:data<=16'd10276;
      105502:data<=16'd9726;
      105503:data<=16'd9098;
      105504:data<=16'd9442;
      105505:data<=16'd9897;
      105506:data<=16'd9451;
      105507:data<=16'd9430;
      105508:data<=16'd8774;
      105509:data<=16'd7368;
      105510:data<=16'd7762;
      105511:data<=16'd8621;
      105512:data<=16'd8392;
      105513:data<=16'd7991;
      105514:data<=16'd7212;
      105515:data<=16'd6536;
      105516:data<=16'd6270;
      105517:data<=16'd5535;
      105518:data<=16'd4928;
      105519:data<=16'd4987;
      105520:data<=16'd4831;
      105521:data<=16'd4087;
      105522:data<=16'd3691;
      105523:data<=16'd3087;
      105524:data<=16'd1095;
      105525:data<=16'd294;
      105526:data<=16'd86;
      105527:data<=-16'd3753;
      105528:data<=-16'd7277;
      105529:data<=-16'd7090;
      105530:data<=-16'd7744;
      105531:data<=-16'd9498;
      105532:data<=-16'd10299;
      105533:data<=-16'd11224;
      105534:data<=-16'd11684;
      105535:data<=-16'd11300;
      105536:data<=-16'd10954;
      105537:data<=-16'd11436;
      105538:data<=-16'd12730;
      105539:data<=-16'd12609;
      105540:data<=-16'd11699;
      105541:data<=-16'd12000;
      105542:data<=-16'd11758;
      105543:data<=-16'd11421;
      105544:data<=-16'd12577;
      105545:data<=-16'd13039;
      105546:data<=-16'd12242;
      105547:data<=-16'd12013;
      105548:data<=-16'd12134;
      105549:data<=-16'd11550;
      105550:data<=-16'd11618;
      105551:data<=-16'd13000;
      105552:data<=-16'd12903;
      105553:data<=-16'd11835;
      105554:data<=-16'd12038;
      105555:data<=-16'd11329;
      105556:data<=-16'd10401;
      105557:data<=-16'd11538;
      105558:data<=-16'd12339;
      105559:data<=-16'd12111;
      105560:data<=-16'd11820;
      105561:data<=-16'd11276;
      105562:data<=-16'd10941;
      105563:data<=-16'd10836;
      105564:data<=-16'd11731;
      105565:data<=-16'd12519;
      105566:data<=-16'd11486;
      105567:data<=-16'd11520;
      105568:data<=-16'd11526;
      105569:data<=-16'd9850;
      105570:data<=-16'd10906;
      105571:data<=-16'd11065;
      105572:data<=-16'd6498;
      105573:data<=-16'd4270;
      105574:data<=-16'd4971;
      105575:data<=-16'd4479;
      105576:data<=-16'd4469;
      105577:data<=-16'd5231;
      105578:data<=-16'd5900;
      105579:data<=-16'd6070;
      105580:data<=-16'd5600;
      105581:data<=-16'd6047;
      105582:data<=-16'd5967;
      105583:data<=-16'd5156;
      105584:data<=-16'd6543;
      105585:data<=-16'd7752;
      105586:data<=-16'd6872;
      105587:data<=-16'd6426;
      105588:data<=-16'd6211;
      105589:data<=-16'd5638;
      105590:data<=-16'd6228;
      105591:data<=-16'd7718;
      105592:data<=-16'd7855;
      105593:data<=-16'd6566;
      105594:data<=-16'd6454;
      105595:data<=-16'd6737;
      105596:data<=-16'd6020;
      105597:data<=-16'd6904;
      105598:data<=-16'd8197;
      105599:data<=-16'd6913;
      105600:data<=-16'd5327;
      105601:data<=-16'd4663;
      105602:data<=-16'd4190;
      105603:data<=-16'd4663;
      105604:data<=-16'd5614;
      105605:data<=-16'd5915;
      105606:data<=-16'd5488;
      105607:data<=-16'd5137;
      105608:data<=-16'd5143;
      105609:data<=-16'd4655;
      105610:data<=-16'd4775;
      105611:data<=-16'd5808;
      105612:data<=-16'd5785;
      105613:data<=-16'd5655;
      105614:data<=-16'd5571;
      105615:data<=-16'd4868;
      105616:data<=-16'd7303;
      105617:data<=-16'd11985;
      105618:data<=-16'd13083;
      105619:data<=-16'd11897;
      105620:data<=-16'd11676;
      105621:data<=-16'd11138;
      105622:data<=-16'd10354;
      105623:data<=-16'd10235;
      105624:data<=-16'd9608;
      105625:data<=-16'd8543;
      105626:data<=-16'd8044;
      105627:data<=-16'd7436;
      105628:data<=-16'd6704;
      105629:data<=-16'd6513;
      105630:data<=-16'd5506;
      105631:data<=-16'd3644;
      105632:data<=-16'd3084;
      105633:data<=-16'd3289;
      105634:data<=-16'd2866;
      105635:data<=-16'd2328;
      105636:data<=-16'd1480;
      105637:data<=-16'd74;
      105638:data<=16'd769;
      105639:data<=16'd763;
      105640:data<=16'd1215;
      105641:data<=16'd2118;
      105642:data<=16'd1917;
      105643:data<=16'd1983;
      105644:data<=16'd3748;
      105645:data<=16'd4482;
      105646:data<=16'd4146;
      105647:data<=16'd4761;
      105648:data<=16'd4701;
      105649:data<=16'd4388;
      105650:data<=16'd5595;
      105651:data<=16'd6646;
      105652:data<=16'd6802;
      105653:data<=16'd6642;
      105654:data<=16'd6546;
      105655:data<=16'd6769;
      105656:data<=16'd6664;
      105657:data<=16'd7501;
      105658:data<=16'd8833;
      105659:data<=16'd8108;
      105660:data<=16'd9056;
      105661:data<=16'd12966;
      105662:data<=16'd14149;
      105663:data<=16'd13864;
      105664:data<=16'd15512;
      105665:data<=16'd15852;
      105666:data<=16'd14058;
      105667:data<=16'd12646;
      105668:data<=16'd11956;
      105669:data<=16'd11711;
      105670:data<=16'd12299;
      105671:data<=16'd13244;
      105672:data<=16'd12883;
      105673:data<=16'd11966;
      105674:data<=16'd12002;
      105675:data<=16'd11365;
      105676:data<=16'd11038;
      105677:data<=16'd12901;
      105678:data<=16'd13700;
      105679:data<=16'd12672;
      105680:data<=16'd12249;
      105681:data<=16'd11762;
      105682:data<=16'd11274;
      105683:data<=16'd12061;
      105684:data<=16'd12950;
      105685:data<=16'd12442;
      105686:data<=16'd11391;
      105687:data<=16'd11406;
      105688:data<=16'd11474;
      105689:data<=16'd11009;
      105690:data<=16'd11576;
      105691:data<=16'd11811;
      105692:data<=16'd10812;
      105693:data<=16'd10624;
      105694:data<=16'd10578;
      105695:data<=16'd9864;
      105696:data<=16'd9812;
      105697:data<=16'd10615;
      105698:data<=16'd11341;
      105699:data<=16'd10666;
      105700:data<=16'd9617;
      105701:data<=16'd9438;
      105702:data<=16'd8378;
      105703:data<=16'd8448;
      105704:data<=16'd10352;
      105705:data<=16'd7902;
      105706:data<=16'd2907;
      105707:data<=16'd2111;
      105708:data<=16'd2701;
      105709:data<=16'd2156;
      105710:data<=16'd2839;
      105711:data<=16'd3624;
      105712:data<=16'd3315;
      105713:data<=16'd3330;
      105714:data<=16'd3386;
      105715:data<=16'd2695;
      105716:data<=16'd2716;
      105717:data<=16'd4190;
      105718:data<=16'd4966;
      105719:data<=16'd4284;
      105720:data<=16'd3735;
      105721:data<=16'd3298;
      105722:data<=16'd2890;
      105723:data<=16'd3601;
      105724:data<=16'd4602;
      105725:data<=16'd4549;
      105726:data<=16'd4197;
      105727:data<=16'd4264;
      105728:data<=16'd3977;
      105729:data<=16'd3313;
      105730:data<=16'd3278;
      105731:data<=16'd3488;
      105732:data<=16'd3219;
      105733:data<=16'd3172;
      105734:data<=16'd3812;
      105735:data<=16'd4470;
      105736:data<=16'd3906;
      105737:data<=16'd2171;
      105738:data<=16'd1139;
      105739:data<=16'd984;
      105740:data<=16'd560;
      105741:data<=16'd293;
      105742:data<=16'd340;
      105743:data<=16'd77;
      105744:data<=-16'd517;
      105745:data<=-16'd920;
      105746:data<=-16'd494;
      105747:data<=-16'd437;
      105748:data<=-16'd1442;
      105749:data<=-16'd798;
      105750:data<=16'd1436;
      105751:data<=16'd1753;
      105752:data<=16'd732;
      105753:data<=16'd675;
      105754:data<=16'd907;
      105755:data<=16'd751;
      105756:data<=16'd92;
      105757:data<=-16'd1395;
      105758:data<=-16'd2396;
      105759:data<=-16'd2015;
      105760:data<=-16'd1829;
      105761:data<=-16'd2234;
      105762:data<=-16'd2214;
      105763:data<=-16'd2863;
      105764:data<=-16'd4487;
      105765:data<=-16'd4702;
      105766:data<=-16'd3768;
      105767:data<=-16'd3847;
      105768:data<=-16'd4176;
      105769:data<=-16'd4360;
      105770:data<=-16'd5582;
      105771:data<=-16'd6526;
      105772:data<=-16'd6249;
      105773:data<=-16'd6322;
      105774:data<=-16'd6337;
      105775:data<=-16'd5708;
      105776:data<=-16'd6501;
      105777:data<=-16'd8255;
      105778:data<=-16'd8261;
      105779:data<=-16'd7359;
      105780:data<=-16'd7520;
      105781:data<=-16'd7768;
      105782:data<=-16'd7406;
      105783:data<=-16'd7830;
      105784:data<=-16'd8799;
      105785:data<=-16'd8601;
      105786:data<=-16'd8003;
      105787:data<=-16'd8164;
      105788:data<=-16'd8075;
      105789:data<=-16'd8029;
      105790:data<=-16'd9097;
      105791:data<=-16'd9643;
      105792:data<=-16'd8705;
      105793:data<=-16'd8787;
      105794:data<=-16'd10898;
      105795:data<=-16'd12427;
      105796:data<=-16'd12762;
      105797:data<=-16'd13524;
      105798:data<=-16'd13628;
      105799:data<=-16'd12998;
      105800:data<=-16'd13885;
      105801:data<=-16'd14592;
      105802:data<=-16'd13769;
      105803:data<=-16'd14029;
      105804:data<=-16'd14804;
      105805:data<=-16'd14322;
      105806:data<=-16'd13863;
      105807:data<=-16'd13209;
      105808:data<=-16'd11988;
      105809:data<=-16'd12128;
      105810:data<=-16'd13373;
      105811:data<=-16'd13517;
      105812:data<=-16'd12557;
      105813:data<=-16'd11767;
      105814:data<=-16'd10974;
      105815:data<=-16'd10094;
      105816:data<=-16'd10499;
      105817:data<=-16'd11583;
      105818:data<=-16'd11339;
      105819:data<=-16'd10663;
      105820:data<=-16'd10525;
      105821:data<=-16'd9821;
      105822:data<=-16'd9219;
      105823:data<=-16'd9814;
      105824:data<=-16'd10120;
      105825:data<=-16'd9523;
      105826:data<=-16'd9256;
      105827:data<=-16'd8997;
      105828:data<=-16'd8335;
      105829:data<=-16'd8775;
      105830:data<=-16'd10044;
      105831:data<=-16'd9884;
      105832:data<=-16'd8552;
      105833:data<=-16'd7997;
      105834:data<=-16'd8032;
      105835:data<=-16'd7413;
      105836:data<=-16'd6939;
      105837:data<=-16'd7090;
      105838:data<=-16'd5450;
      105839:data<=-16'd2097;
      105840:data<=-16'd655;
      105841:data<=-16'd928;
      105842:data<=-16'd341;
      105843:data<=16'd904;
      105844:data<=16'd1924;
      105845:data<=16'd2317;
      105846:data<=16'd2332;
      105847:data<=16'd2616;
      105848:data<=16'd2487;
      105849:data<=16'd2575;
      105850:data<=16'd4046;
      105851:data<=16'd4981;
      105852:data<=16'd4783;
      105853:data<=16'd4913;
      105854:data<=16'd4754;
      105855:data<=16'd4560;
      105856:data<=16'd5738;
      105857:data<=16'd7007;
      105858:data<=16'd6995;
      105859:data<=16'd6673;
      105860:data<=16'd6658;
      105861:data<=16'd6517;
      105862:data<=16'd6707;
      105863:data<=16'd7794;
      105864:data<=16'd8636;
      105865:data<=16'd8298;
      105866:data<=16'd7959;
      105867:data<=16'd8625;
      105868:data<=16'd9370;
      105869:data<=16'd9591;
      105870:data<=16'd10264;
      105871:data<=16'd11101;
      105872:data<=16'd10809;
      105873:data<=16'd10182;
      105874:data<=16'd9964;
      105875:data<=16'd9885;
      105876:data<=16'd10689;
      105877:data<=16'd11671;
      105878:data<=16'd11201;
      105879:data<=16'd10331;
      105880:data<=16'd10398;
      105881:data<=16'd10643;
      105882:data<=16'd9812;
      105883:data<=16'd8140;
      105884:data<=16'd7004;
      105885:data<=16'd6514;
      105886:data<=16'd6299;
      105887:data<=16'd6131;
      105888:data<=16'd5510;
      105889:data<=16'd5877;
      105890:data<=16'd7489;
      105891:data<=16'd7708;
      105892:data<=16'd7009;
      105893:data<=16'd7069;
      105894:data<=16'd6980;
      105895:data<=16'd6789;
      105896:data<=16'd7280;
      105897:data<=16'd7915;
      105898:data<=16'd7700;
      105899:data<=16'd6902;
      105900:data<=16'd6843;
      105901:data<=16'd6793;
      105902:data<=16'd6610;
      105903:data<=16'd7668;
      105904:data<=16'd8029;
      105905:data<=16'd7219;
      105906:data<=16'd7294;
      105907:data<=16'd6760;
      105908:data<=16'd5852;
      105909:data<=16'd6878;
      105910:data<=16'd8040;
      105911:data<=16'd7758;
      105912:data<=16'd7141;
      105913:data<=16'd6975;
      105914:data<=16'd6751;
      105915:data<=16'd6140;
      105916:data<=16'd6576;
      105917:data<=16'd7436;
      105918:data<=16'd7119;
      105919:data<=16'd6939;
      105920:data<=16'd6484;
      105921:data<=16'd5483;
      105922:data<=16'd5911;
      105923:data<=16'd6711;
      105924:data<=16'd6942;
      105925:data<=16'd6675;
      105926:data<=16'd5780;
      105927:data<=16'd6810;
      105928:data<=16'd9171;
      105929:data<=16'd10275;
      105930:data<=16'd10948;
      105931:data<=16'd10384;
      105932:data<=16'd9351;
      105933:data<=16'd9556;
      105934:data<=16'd7893;
      105935:data<=16'd5930;
      105936:data<=16'd7130;
      105937:data<=16'd7794;
      105938:data<=16'd6766;
      105939:data<=16'd6266;
      105940:data<=16'd5702;
      105941:data<=16'd5375;
      105942:data<=16'd5729;
      105943:data<=16'd5532;
      105944:data<=16'd4805;
      105945:data<=16'd4405;
      105946:data<=16'd4003;
      105947:data<=16'd3486;
      105948:data<=16'd3647;
      105949:data<=16'd2886;
      105950:data<=16'd464;
      105951:data<=-16'd302;
      105952:data<=16'd321;
      105953:data<=16'd14;
      105954:data<=-16'd258;
      105955:data<=-16'd1063;
      105956:data<=-16'd2537;
      105957:data<=-16'd3022;
      105958:data<=-16'd3248;
      105959:data<=-16'd3565;
      105960:data<=-16'd3759;
      105961:data<=-16'd3679;
      105962:data<=-16'd3386;
      105963:data<=-16'd4921;
      105964:data<=-16'd6555;
      105965:data<=-16'd5853;
      105966:data<=-16'd5582;
      105967:data<=-16'd5671;
      105968:data<=-16'd5447;
      105969:data<=-16'd6558;
      105970:data<=-16'd7115;
      105971:data<=-16'd7949;
      105972:data<=-16'd10903;
      105973:data<=-16'd12140;
      105974:data<=-16'd11359;
      105975:data<=-16'd11693;
      105976:data<=-16'd12701;
      105977:data<=-16'd13010;
      105978:data<=-16'd12487;
      105979:data<=-16'd12240;
      105980:data<=-16'd12113;
      105981:data<=-16'd11364;
      105982:data<=-16'd11796;
      105983:data<=-16'd12915;
      105984:data<=-16'd12813;
      105985:data<=-16'd12480;
      105986:data<=-16'd12107;
      105987:data<=-16'd11703;
      105988:data<=-16'd11861;
      105989:data<=-16'd12126;
      105990:data<=-16'd12604;
      105991:data<=-16'd12558;
      105992:data<=-16'd11864;
      105993:data<=-16'd11699;
      105994:data<=-16'd11119;
      105995:data<=-16'd10904;
      105996:data<=-16'd12232;
      105997:data<=-16'd12487;
      105998:data<=-16'd11684;
      105999:data<=-16'd11690;
      106000:data<=-16'd11036;
      106001:data<=-16'd9192;
      106002:data<=-16'd8364;
      106003:data<=-16'd9327;
      106004:data<=-16'd9781;
      106005:data<=-16'd9068;
      106006:data<=-16'd9144;
      106007:data<=-16'd9021;
      106008:data<=-16'd8296;
      106009:data<=-16'd9000;
      106010:data<=-16'd9489;
      106011:data<=-16'd8828;
      106012:data<=-16'd8637;
      106013:data<=-16'd8207;
      106014:data<=-16'd7882;
      106015:data<=-16'd8012;
      106016:data<=-16'd6558;
      106017:data<=-16'd4419;
      106018:data<=-16'd3726;
      106019:data<=-16'd3853;
      106020:data<=-16'd3533;
      106021:data<=-16'd2837;
      106022:data<=-16'd3236;
      106023:data<=-16'd4561;
      106024:data<=-16'd4846;
      106025:data<=-16'd4408;
      106026:data<=-16'd4319;
      106027:data<=-16'd4073;
      106028:data<=-16'd3876;
      106029:data<=-16'd4657;
      106030:data<=-16'd5560;
      106031:data<=-16'd5175;
      106032:data<=-16'd4557;
      106033:data<=-16'd4538;
      106034:data<=-16'd4149;
      106035:data<=-16'd4482;
      106036:data<=-16'd5923;
      106037:data<=-16'd6053;
      106038:data<=-16'd5433;
      106039:data<=-16'd5570;
      106040:data<=-16'd5115;
      106041:data<=-16'd4316;
      106042:data<=-16'd4869;
      106043:data<=-16'd5967;
      106044:data<=-16'd5984;
      106045:data<=-16'd5419;
      106046:data<=-16'd5356;
      106047:data<=-16'd5068;
      106048:data<=-16'd4384;
      106049:data<=-16'd4184;
      106050:data<=-16'd3867;
      106051:data<=-16'd3489;
      106052:data<=-16'd3620;
      106053:data<=-16'd3371;
      106054:data<=-16'd2990;
      106055:data<=-16'd2334;
      106056:data<=-16'd702;
      106057:data<=-16'd194;
      106058:data<=-16'd444;
      106059:data<=16'd513;
      106060:data<=-16'd555;
      106061:data<=-16'd3774;
      106062:data<=-16'd3780;
      106063:data<=-16'd1507;
      106064:data<=-16'd1134;
      106065:data<=-16'd1583;
      106066:data<=-16'd1248;
      106067:data<=-16'd1010;
      106068:data<=-16'd1134;
      106069:data<=-16'd884;
      106070:data<=-16'd79;
      106071:data<=16'd491;
      106072:data<=16'd591;
      106073:data<=16'd746;
      106074:data<=16'd936;
      106075:data<=16'd1477;
      106076:data<=16'd2572;
      106077:data<=16'd3104;
      106078:data<=16'd2984;
      106079:data<=16'd3196;
      106080:data<=16'd3451;
      106081:data<=16'd3670;
      106082:data<=16'd4639;
      106083:data<=16'd5700;
      106084:data<=16'd5720;
      106085:data<=16'd5395;
      106086:data<=16'd5474;
      106087:data<=16'd5476;
      106088:data<=16'd5826;
      106089:data<=16'd6987;
      106090:data<=16'd7550;
      106091:data<=16'd7230;
      106092:data<=16'd7409;
      106093:data<=16'd7638;
      106094:data<=16'd7162;
      106095:data<=16'd7444;
      106096:data<=16'd8739;
      106097:data<=16'd8919;
      106098:data<=16'd8214;
      106099:data<=16'd8436;
      106100:data<=16'd8504;
      106101:data<=16'd8155;
      106102:data<=16'd9081;
      106103:data<=16'd9894;
      106104:data<=16'd10358;
      106105:data<=16'd12663;
      106106:data<=16'd14407;
      106107:data<=16'd13702;
      106108:data<=16'd13537;
      106109:data<=16'd14330;
      106110:data<=16'd14378;
      106111:data<=16'd14005;
      106112:data<=16'd13577;
      106113:data<=16'd12941;
      106114:data<=16'd12251;
      106115:data<=16'd12483;
      106116:data<=16'd13612;
      106117:data<=16'd13421;
      106118:data<=16'd12225;
      106119:data<=16'd12031;
      106120:data<=16'd12057;
      106121:data<=16'd11993;
      106122:data<=16'd12478;
      106123:data<=16'd12634;
      106124:data<=16'd12202;
      106125:data<=16'd11773;
      106126:data<=16'd11395;
      106127:data<=16'd10722;
      106128:data<=16'd10336;
      106129:data<=16'd11301;
      106130:data<=16'd11835;
      106131:data<=16'd10839;
      106132:data<=16'd10564;
      106133:data<=16'd10408;
      106134:data<=16'd9706;
      106135:data<=16'd11054;
      106136:data<=16'd12989;
      106137:data<=16'd12660;
      106138:data<=16'd11817;
      106139:data<=16'd11767;
      106140:data<=16'd11449;
      106141:data<=16'd11010;
      106142:data<=16'd11550;
      106143:data<=16'd12060;
      106144:data<=16'd11370;
      106145:data<=16'd10981;
      106146:data<=16'd10457;
      106147:data<=16'd9230;
      106148:data<=16'd9929;
      106149:data<=16'd9934;
      106150:data<=16'd6443;
      106151:data<=16'd4608;
      106152:data<=16'd5307;
      106153:data<=16'd4981;
      106154:data<=16'd4472;
      106155:data<=16'd3949;
      106156:data<=16'd3338;
      106157:data<=16'd3656;
      106158:data<=16'd3521;
      106159:data<=16'd3236;
      106160:data<=16'd3538;
      106161:data<=16'd2598;
      106162:data<=16'd908;
      106163:data<=16'd105;
      106164:data<=-16'd167;
      106165:data<=-16'd573;
      106166:data<=-16'd1013;
      106167:data<=-16'd834;
      106168:data<=-16'd1005;
      106169:data<=-16'd2537;
      106170:data<=-16'd3563;
      106171:data<=-16'd3212;
      106172:data<=-16'd2754;
      106173:data<=-16'd2757;
      106174:data<=-16'd3409;
      106175:data<=-16'd4587;
      106176:data<=-16'd5406;
      106177:data<=-16'd5266;
      106178:data<=-16'd4984;
      106179:data<=-16'd5292;
      106180:data<=-16'd5333;
      106181:data<=-16'd5509;
      106182:data<=-16'd6570;
      106183:data<=-16'd7127;
      106184:data<=-16'd7141;
      106185:data<=-16'd7289;
      106186:data<=-16'd7063;
      106187:data<=-16'd6771;
      106188:data<=-16'd6918;
      106189:data<=-16'd7935;
      106190:data<=-16'd8739;
      106191:data<=-16'd8035;
      106192:data<=-16'd8037;
      106193:data<=-16'd7606;
      106194:data<=-16'd4484;
      106195:data<=-16'd3571;
      106196:data<=-16'd5098;
      106197:data<=-16'd4454;
      106198:data<=-16'd4197;
      106199:data<=-16'd5222;
      106200:data<=-16'd4764;
      106201:data<=-16'd5049;
      106202:data<=-16'd7448;
      106203:data<=-16'd9048;
      106204:data<=-16'd8637;
      106205:data<=-16'd8299;
      106206:data<=-16'd8470;
      106207:data<=-16'd7483;
      106208:data<=-16'd7470;
      106209:data<=-16'd9280;
      106210:data<=-16'd9386;
      106211:data<=-16'd8690;
      106212:data<=-16'd8807;
      106213:data<=-16'd8354;
      106214:data<=-16'd8395;
      106215:data<=-16'd9083;
      106216:data<=-16'd9403;
      106217:data<=-16'd9559;
      106218:data<=-16'd9015;
      106219:data<=-16'd8611;
      106220:data<=-16'd8484;
      106221:data<=-16'd8129;
      106222:data<=-16'd9179;
      106223:data<=-16'd9902;
      106224:data<=-16'd8998;
      106225:data<=-16'd9068;
      106226:data<=-16'd8975;
      106227:data<=-16'd8015;
      106228:data<=-16'd8445;
      106229:data<=-16'd9165;
      106230:data<=-16'd8916;
      106231:data<=-16'd8502;
      106232:data<=-16'd8310;
      106233:data<=-16'd8035;
      106234:data<=-16'd7612;
      106235:data<=-16'd8395;
      106236:data<=-16'd9335;
      106237:data<=-16'd8795;
      106238:data<=-16'd9925;
      106239:data<=-16'd12568;
      106240:data<=-16'd12666;
      106241:data<=-16'd11999;
      106242:data<=-16'd13098;
      106243:data<=-16'd13509;
      106244:data<=-16'd12196;
      106245:data<=-16'd11620;
      106246:data<=-16'd11617;
      106247:data<=-16'd10360;
      106248:data<=-16'd10373;
      106249:data<=-16'd11997;
      106250:data<=-16'd11332;
      106251:data<=-16'd10252;
      106252:data<=-16'd10669;
      106253:data<=-16'd9699;
      106254:data<=-16'd8813;
      106255:data<=-16'd9911;
      106256:data<=-16'd10307;
      106257:data<=-16'd9309;
      106258:data<=-16'd8733;
      106259:data<=-16'd8746;
      106260:data<=-16'd8005;
      106261:data<=-16'd7195;
      106262:data<=-16'd7195;
      106263:data<=-16'd6370;
      106264:data<=-16'd5759;
      106265:data<=-16'd6029;
      106266:data<=-16'd5150;
      106267:data<=-16'd4734;
      106268:data<=-16'd3788;
      106269:data<=-16'd459;
      106270:data<=16'd684;
      106271:data<=16'd456;
      106272:data<=16'd1562;
      106273:data<=16'd1125;
      106274:data<=16'd1372;
      106275:data<=16'd3366;
      106276:data<=16'd3750;
      106277:data<=16'd3993;
      106278:data<=16'd4246;
      106279:data<=16'd4065;
      106280:data<=16'd4645;
      106281:data<=16'd4557;
      106282:data<=16'd6576;
      106283:data<=16'd10939;
      106284:data<=16'd11358;
      106285:data<=16'd10126;
      106286:data<=16'd10725;
      106287:data<=16'd10571;
      106288:data<=16'd11015;
      106289:data<=16'd12164;
      106290:data<=16'd11909;
      106291:data<=16'd11838;
      106292:data<=16'd11721;
      106293:data<=16'd11003;
      106294:data<=16'd11230;
      106295:data<=16'd11906;
      106296:data<=16'd12066;
      106297:data<=16'd11828;
      106298:data<=16'd11731;
      106299:data<=16'd11614;
      106300:data<=16'd10859;
      106301:data<=16'd11018;
      106302:data<=16'd12117;
      106303:data<=16'd12098;
      106304:data<=16'd11784;
      106305:data<=16'd11562;
      106306:data<=16'd10704;
      106307:data<=16'd10578;
      106308:data<=16'd11341;
      106309:data<=16'd11634;
      106310:data<=16'd11383;
      106311:data<=16'd11414;
      106312:data<=16'd11398;
      106313:data<=16'd10088;
      106314:data<=16'd9482;
      106315:data<=16'd11217;
      106316:data<=16'd11981;
      106317:data<=16'd11198;
      106318:data<=16'd11151;
      106319:data<=16'd10693;
      106320:data<=16'd9547;
      106321:data<=16'd9790;
      106322:data<=16'd11227;
      106323:data<=16'd11417;
      106324:data<=16'd10108;
      106325:data<=16'd9905;
      106326:data<=16'd9639;
      106327:data<=16'd7206;
      106328:data<=16'd5940;
      106329:data<=16'd6240;
      106330:data<=16'd5497;
      106331:data<=16'd5260;
      106332:data<=16'd5377;
      106333:data<=16'd4690;
      106334:data<=16'd4977;
      106335:data<=16'd5470;
      106336:data<=16'd4740;
      106337:data<=16'd3874;
      106338:data<=16'd3463;
      106339:data<=16'd3425;
      106340:data<=16'd3422;
      106341:data<=16'd3777;
      106342:data<=16'd4698;
      106343:data<=16'd4660;
      106344:data<=16'd3982;
      106345:data<=16'd4061;
      106346:data<=16'd4225;
      106347:data<=16'd4244;
      106348:data<=16'd4602;
      106349:data<=16'd5183;
      106350:data<=16'd5357;
      106351:data<=16'd4796;
      106352:data<=16'd4431;
      106353:data<=16'd4240;
      106354:data<=16'd4347;
      106355:data<=16'd5488;
      106356:data<=16'd5483;
      106357:data<=16'd4434;
      106358:data<=16'd4852;
      106359:data<=16'd4758;
      106360:data<=16'd3829;
      106361:data<=16'd4399;
      106362:data<=16'd5096;
      106363:data<=16'd5151;
      106364:data<=16'd5093;
      106365:data<=16'd4716;
      106366:data<=16'd4605;
      106367:data<=16'd4199;
      106368:data<=16'd3724;
      106369:data<=16'd3756;
      106370:data<=16'd2986;
      106371:data<=16'd3624;
      106372:data<=16'd6575;
      106373:data<=16'd7121;
      106374:data<=16'd5351;
      106375:data<=16'd4396;
      106376:data<=16'd3504;
      106377:data<=16'd2634;
      106378:data<=16'd2411;
      106379:data<=16'd2282;
      106380:data<=16'd2105;
      106381:data<=16'd1157;
      106382:data<=-16'd388;
      106383:data<=-16'd1005;
      106384:data<=-16'd925;
      106385:data<=-16'd1113;
      106386:data<=-16'd1374;
      106387:data<=-16'd1688;
      106388:data<=-16'd2573;
      106389:data<=-16'd3709;
      106390:data<=-16'd4244;
      106391:data<=-16'd4226;
      106392:data<=-16'd4029;
      106393:data<=-16'd3877;
      106394:data<=-16'd4349;
      106395:data<=-16'd5453;
      106396:data<=-16'd6081;
      106397:data<=-16'd5714;
      106398:data<=-16'd5606;
      106399:data<=-16'd5927;
      106400:data<=-16'd5629;
      106401:data<=-16'd6197;
      106402:data<=-16'd7285;
      106403:data<=-16'd6137;
      106404:data<=-16'd5438;
      106405:data<=-16'd6488;
      106406:data<=-16'd5758;
      106407:data<=-16'd5272;
      106408:data<=-16'd6748;
      106409:data<=-16'd7191;
      106410:data<=-16'd7295;
      106411:data<=-16'd7363;
      106412:data<=-16'd6385;
      106413:data<=-16'd6287;
      106414:data<=-16'd6953;
      106415:data<=-16'd8469;
      106416:data<=-16'd11335;
      106417:data<=-16'd12472;
      106418:data<=-16'd11994;
      106419:data<=-16'd11741;
      106420:data<=-16'd11412;
      106421:data<=-16'd12489;
      106422:data<=-16'd13567;
      106423:data<=-16'd12577;
      106424:data<=-16'd12263;
      106425:data<=-16'd12229;
      106426:data<=-16'd11323;
      106427:data<=-16'd11925;
      106428:data<=-16'd12948;
      106429:data<=-16'd12790;
      106430:data<=-16'd12413;
      106431:data<=-16'd11721;
      106432:data<=-16'd11141;
      106433:data<=-16'd11101;
      106434:data<=-16'd11345;
      106435:data<=-16'd11829;
      106436:data<=-16'd11624;
      106437:data<=-16'd11179;
      106438:data<=-16'd11191;
      106439:data<=-16'd10677;
      106440:data<=-16'd10419;
      106441:data<=-16'd11082;
      106442:data<=-16'd11406;
      106443:data<=-16'd11101;
      106444:data<=-16'd10637;
      106445:data<=-16'd10336;
      106446:data<=-16'd9705;
      106447:data<=-16'd9274;
      106448:data<=-16'd10517;
      106449:data<=-16'd11085;
      106450:data<=-16'd9938;
      106451:data<=-16'd9768;
      106452:data<=-16'd9447;
      106453:data<=-16'd8511;
      106454:data<=-16'd9085;
      106455:data<=-16'd9922;
      106456:data<=-16'd10238;
      106457:data<=-16'd9923;
      106458:data<=-16'd8812;
      106459:data<=-16'd8610;
      106460:data<=-16'd7558;
      106461:data<=-16'd5209;
      106462:data<=-16'd5059;
      106463:data<=-16'd5184;
      106464:data<=-16'd4225;
      106465:data<=-16'd4231;
      106466:data<=-16'd3865;
      106467:data<=-16'd4091;
      106468:data<=-16'd5783;
      106469:data<=-16'd5709;
      106470:data<=-16'd4778;
      106471:data<=-16'd4538;
      106472:data<=-16'd4073;
      106473:data<=-16'd4153;
      106474:data<=-16'd3842;
      106475:data<=-16'd3074;
      106476:data<=-16'd3604;
      106477:data<=-16'd3456;
      106478:data<=-16'd2513;
      106479:data<=-16'd2620;
      106480:data<=-16'd1820;
      106481:data<=-16'd438;
      106482:data<=-16'd417;
      106483:data<=-16'd97;
      106484:data<=16'd585;
      106485:data<=16'd497;
      106486:data<=16'd875;
      106487:data<=16'd1698;
      106488:data<=16'd2288;
      106489:data<=16'd3028;
      106490:data<=16'd3262;
      106491:data<=16'd3033;
      106492:data<=16'd3087;
      106493:data<=16'd3153;
      106494:data<=16'd3947;
      106495:data<=16'd5181;
      106496:data<=16'd5330;
      106497:data<=16'd5441;
      106498:data<=16'd5547;
      106499:data<=16'd4936;
      106500:data<=16'd5548;
      106501:data<=16'd6531;
      106502:data<=16'd6570;
      106503:data<=16'd7197;
      106504:data<=16'd6276;
      106505:data<=16'd3068;
      106506:data<=16'd1780;
      106507:data<=16'd2695;
      106508:data<=16'd3829;
      106509:data<=16'd4584;
      106510:data<=16'd4269;
      106511:data<=16'd4131;
      106512:data<=16'd4443;
      106513:data<=16'd4244;
      106514:data<=16'd4952;
      106515:data<=16'd5965;
      106516:data<=16'd5671;
      106517:data<=16'd5677;
      106518:data<=16'd6028;
      106519:data<=16'd5251;
      106520:data<=16'd4884;
      106521:data<=16'd6264;
      106522:data<=16'd7535;
      106523:data<=16'd7680;
      106524:data<=16'd7700;
      106525:data<=16'd6865;
      106526:data<=16'd5489;
      106527:data<=16'd6451;
      106528:data<=16'd8711;
      106529:data<=16'd9433;
      106530:data<=16'd9007;
      106531:data<=16'd8090;
      106532:data<=16'd7450;
      106533:data<=16'd7830;
      106534:data<=16'd8624;
      106535:data<=16'd9374;
      106536:data<=16'd9226;
      106537:data<=16'd8640;
      106538:data<=16'd8671;
      106539:data<=16'd7747;
      106540:data<=16'd7236;
      106541:data<=16'd9031;
      106542:data<=16'd9641;
      106543:data<=16'd8739;
      106544:data<=16'd8661;
      106545:data<=16'd8155;
      106546:data<=16'd7629;
      106547:data<=16'd8100;
      106548:data<=16'd8828;
      106549:data<=16'd10313;
      106550:data<=16'd11890;
      106551:data<=16'd12407;
      106552:data<=16'd12090;
      106553:data<=16'd11301;
      106554:data<=16'd11465;
      106555:data<=16'd12184;
      106556:data<=16'd11799;
      106557:data<=16'd11505;
      106558:data<=16'd11113;
      106559:data<=16'd9767;
      106560:data<=16'd9514;
      106561:data<=16'd10363;
      106562:data<=16'd10592;
      106563:data<=16'd10255;
      106564:data<=16'd9797;
      106565:data<=16'd9453;
      106566:data<=16'd9016;
      106567:data<=16'd8849;
      106568:data<=16'd9474;
      106569:data<=16'd9565;
      106570:data<=16'd8968;
      106571:data<=16'd8575;
      106572:data<=16'd8003;
      106573:data<=16'd8087;
      106574:data<=16'd9024;
      106575:data<=16'd9306;
      106576:data<=16'd9128;
      106577:data<=16'd8658;
      106578:data<=16'd7444;
      106579:data<=16'd6390;
      106580:data<=16'd6244;
      106581:data<=16'd6476;
      106582:data<=16'd6159;
      106583:data<=16'd5651;
      106584:data<=16'd5350;
      106585:data<=16'd4640;
      106586:data<=16'd4335;
      106587:data<=16'd3826;
      106588:data<=16'd1977;
      106589:data<=16'd1433;
      106590:data<=16'd1524;
      106591:data<=16'd537;
      106592:data<=16'd949;
      106593:data<=-16'd282;
      106594:data<=-16'd4745;
      106595:data<=-16'd6097;
      106596:data<=-16'd5383;
      106597:data<=-16'd6213;
      106598:data<=-16'd6096;
      106599:data<=-16'd5841;
      106600:data<=-16'd6539;
      106601:data<=-16'd7100;
      106602:data<=-16'd8147;
      106603:data<=-16'd8231;
      106604:data<=-16'd7454;
      106605:data<=-16'd7785;
      106606:data<=-16'd7696;
      106607:data<=-16'd7680;
      106608:data<=-16'd8851;
      106609:data<=-16'd8922;
      106610:data<=-16'd8241;
      106611:data<=-16'd8272;
      106612:data<=-16'd8066;
      106613:data<=-16'd7808;
      106614:data<=-16'd8522;
      106615:data<=-16'd9309;
      106616:data<=-16'd9068;
      106617:data<=-16'd8846;
      106618:data<=-16'd8652;
      106619:data<=-16'd7733;
      106620:data<=-16'd8307;
      106621:data<=-16'd9729;
      106622:data<=-16'd9180;
      106623:data<=-16'd8593;
      106624:data<=-16'd8511;
      106625:data<=-16'd7846;
      106626:data<=-16'd8247;
      106627:data<=-16'd9044;
      106628:data<=-16'd9229;
      106629:data<=-16'd9327;
      106630:data<=-16'd8954;
      106631:data<=-16'd8960;
      106632:data<=-16'd8825;
      106633:data<=-16'd8252;
      106634:data<=-16'd9447;
      106635:data<=-16'd10662;
      106636:data<=-16'd10214;
      106637:data<=-16'd9081;
      106638:data<=-16'd6378;
      106639:data<=-16'd4206;
      106640:data<=-16'd4984;
      106641:data<=-16'd6475;
      106642:data<=-16'd6907;
      106643:data<=-16'd5961;
      106644:data<=-16'd5382;
      106645:data<=-16'd5914;
      106646:data<=-16'd5269;
      106647:data<=-16'd5436;
      106648:data<=-16'd6702;
      106649:data<=-16'd5661;
      106650:data<=-16'd5316;
      106651:data<=-16'd6307;
      106652:data<=-16'd5409;
      106653:data<=-16'd5422;
      106654:data<=-16'd6893;
      106655:data<=-16'd7172;
      106656:data<=-16'd7021;
      106657:data<=-16'd6611;
      106658:data<=-16'd5912;
      106659:data<=-16'd5733;
      106660:data<=-16'd6190;
      106661:data<=-16'd6678;
      106662:data<=-16'd6070;
      106663:data<=-16'd5930;
      106664:data<=-16'd6672;
      106665:data<=-16'd5705;
      106666:data<=-16'd4824;
      106667:data<=-16'd5777;
      106668:data<=-16'd6623;
      106669:data<=-16'd6910;
      106670:data<=-16'd6549;
      106671:data<=-16'd6203;
      106672:data<=-16'd6096;
      106673:data<=-16'd5416;
      106674:data<=-16'd6185;
      106675:data<=-16'd7131;
      106676:data<=-16'd5946;
      106677:data<=-16'd5709;
      106678:data<=-16'd5668;
      106679:data<=-16'd4743;
      106680:data<=-16'd5697;
      106681:data<=-16'd6223;
      106682:data<=-16'd6352;
      106683:data<=-16'd8874;
      106684:data<=-16'd9855;
      106685:data<=-16'd8539;
      106686:data<=-16'd8399;
      106687:data<=-16'd8464;
      106688:data<=-16'd7914;
      106689:data<=-16'd7356;
      106690:data<=-16'd6604;
      106691:data<=-16'd5964;
      106692:data<=-16'd5498;
      106693:data<=-16'd4716;
      106694:data<=-16'd3121;
      106695:data<=-16'd1765;
      106696:data<=-16'd1621;
      106697:data<=-16'd1413;
      106698:data<=-16'd1592;
      106699:data<=-16'd2188;
      106700:data<=-16'd785;
      106701:data<=16'd1160;
      106702:data<=16'd1612;
      106703:data<=16'd1917;
      106704:data<=16'd2017;
      106705:data<=16'd1694;
      106706:data<=16'd2267;
      106707:data<=16'd3664;
      106708:data<=16'd4399;
      106709:data<=16'd4071;
      106710:data<=16'd4208;
      106711:data<=16'd4669;
      106712:data<=16'd4338;
      106713:data<=16'd4833;
      106714:data<=16'd6258;
      106715:data<=16'd6651;
      106716:data<=16'd6469;
      106717:data<=16'd6434;
      106718:data<=16'd5890;
      106719:data<=16'd5198;
      106720:data<=16'd6250;
      106721:data<=16'd8087;
      106722:data<=16'd7498;
      106723:data<=16'd6956;
      106724:data<=16'd7931;
      106725:data<=16'd6757;
      106726:data<=16'd7145;
      106727:data<=16'd11438;
      106728:data<=16'd12774;
      106729:data<=16'd11788;
      106730:data<=16'd12314;
      106731:data<=16'd11984;
      106732:data<=16'd11311;
      106733:data<=16'd11509;
      106734:data<=16'd11794;
      106735:data<=16'd12222;
      106736:data<=16'd11602;
      106737:data<=16'd10925;
      106738:data<=16'd11197;
      106739:data<=16'd10672;
      106740:data<=16'd10840;
      106741:data<=16'd11941;
      106742:data<=16'd11549;
      106743:data<=16'd10921;
      106744:data<=16'd10909;
      106745:data<=16'd10592;
      106746:data<=16'd10249;
      106747:data<=16'd10566;
      106748:data<=16'd11577;
      106749:data<=16'd11345;
      106750:data<=16'd10152;
      106751:data<=16'd9837;
      106752:data<=16'd8883;
      106753:data<=16'd8771;
      106754:data<=16'd10734;
      106755:data<=16'd10520;
      106756:data<=16'd9136;
      106757:data<=16'd9210;
      106758:data<=16'd8830;
      106759:data<=16'd9063;
      106760:data<=16'd10103;
      106761:data<=16'd9741;
      106762:data<=16'd8987;
      106763:data<=16'd8634;
      106764:data<=16'd8443;
      106765:data<=16'd7978;
      106766:data<=16'd7650;
      106767:data<=16'd8877;
      106768:data<=16'd8866;
      106769:data<=16'd7470;
      106770:data<=16'd8129;
      106771:data<=16'd6561;
      106772:data<=16'd2238;
      106773:data<=16'd1999;
      106774:data<=16'd3777;
      106775:data<=16'd3756;
      106776:data<=16'd3576;
      106777:data<=16'd3055;
      106778:data<=16'd2314;
      106779:data<=16'd2055;
      106780:data<=16'd2605;
      106781:data<=16'd4138;
      106782:data<=16'd4102;
      106783:data<=16'd3095;
      106784:data<=16'd3260;
      106785:data<=16'd2570;
      106786:data<=16'd2511;
      106787:data<=16'd4366;
      106788:data<=16'd4309;
      106789:data<=16'd3383;
      106790:data<=16'd3874;
      106791:data<=16'd3941;
      106792:data<=16'd3745;
      106793:data<=16'd3506;
      106794:data<=16'd2643;
      106795:data<=16'd2094;
      106796:data<=16'd1548;
      106797:data<=16'd1218;
      106798:data<=16'd1844;
      106799:data<=16'd1524;
      106800:data<=-16'd297;
      106801:data<=-16'd1475;
      106802:data<=-16'd1545;
      106803:data<=-16'd1804;
      106804:data<=-16'd2446;
      106805:data<=-16'd2811;
      106806:data<=-16'd3218;
      106807:data<=-16'd3947;
      106808:data<=-16'd4508;
      106809:data<=-16'd4723;
      106810:data<=-16'd4664;
      106811:data<=-16'd4532;
      106812:data<=-16'd4340;
      106813:data<=-16'd4877;
      106814:data<=-16'd6702;
      106815:data<=-16'd6147;
      106816:data<=-16'd2476;
      106817:data<=-16'd1545;
      106818:data<=-16'd2863;
      106819:data<=-16'd2645;
      106820:data<=-16'd3366;
      106821:data<=-16'd4640;
      106822:data<=-16'd4363;
      106823:data<=-16'd4793;
      106824:data<=-16'd5025;
      106825:data<=-16'd4009;
      106826:data<=-16'd4730;
      106827:data<=-16'd6479;
      106828:data<=-16'd6683;
      106829:data<=-16'd6117;
      106830:data<=-16'd5926;
      106831:data<=-16'd5926;
      106832:data<=-16'd6135;
      106833:data<=-16'd7165;
      106834:data<=-16'd8228;
      106835:data<=-16'd8150;
      106836:data<=-16'd7873;
      106837:data<=-16'd7682;
      106838:data<=-16'd7185;
      106839:data<=-16'd7548;
      106840:data<=-16'd8577;
      106841:data<=-16'd8624;
      106842:data<=-16'd8015;
      106843:data<=-16'd8244;
      106844:data<=-16'd8469;
      106845:data<=-16'd7450;
      106846:data<=-16'd7732;
      106847:data<=-16'd9659;
      106848:data<=-16'd9624;
      106849:data<=-16'd8742;
      106850:data<=-16'd8777;
      106851:data<=-16'd8079;
      106852:data<=-16'd8008;
      106853:data<=-16'd9427;
      106854:data<=-16'd10266;
      106855:data<=-16'd10175;
      106856:data<=-16'd9738;
      106857:data<=-16'd9336;
      106858:data<=-16'd8269;
      106859:data<=-16'd7756;
      106860:data<=-16'd11118;
      106861:data<=-16'd14266;
      106862:data<=-16'd13256;
      106863:data<=-16'd12801;
      106864:data<=-16'd13107;
      106865:data<=-16'd11847;
      106866:data<=-16'd11764;
      106867:data<=-16'd12434;
      106868:data<=-16'd12275;
      106869:data<=-16'd12013;
      106870:data<=-16'd11315;
      106871:data<=-16'd11060;
      106872:data<=-16'd11559;
      106873:data<=-16'd11702;
      106874:data<=-16'd11744;
      106875:data<=-16'd11397;
      106876:data<=-16'd10663;
      106877:data<=-16'd10067;
      106878:data<=-16'd9461;
      106879:data<=-16'd9492;
      106880:data<=-16'd9972;
      106881:data<=-16'd10025;
      106882:data<=-16'd9621;
      106883:data<=-16'd8995;
      106884:data<=-16'd8740;
      106885:data<=-16'd8490;
      106886:data<=-16'd8769;
      106887:data<=-16'd9928;
      106888:data<=-16'd9397;
      106889:data<=-16'd8631;
      106890:data<=-16'd9180;
      106891:data<=-16'd7721;
      106892:data<=-16'd6687;
      106893:data<=-16'd8261;
      106894:data<=-16'd8520;
      106895:data<=-16'd8050;
      106896:data<=-16'd7765;
      106897:data<=-16'd6836;
      106898:data<=-16'd6843;
      106899:data<=-16'd6551;
      106900:data<=-16'd5741;
      106901:data<=-16'd5680;
      106902:data<=-16'd5181;
      106903:data<=-16'd5163;
      106904:data<=-16'd4219;
      106905:data<=-16'd796;
      106906:data<=16'd1169;
      106907:data<=16'd2005;
      106908:data<=16'd3054;
      106909:data<=16'd2547;
      106910:data<=16'd2547;
      106911:data<=16'd3118;
      106912:data<=16'd3046;
      106913:data<=16'd4061;
      106914:data<=16'd4813;
      106915:data<=16'd4955;
      106916:data<=16'd5527;
      106917:data<=16'd4898;
      106918:data<=16'd4261;
      106919:data<=16'd5057;
      106920:data<=16'd6122;
      106921:data<=16'd6836;
      106922:data<=16'd6598;
      106923:data<=16'd6246;
      106924:data<=16'd6061;
      106925:data<=16'd5395;
      106926:data<=16'd6187;
      106927:data<=16'd7820;
      106928:data<=16'd8076;
      106929:data<=16'd7896;
      106930:data<=16'd7635;
      106931:data<=16'd7577;
      106932:data<=16'd8181;
      106933:data<=16'd8771;
      106934:data<=16'd9232;
      106935:data<=16'd8816;
      106936:data<=16'd8408;
      106937:data<=16'd8869;
      106938:data<=16'd7979;
      106939:data<=16'd7626;
      106940:data<=16'd9488;
      106941:data<=16'd9705;
      106942:data<=16'd8789;
      106943:data<=16'd8954;
      106944:data<=16'd8443;
      106945:data<=16'd7899;
      106946:data<=16'd9229;
      106947:data<=16'd10833;
      106948:data<=16'd9829;
      106949:data<=16'd6890;
      106950:data<=16'd5218;
      106951:data<=16'd4804;
      106952:data<=16'd5012;
      106953:data<=16'd6179;
      106954:data<=16'd6739;
      106955:data<=16'd6783;
      106956:data<=16'd6940;
      106957:data<=16'd5905;
      106958:data<=16'd4394;
      106959:data<=16'd4783;
      106960:data<=16'd7482;
      106961:data<=16'd8693;
      106962:data<=16'd6687;
      106963:data<=16'd6034;
      106964:data<=16'd6479;
      106965:data<=16'd5950;
      106966:data<=16'd7248;
      106967:data<=16'd7935;
      106968:data<=16'd7098;
      106969:data<=16'd8272;
      106970:data<=16'd7890;
      106971:data<=16'd6067;
      106972:data<=16'd7056;
      106973:data<=16'd7850;
      106974:data<=16'd7448;
      106975:data<=16'd7256;
      106976:data<=16'd6884;
      106977:data<=16'd7106;
      106978:data<=16'd6836;
      106979:data<=16'd7244;
      106980:data<=16'd9288;
      106981:data<=16'd8698;
      106982:data<=16'd6837;
      106983:data<=16'd6725;
      106984:data<=16'd6648;
      106985:data<=16'd7084;
      106986:data<=16'd7379;
      106987:data<=16'd7098;
      106988:data<=16'd7727;
      106989:data<=16'd7316;
      106990:data<=16'd6587;
      106991:data<=16'd6680;
      106992:data<=16'd6228;
      106993:data<=16'd8304;
      106994:data<=16'd11512;
      106995:data<=16'd11253;
      106996:data<=16'd10684;
      106997:data<=16'd10675;
      106998:data<=16'd9456;
      106999:data<=16'd9603;
      107000:data<=16'd10881;
      107001:data<=16'd11154;
      107002:data<=16'd10634;
      107003:data<=16'd9758;
      107004:data<=16'd9036;
      107005:data<=16'd8721;
      107006:data<=16'd8822;
      107007:data<=16'd8319;
      107008:data<=16'd6716;
      107009:data<=16'd6250;
      107010:data<=16'd6686;
      107011:data<=16'd6399;
      107012:data<=16'd5879;
      107013:data<=16'd4426;
      107014:data<=16'd3102;
      107015:data<=16'd3312;
      107016:data<=16'd2936;
      107017:data<=16'd2587;
      107018:data<=16'd2846;
      107019:data<=16'd1486;
      107020:data<=-16'd30;
      107021:data<=-16'd428;
      107022:data<=-16'd795;
      107023:data<=-16'd660;
      107024:data<=-16'd494;
      107025:data<=-16'd1149;
      107026:data<=-16'd1989;
      107027:data<=-16'd2329;
      107028:data<=-16'd2312;
      107029:data<=-16'd3096;
      107030:data<=-16'd3680;
      107031:data<=-16'd3110;
      107032:data<=-16'd3747;
      107033:data<=-16'd5104;
      107034:data<=-16'd5386;
      107035:data<=-16'd5562;
      107036:data<=-16'd5527;
      107037:data<=-16'd6176;
      107038:data<=-16'd8120;
      107039:data<=-16'd9339;
      107040:data<=-16'd10696;
      107041:data<=-16'd11887;
      107042:data<=-16'd10828;
      107043:data<=-16'd10210;
      107044:data<=-16'd10336;
      107045:data<=-16'd9357;
      107046:data<=-16'd9790;
      107047:data<=-16'd10792;
      107048:data<=-16'd9861;
      107049:data<=-16'd9445;
      107050:data<=-16'd9782;
      107051:data<=-16'd9088;
      107052:data<=-16'd9147;
      107053:data<=-16'd10489;
      107054:data<=-16'd10472;
      107055:data<=-16'd9092;
      107056:data<=-16'd8683;
      107057:data<=-16'd8681;
      107058:data<=-16'd8298;
      107059:data<=-16'd9109;
      107060:data<=-16'd10342;
      107061:data<=-16'd10566;
      107062:data<=-16'd10314;
      107063:data<=-16'd9247;
      107064:data<=-16'd8536;
      107065:data<=-16'd9456;
      107066:data<=-16'd10056;
      107067:data<=-16'd10129;
      107068:data<=-16'd10152;
      107069:data<=-16'd9391;
      107070:data<=-16'd8984;
      107071:data<=-16'd8862;
      107072:data<=-16'd8900;
      107073:data<=-16'd10123;
      107074:data<=-16'd10175;
      107075:data<=-16'd8857;
      107076:data<=-16'd8869;
      107077:data<=-16'd9054;
      107078:data<=-16'd8783;
      107079:data<=-16'd8994;
      107080:data<=-16'd9356;
      107081:data<=-16'd9354;
      107082:data<=-16'd6865;
      107083:data<=-16'd3410;
      107084:data<=-16'd3576;
      107085:data<=-16'd4851;
      107086:data<=-16'd4610;
      107087:data<=-16'd4851;
      107088:data<=-16'd4981;
      107089:data<=-16'd5068;
      107090:data<=-16'd5259;
      107091:data<=-16'd4214;
      107092:data<=-16'd4479;
      107093:data<=-16'd5626;
      107094:data<=-16'd4475;
      107095:data<=-16'd4129;
      107096:data<=-16'd5424;
      107097:data<=-16'd5083;
      107098:data<=-16'd4551;
      107099:data<=-16'd5333;
      107100:data<=-16'd5970;
      107101:data<=-16'd5849;
      107102:data<=-16'd5272;
      107103:data<=-16'd4681;
      107104:data<=-16'd3947;
      107105:data<=-16'd4115;
      107106:data<=-16'd5811;
      107107:data<=-16'd6075;
      107108:data<=-16'd5096;
      107109:data<=-16'd5506;
      107110:data<=-16'd5371;
      107111:data<=-16'd4334;
      107112:data<=-16'd4126;
      107113:data<=-16'd3733;
      107114:data<=-16'd3580;
      107115:data<=-16'd3783;
      107116:data<=-16'd3154;
      107117:data<=-16'd2963;
      107118:data<=-16'd2481;
      107119:data<=-16'd419;
      107120:data<=16'd755;
      107121:data<=16'd458;
      107122:data<=16'd92;
      107123:data<=-16'd517;
      107124:data<=-16'd755;
      107125:data<=16'd534;
      107126:data<=16'd1513;
      107127:data<=-16'd179;
      107128:data<=-16'd1676;
      107129:data<=-16'd1134;
      107130:data<=-16'd1732;
      107131:data<=-16'd1668;
      107132:data<=16'd610;
      107133:data<=16'd1556;
      107134:data<=16'd2428;
      107135:data<=16'd2614;
      107136:data<=16'd1228;
      107137:data<=16'd2279;
      107138:data<=16'd425;
      107139:data<=-16'd4543;
      107140:data<=-16'd4676;
      107141:data<=-16'd4223;
      107142:data<=16'd3779;
      107143:data<=16'd21062;
      107144:data<=16'd17946;
      107145:data<=-16'd1300;
      107146:data<=-16'd5891;
      107147:data<=-16'd4299;
      107148:data<=-16'd5571;
      107149:data<=-16'd3231;
      107150:data<=-16'd2987;
      107151:data<=-16'd3122;
      107152:data<=-16'd2026;
      107153:data<=-16'd3034;
      107154:data<=-16'd611;
      107155:data<=-16'd3726;
      107156:data<=-16'd16222;
      107157:data<=-16'd16130;
      107158:data<=-16'd2581;
      107159:data<=16'd5736;
      107160:data<=16'd6537;
      107161:data<=16'd5224;
      107162:data<=16'd4581;
      107163:data<=16'd4511;
      107164:data<=16'd4276;
      107165:data<=16'd5195;
      107166:data<=16'd5680;
      107167:data<=16'd5548;
      107168:data<=16'd6052;
      107169:data<=16'd5617;
      107170:data<=16'd6062;
      107171:data<=16'd7659;
      107172:data<=16'd7160;
      107173:data<=16'd6100;
      107174:data<=16'd6399;
      107175:data<=16'd7480;
      107176:data<=16'd8085;
      107177:data<=16'd7156;
      107178:data<=16'd6256;
      107179:data<=16'd5679;
      107180:data<=16'd4840;
      107181:data<=16'd4637;
      107182:data<=16'd4726;
      107183:data<=16'd5137;
      107184:data<=16'd4708;
      107185:data<=16'd3077;
      107186:data<=16'd2916;
      107187:data<=16'd2670;
      107188:data<=16'd2088;
      107189:data<=16'd2541;
      107190:data<=16'd1319;
      107191:data<=16'd3245;
      107192:data<=16'd9953;
      107193:data<=16'd11653;
      107194:data<=16'd10097;
      107195:data<=16'd10395;
      107196:data<=16'd9169;
      107197:data<=16'd8219;
      107198:data<=16'd8152;
      107199:data<=16'd6969;
      107200:data<=16'd6751;
      107201:data<=16'd6209;
      107202:data<=16'd5479;
      107203:data<=16'd6484;
      107204:data<=16'd6481;
      107205:data<=16'd5507;
      107206:data<=16'd4983;
      107207:data<=16'd4687;
      107208:data<=16'd5389;
      107209:data<=16'd5500;
      107210:data<=16'd4168;
      107211:data<=16'd2613;
      107212:data<=16'd1410;
      107213:data<=16'd1918;
      107214:data<=16'd2684;
      107215:data<=16'd1166;
      107216:data<=-16'd1748;
      107217:data<=-16'd3797;
      107218:data<=-16'd2949;
      107219:data<=-16'd1877;
      107220:data<=-16'd3001;
      107221:data<=-16'd2669;
      107222:data<=-16'd1647;
      107223:data<=-16'd1917;
      107224:data<=-16'd1662;
      107225:data<=-16'd2984;
      107226:data<=-16'd4491;
      107227:data<=-16'd2855;
      107228:data<=-16'd2147;
      107229:data<=-16'd3175;
      107230:data<=-16'd3362;
      107231:data<=-16'd3065;
      107232:data<=-16'd2118;
      107233:data<=-16'd1751;
      107234:data<=-16'd2036;
      107235:data<=-16'd1691;
      107236:data<=-16'd2135;
      107237:data<=-16'd2740;
      107238:data<=-16'd3239;
      107239:data<=-16'd3714;
      107240:data<=-16'd2188;
      107241:data<=-16'd2253;
      107242:data<=-16'd4026;
      107243:data<=-16'd2810;
      107244:data<=-16'd4570;
      107245:data<=-16'd10310;
      107246:data<=-16'd10969;
      107247:data<=-16'd9479;
      107248:data<=-16'd10295;
      107249:data<=-16'd9567;
      107250:data<=-16'd8901;
      107251:data<=-16'd9970;
      107252:data<=-16'd9843;
      107253:data<=-16'd9421;
      107254:data<=-16'd9770;
      107255:data<=-16'd9461;
      107256:data<=-16'd8173;
      107257:data<=-16'd6513;
      107258:data<=-16'd6297;
      107259:data<=-16'd7007;
      107260:data<=-16'd5259;
      107261:data<=-16'd2549;
      107262:data<=-16'd1870;
      107263:data<=-16'd1794;
      107264:data<=-16'd1964;
      107265:data<=-16'd2623;
      107266:data<=-16'd2554;
      107267:data<=-16'd2626;
      107268:data<=-16'd2834;
      107269:data<=-16'd2322;
      107270:data<=-16'd2182;
      107271:data<=-16'd1800;
      107272:data<=-16'd1277;
      107273:data<=-16'd2052;
      107274:data<=-16'd2127;
      107275:data<=-16'd1021;
      107276:data<=-16'd726;
      107277:data<=-16'd1451;
      107278:data<=-16'd3247;
      107279:data<=-16'd4179;
      107280:data<=-16'd2869;
      107281:data<=-16'd2353;
      107282:data<=-16'd2431;
      107283:data<=-16'd1351;
      107284:data<=-16'd1410;
      107285:data<=-16'd1914;
      107286:data<=-16'd1189;
      107287:data<=-16'd1401;
      107288:data<=-16'd1624;
      107289:data<=-16'd587;
      107290:data<=-16'd1101;
      107291:data<=-16'd2096;
      107292:data<=-16'd1695;
      107293:data<=-16'd2270;
      107294:data<=-16'd2355;
      107295:data<=-16'd1519;
      107296:data<=-16'd2998;
      107297:data<=-16'd1195;
      107298:data<=16'd5835;
      107299:data<=16'd8170;
      107300:data<=16'd6391;
      107301:data<=16'd6733;
      107302:data<=16'd6737;
      107303:data<=16'd6191;
      107304:data<=16'd5162;
      107305:data<=16'd2024;
      107306:data<=16'd506;
      107307:data<=16'd819;
      107308:data<=16'd277;
      107309:data<=16'd252;
      107310:data<=16'd581;
      107311:data<=16'd688;
      107312:data<=16'd887;
      107313:data<=16'd810;
      107314:data<=16'd1163;
      107315:data<=16'd1266;
      107316:data<=16'd878;
      107317:data<=16'd566;
      107318:data<=-16'd644;
      107319:data<=-16'd836;
      107320:data<=16'd414;
      107321:data<=16'd126;
      107322:data<=-16'd494;
      107323:data<=-16'd247;
      107324:data<=-16'd71;
      107325:data<=16'd241;
      107326:data<=16'd94;
      107327:data<=-16'd173;
      107328:data<=16'd203;
      107329:data<=16'd823;
      107330:data<=16'd787;
      107331:data<=-16'd943;
      107332:data<=-16'd1448;
      107333:data<=-16'd8;
      107334:data<=-16'd449;
      107335:data<=-16'd608;
      107336:data<=16'd302;
      107337:data<=-16'd212;
      107338:data<=16'd540;
      107339:data<=16'd1043;
      107340:data<=-16'd409;
      107341:data<=-16'd234;
      107342:data<=16'd42;
      107343:data<=-16'd171;
      107344:data<=-16'd570;
      107345:data<=-16'd2572;
      107346:data<=-16'd1530;
      107347:data<=16'd459;
      107348:data<=-16'd1196;
      107349:data<=16'd176;
      107350:data<=16'd1847;
      107351:data<=-16'd2766;
      107352:data<=-16'd5812;
      107353:data<=-16'd4520;
      107354:data<=-16'd3548;
      107355:data<=-16'd2717;
      107356:data<=-16'd2638;
      107357:data<=-16'd3375;
      107358:data<=-16'd3040;
      107359:data<=-16'd2475;
      107360:data<=-16'd2535;
      107361:data<=-16'd2416;
      107362:data<=-16'd1867;
      107363:data<=-16'd1651;
      107364:data<=-16'd1325;
      107365:data<=-16'd522;
      107366:data<=-16'd978;
      107367:data<=-16'd1902;
      107368:data<=-16'd1905;
      107369:data<=-16'd1856;
      107370:data<=-16'd235;
      107371:data<=16'd2167;
      107372:data<=16'd2164;
      107373:data<=16'd1988;
      107374:data<=16'd2786;
      107375:data<=16'd2453;
      107376:data<=16'd2267;
      107377:data<=16'd3068;
      107378:data<=16'd3036;
      107379:data<=16'd2199;
      107380:data<=16'd2311;
      107381:data<=16'd3116;
      107382:data<=16'd3089;
      107383:data<=16'd3115;
      107384:data<=16'd3958;
      107385:data<=16'd4595;
      107386:data<=16'd4745;
      107387:data<=16'd4288;
      107388:data<=16'd4434;
      107389:data<=16'd5829;
      107390:data<=16'd5709;
      107391:data<=16'd4451;
      107392:data<=16'd4645;
      107393:data<=16'd4496;
      107394:data<=16'd2352;
      107395:data<=16'd127;
      107396:data<=16'd182;
      107397:data<=16'd2076;
      107398:data<=16'd2842;
      107399:data<=16'd2079;
      107400:data<=16'd2190;
      107401:data<=16'd3306;
      107402:data<=16'd3236;
      107403:data<=16'd3374;
      107404:data<=16'd7436;
      107405:data<=16'd11544;
      107406:data<=16'd11194;
      107407:data<=16'd10702;
      107408:data<=16'd10981;
      107409:data<=16'd10020;
      107410:data<=16'd10572;
      107411:data<=16'd11353;
      107412:data<=16'd10604;
      107413:data<=16'd10777;
      107414:data<=16'd11079;
      107415:data<=16'd10549;
      107416:data<=16'd9785;
      107417:data<=16'd9213;
      107418:data<=16'd9721;
      107419:data<=16'd9511;
      107420:data<=16'd8696;
      107421:data<=16'd8950;
      107422:data<=16'd8467;
      107423:data<=16'd8742;
      107424:data<=16'd10619;
      107425:data<=16'd10749;
      107426:data<=16'd10213;
      107427:data<=16'd9603;
      107428:data<=16'd8072;
      107429:data<=16'd8219;
      107430:data<=16'd8906;
      107431:data<=16'd7924;
      107432:data<=16'd7288;
      107433:data<=16'd7450;
      107434:data<=16'd7224;
      107435:data<=16'd6752;
      107436:data<=16'd6749;
      107437:data<=16'd7285;
      107438:data<=16'd8771;
      107439:data<=16'd11362;
      107440:data<=16'd11905;
      107441:data<=16'd10314;
      107442:data<=16'd10320;
      107443:data<=16'd10419;
      107444:data<=16'd9633;
      107445:data<=16'd9700;
      107446:data<=16'd9447;
      107447:data<=16'd9027;
      107448:data<=16'd8296;
      107449:data<=16'd7668;
      107450:data<=16'd9477;
      107451:data<=16'd9887;
      107452:data<=16'd8328;
      107453:data<=16'd9007;
      107454:data<=16'd8163;
      107455:data<=16'd6449;
      107456:data<=16'd7671;
      107457:data<=16'd5315;
      107458:data<=-16'd616;
      107459:data<=-16'd2587;
      107460:data<=-16'd1932;
      107461:data<=-16'd1865;
      107462:data<=-16'd1929;
      107463:data<=-16'd1434;
      107464:data<=16'd80;
      107465:data<=16'd967;
      107466:data<=16'd567;
      107467:data<=16'd717;
      107468:data<=16'd836;
      107469:data<=16'd53;
      107470:data<=16'd208;
      107471:data<=16'd789;
      107472:data<=16'd0;
      107473:data<=-16'd197;
      107474:data<=-16'd47;
      107475:data<=-16'd1483;
      107476:data<=-16'd1075;
      107477:data<=16'd1210;
      107478:data<=16'd1685;
      107479:data<=16'd1721;
      107480:data<=16'd1216;
      107481:data<=16'd325;
      107482:data<=16'd1289;
      107483:data<=16'd188;
      107484:data<=-16'd2943;
      107485:data<=-16'd3143;
      107486:data<=-16'd2789;
      107487:data<=-16'd3286;
      107488:data<=-16'd2910;
      107489:data<=-16'd2376;
      107490:data<=-16'd1263;
      107491:data<=-16'd684;
      107492:data<=-16'd1398;
      107493:data<=-16'd1187;
      107494:data<=-16'd732;
      107495:data<=-16'd267;
      107496:data<=16'd955;
      107497:data<=16'd925;
      107498:data<=-16'd168;
      107499:data<=-16'd816;
      107500:data<=-16'd1240;
      107501:data<=-16'd1284;
      107502:data<=-16'd807;
      107503:data<=-16'd44;
      107504:data<=16'd591;
      107505:data<=16'd778;
      107506:data<=16'd532;
      107507:data<=16'd92;
      107508:data<=-16'd205;
      107509:data<=-16'd296;
      107510:data<=16'd2432;
      107511:data<=16'd7865;
      107512:data<=16'd9342;
      107513:data<=16'd7855;
      107514:data<=16'd7970;
      107515:data<=16'd6981;
      107516:data<=16'd7013;
      107517:data<=16'd8972;
      107518:data<=16'd7726;
      107519:data<=16'd6672;
      107520:data<=16'd7386;
      107521:data<=16'd6466;
      107522:data<=16'd6067;
      107523:data<=16'd5336;
      107524:data<=16'd3924;
      107525:data<=16'd3990;
      107526:data<=16'd3242;
      107527:data<=16'd3935;
      107528:data<=16'd6921;
      107529:data<=16'd7736;
      107530:data<=16'd8369;
      107531:data<=16'd9016;
      107532:data<=16'd7871;
      107533:data<=16'd7636;
      107534:data<=16'd7012;
      107535:data<=16'd5844;
      107536:data<=16'd6472;
      107537:data<=16'd6307;
      107538:data<=16'd5098;
      107539:data<=16'd4881;
      107540:data<=16'd4871;
      107541:data<=16'd4258;
      107542:data<=16'd3847;
      107543:data<=16'd4936;
      107544:data<=16'd5321;
      107545:data<=16'd4049;
      107546:data<=16'd3927;
      107547:data<=16'd3322;
      107548:data<=16'd2120;
      107549:data<=16'd2729;
      107550:data<=16'd2599;
      107551:data<=16'd1774;
      107552:data<=16'd1489;
      107553:data<=16'd1142;
      107554:data<=16'd2032;
      107555:data<=16'd1839;
      107556:data<=16'd651;
      107557:data<=16'd1630;
      107558:data<=16'd1908;
      107559:data<=16'd1632;
      107560:data<=16'd1651;
      107561:data<=16'd435;
      107562:data<=16'd1139;
      107563:data<=-16'd241;
      107564:data<=-16'd6617;
      107565:data<=-16'd8947;
      107566:data<=-16'd8143;
      107567:data<=-16'd8990;
      107568:data<=-16'd8100;
      107569:data<=-16'd7511;
      107570:data<=-16'd7912;
      107571:data<=-16'd6781;
      107572:data<=-16'd7865;
      107573:data<=-16'd10898;
      107574:data<=-16'd11879;
      107575:data<=-16'd11453;
      107576:data<=-16'd10809;
      107577:data<=-16'd10328;
      107578:data<=-16'd10187;
      107579:data<=-16'd10310;
      107580:data<=-16'd10505;
      107581:data<=-16'd10272;
      107582:data<=-16'd10590;
      107583:data<=-16'd11600;
      107584:data<=-16'd11920;
      107585:data<=-16'd11659;
      107586:data<=-16'd11402;
      107587:data<=-16'd11367;
      107588:data<=-16'd10847;
      107589:data<=-16'd10032;
      107590:data<=-16'd10502;
      107591:data<=-16'd10475;
      107592:data<=-16'd9336;
      107593:data<=-16'd9429;
      107594:data<=-16'd9418;
      107595:data<=-16'd9288;
      107596:data<=-16'd10452;
      107597:data<=-16'd10605;
      107598:data<=-16'd9946;
      107599:data<=-16'd9894;
      107600:data<=-16'd9547;
      107601:data<=-16'd9245;
      107602:data<=-16'd8898;
      107603:data<=-16'd8649;
      107604:data<=-16'd9004;
      107605:data<=-16'd8692;
      107606:data<=-16'd8422;
      107607:data<=-16'd8478;
      107608:data<=-16'd7803;
      107609:data<=-16'd8502;
      107610:data<=-16'd10009;
      107611:data<=-16'd9583;
      107612:data<=-16'd8898;
      107613:data<=-16'd8583;
      107614:data<=-16'd8440;
      107615:data<=-16'd9447;
      107616:data<=-16'd6743;
      107617:data<=16'd1434;
      107618:data<=16'd5937;
      107619:data<=16'd4579;
      107620:data<=16'd4170;
      107621:data<=16'd4087;
      107622:data<=16'd2158;
      107623:data<=16'd940;
      107624:data<=16'd423;
      107625:data<=16'd461;
      107626:data<=16'd1181;
      107627:data<=16'd998;
      107628:data<=16'd666;
      107629:data<=16'd70;
      107630:data<=-16'd792;
      107631:data<=16'd188;
      107632:data<=16'd616;
      107633:data<=-16'd472;
      107634:data<=-16'd234;
      107635:data<=-16'd277;
      107636:data<=-16'd1453;
      107637:data<=-16'd2241;
      107638:data<=-16'd2779;
      107639:data<=-16'd2458;
      107640:data<=-16'd2276;
      107641:data<=-16'd2946;
      107642:data<=-16'd3057;
      107643:data<=-16'd3432;
      107644:data<=-16'd3488;
      107645:data<=-16'd2358;
      107646:data<=-16'd2167;
      107647:data<=-16'd2814;
      107648:data<=-16'd3627;
      107649:data<=-16'd4623;
      107650:data<=-16'd4987;
      107651:data<=-16'd5190;
      107652:data<=-16'd5028;
      107653:data<=-16'd4566;
      107654:data<=-16'd4686;
      107655:data<=-16'd4716;
      107656:data<=-16'd4927;
      107657:data<=-16'd4843;
      107658:data<=-16'd4238;
      107659:data<=-16'd4299;
      107660:data<=-16'd3513;
      107661:data<=-16'd4143;
      107662:data<=-16'd8257;
      107663:data<=-16'd10003;
      107664:data<=-16'd9081;
      107665:data<=-16'd8884;
      107666:data<=-16'd8464;
      107667:data<=-16'd8504;
      107668:data<=-16'd8056;
      107669:data<=-16'd8661;
      107670:data<=-16'd13559;
      107671:data<=-16'd16489;
      107672:data<=-16'd15849;
      107673:data<=-16'd15861;
      107674:data<=-16'd14366;
      107675:data<=-16'd13658;
      107676:data<=-16'd15620;
      107677:data<=-16'd15620;
      107678:data<=-16'd14580;
      107679:data<=-16'd14061;
      107680:data<=-16'd13494;
      107681:data<=-16'd13438;
      107682:data<=-16'd12266;
      107683:data<=-16'd11059;
      107684:data<=-16'd11035;
      107685:data<=-16'd10348;
      107686:data<=-16'd9699;
      107687:data<=-16'd9144;
      107688:data<=-16'd9051;
      107689:data<=-16'd10452;
      107690:data<=-16'd11083;
      107691:data<=-16'd10922;
      107692:data<=-16'd10199;
      107693:data<=-16'd8378;
      107694:data<=-16'd7928;
      107695:data<=-16'd7867;
      107696:data<=-16'd7141;
      107697:data<=-16'd7362;
      107698:data<=-16'd6983;
      107699:data<=-16'd6247;
      107700:data<=-16'd6021;
      107701:data<=-16'd5777;
      107702:data<=-16'd6795;
      107703:data<=-16'd7279;
      107704:data<=-16'd6852;
      107705:data<=-16'd6937;
      107706:data<=-16'd4555;
      107707:data<=-16'd1551;
      107708:data<=-16'd1108;
      107709:data<=-16'd940;
      107710:data<=-16'd1136;
      107711:data<=-16'd1045;
      107712:data<=-16'd130;
      107713:data<=-16'd456;
      107714:data<=-16'd384;
      107715:data<=-16'd729;
      107716:data<=-16'd2443;
      107717:data<=-16'd1868;
      107718:data<=-16'd1169;
      107719:data<=-16'd1851;
      107720:data<=-16'd978;
      107721:data<=-16'd726;
      107722:data<=-16'd444;
      107723:data<=16'd3664;
      107724:data<=16'd7914;
      107725:data<=16'd8301;
      107726:data<=16'd7444;
      107727:data<=16'd7787;
      107728:data<=16'd7250;
      107729:data<=16'd5456;
      107730:data<=16'd4830;
      107731:data<=16'd4581;
      107732:data<=16'd4414;
      107733:data<=16'd4836;
      107734:data<=16'd4299;
      107735:data<=16'd4293;
      107736:data<=16'd5013;
      107737:data<=16'd4513;
      107738:data<=16'd4531;
      107739:data<=16'd4672;
      107740:data<=16'd4350;
      107741:data<=16'd4579;
      107742:data<=16'd3253;
      107743:data<=16'd2237;
      107744:data<=16'd3166;
      107745:data<=16'd2692;
      107746:data<=16'd2353;
      107747:data<=16'd2971;
      107748:data<=16'd2726;
      107749:data<=16'd3148;
      107750:data<=16'd2406;
      107751:data<=-16'd132;
      107752:data<=-16'd1084;
      107753:data<=-16'd1215;
      107754:data<=-16'd999;
      107755:data<=-16'd775;
      107756:data<=-16'd2003;
      107757:data<=-16'd1973;
      107758:data<=-16'd967;
      107759:data<=-16'd1955;
      107760:data<=-16'd2667;
      107761:data<=-16'd1886;
      107762:data<=-16'd1468;
      107763:data<=-16'd1468;
      107764:data<=-16'd1289;
      107765:data<=-16'd1151;
      107766:data<=-16'd1011;
      107767:data<=-16'd361;
      107768:data<=-16'd252;
      107769:data<=-16'd1312;
      107770:data<=-16'd1459;
      107771:data<=-16'd537;
      107772:data<=-16'd177;
      107773:data<=-16'd429;
      107774:data<=-16'd271;
      107775:data<=16'd370;
      107776:data<=-16'd2228;
      107777:data<=-16'd7577;
      107778:data<=-16'd8619;
      107779:data<=-16'd6854;
      107780:data<=-16'd7021;
      107781:data<=-16'd6655;
      107782:data<=-16'd6216;
      107783:data<=-16'd6488;
      107784:data<=-16'd5075;
      107785:data<=-16'd4164;
      107786:data<=-16'd4652;
      107787:data<=-16'd4508;
      107788:data<=-16'd4067;
      107789:data<=-16'd3133;
      107790:data<=-16'd2526;
      107791:data<=-16'd2928;
      107792:data<=-16'd2482;
      107793:data<=-16'd2238;
      107794:data<=-16'd2309;
      107795:data<=16'd444;
      107796:data<=16'd4143;
      107797:data<=16'd5168;
      107798:data<=16'd5063;
      107799:data<=16'd5510;
      107800:data<=16'd5397;
      107801:data<=16'd4817;
      107802:data<=16'd4905;
      107803:data<=16'd5231;
      107804:data<=16'd5421;
      107805:data<=16'd5547;
      107806:data<=16'd5325;
      107807:data<=16'd5382;
      107808:data<=16'd6191;
      107809:data<=16'd7536;
      107810:data<=16'd8437;
      107811:data<=16'd7432;
      107812:data<=16'd6619;
      107813:data<=16'd7636;
      107814:data<=16'd7215;
      107815:data<=16'd5586;
      107816:data<=16'd5689;
      107817:data<=16'd6246;
      107818:data<=16'd6269;
      107819:data<=16'd6062;
      107820:data<=16'd5662;
      107821:data<=16'd6305;
      107822:data<=16'd7597;
      107823:data<=16'd8285;
      107824:data<=16'd8011;
      107825:data<=16'd6666;
      107826:data<=16'd6352;
      107827:data<=16'd6857;
      107828:data<=16'd6143;
      107829:data<=16'd8355;
      107830:data<=16'd13905;
      107831:data<=16'd15526;
      107832:data<=16'd14187;
      107833:data<=16'd14289;
      107834:data<=16'd13864;
      107835:data<=16'd13891;
      107836:data<=16'd15076;
      107837:data<=16'd14254;
      107838:data<=16'd13547;
      107839:data<=16'd13095;
      107840:data<=16'd9808;
      107841:data<=16'd7953;
      107842:data<=16'd8502;
      107843:data<=16'd7464;
      107844:data<=16'd7172;
      107845:data<=16'd7777;
      107846:data<=16'd7151;
      107847:data<=16'd7835;
      107848:data<=16'd8951;
      107849:data<=16'd8689;
      107850:data<=16'd8516;
      107851:data<=16'd7891;
      107852:data<=16'd7280;
      107853:data<=16'd7313;
      107854:data<=16'd6586;
      107855:data<=16'd6102;
      107856:data<=16'd6237;
      107857:data<=16'd5896;
      107858:data<=16'd5595;
      107859:data<=16'd5442;
      107860:data<=16'd5887;
      107861:data<=16'd7106;
      107862:data<=16'd7750;
      107863:data<=16'd7545;
      107864:data<=16'd6936;
      107865:data<=16'd6683;
      107866:data<=16'd6766;
      107867:data<=16'd6153;
      107868:data<=16'd5812;
      107869:data<=16'd5796;
      107870:data<=16'd5238;
      107871:data<=16'd5385;
      107872:data<=16'd5418;
      107873:data<=16'd4681;
      107874:data<=16'd5532;
      107875:data<=16'd7353;
      107876:data<=16'd7501;
      107877:data<=16'd6498;
      107878:data<=16'd6499;
      107879:data<=16'd6560;
      107880:data<=16'd5624;
      107881:data<=16'd5923;
      107882:data<=16'd3783;
      107883:data<=-16'd2975;
      107884:data<=-16'd3935;
      107885:data<=16'd617;
      107886:data<=16'd423;
      107887:data<=16'd36;
      107888:data<=16'd2839;
      107889:data<=16'd3480;
      107890:data<=16'd3441;
      107891:data<=16'd3573;
      107892:data<=16'd2798;
      107893:data<=16'd3007;
      107894:data<=16'd3080;
      107895:data<=16'd2767;
      107896:data<=16'd2793;
      107897:data<=16'd2179;
      107898:data<=16'd2100;
      107899:data<=16'd2000;
      107900:data<=16'd1438;
      107901:data<=16'd2394;
      107902:data<=16'd3415;
      107903:data<=16'd3774;
      107904:data<=16'd4191;
      107905:data<=16'd3641;
      107906:data<=16'd3280;
      107907:data<=16'd3334;
      107908:data<=16'd2943;
      107909:data<=16'd3271;
      107910:data<=16'd3146;
      107911:data<=16'd2185;
      107912:data<=16'd2196;
      107913:data<=16'd2334;
      107914:data<=16'd2613;
      107915:data<=16'd3779;
      107916:data<=16'd4209;
      107917:data<=16'd3568;
      107918:data<=16'd3206;
      107919:data<=16'd3289;
      107920:data<=16'd2949;
      107921:data<=16'd2450;
      107922:data<=16'd2420;
      107923:data<=16'd2146;
      107924:data<=16'd2059;
      107925:data<=16'd2064;
      107926:data<=16'd1204;
      107927:data<=16'd1627;
      107928:data<=16'd2617;
      107929:data<=16'd1001;
      107930:data<=-16'd1063;
      107931:data<=-16'd1626;
      107932:data<=-16'd1257;
      107933:data<=-16'd908;
      107934:data<=-16'd1839;
      107935:data<=-16'd240;
      107936:data<=16'd5071;
      107937:data<=16'd7547;
      107938:data<=16'd6737;
      107939:data<=16'd6035;
      107940:data<=16'd5527;
      107941:data<=16'd6451;
      107942:data<=16'd7509;
      107943:data<=16'd6698;
      107944:data<=16'd6082;
      107945:data<=16'd5764;
      107946:data<=16'd5081;
      107947:data<=16'd4895;
      107948:data<=16'd4737;
      107949:data<=16'd4393;
      107950:data<=16'd3943;
      107951:data<=16'd3629;
      107952:data<=16'd3462;
      107953:data<=16'd2964;
      107954:data<=16'd3712;
      107955:data<=16'd5054;
      107956:data<=16'd4702;
      107957:data<=16'd4570;
      107958:data<=16'd4599;
      107959:data<=16'd3277;
      107960:data<=16'd2699;
      107961:data<=16'd2870;
      107962:data<=16'd2584;
      107963:data<=16'd2094;
      107964:data<=16'd1485;
      107965:data<=16'd1480;
      107966:data<=16'd1351;
      107967:data<=16'd1577;
      107968:data<=16'd3284;
      107969:data<=16'd3218;
      107970:data<=16'd2303;
      107971:data<=16'd3122;
      107972:data<=16'd2482;
      107973:data<=16'd2500;
      107974:data<=16'd5318;
      107975:data<=16'd5964;
      107976:data<=16'd5040;
      107977:data<=16'd4855;
      107978:data<=16'd3970;
      107979:data<=16'd3366;
      107980:data<=16'd3615;
      107981:data<=16'd4676;
      107982:data<=16'd5476;
      107983:data<=16'd4284;
      107984:data<=16'd4014;
      107985:data<=16'd4541;
      107986:data<=16'd3701;
      107987:data<=16'd3950;
      107988:data<=16'd2161;
      107989:data<=-16'd3715;
      107990:data<=-16'd6918;
      107991:data<=-16'd6802;
      107992:data<=-16'd6731;
      107993:data<=-16'd6467;
      107994:data<=-16'd6467;
      107995:data<=-16'd6144;
      107996:data<=-16'd5712;
      107997:data<=-16'd6250;
      107998:data<=-16'd6158;
      107999:data<=-16'd5923;
      108000:data<=-16'd6290;
      108001:data<=-16'd6219;
      108002:data<=-16'd6396;
      108003:data<=-16'd6523;
      108004:data<=-16'd6308;
      108005:data<=-16'd6203;
      108006:data<=-16'd5792;
      108007:data<=-16'd6664;
      108008:data<=-16'd8360;
      108009:data<=-16'd8369;
      108010:data<=-16'd7834;
      108011:data<=-16'd7471;
      108012:data<=-16'd7345;
      108013:data<=-16'd7811;
      108014:data<=-16'd7470;
      108015:data<=-16'd7224;
      108016:data<=-16'd7412;
      108017:data<=-16'd7036;
      108018:data<=-16'd8408;
      108019:data<=-16'd10666;
      108020:data<=-16'd11536;
      108021:data<=-16'd12662;
      108022:data<=-16'd13042;
      108023:data<=-16'd12085;
      108024:data<=-16'd11949;
      108025:data<=-16'd11771;
      108026:data<=-16'd11332;
      108027:data<=-16'd11344;
      108028:data<=-16'd10927;
      108029:data<=-16'd10502;
      108030:data<=-16'd10147;
      108031:data<=-16'd9812;
      108032:data<=-16'd10058;
      108033:data<=-16'd10081;
      108034:data<=-16'd10546;
      108035:data<=-16'd11524;
      108036:data<=-16'd11015;
      108037:data<=-16'd10346;
      108038:data<=-16'd10298;
      108039:data<=-16'd9389;
      108040:data<=-16'd9395;
      108041:data<=-16'd9236;
      108042:data<=-16'd4761;
      108043:data<=16'd159;
      108044:data<=16'd517;
      108045:data<=-16'd329;
      108046:data<=-16'd271;
      108047:data<=-16'd1142;
      108048:data<=-16'd2017;
      108049:data<=-16'd2385;
      108050:data<=-16'd2993;
      108051:data<=-16'd2874;
      108052:data<=-16'd2247;
      108053:data<=-16'd2049;
      108054:data<=-16'd2362;
      108055:data<=-16'd3058;
      108056:data<=-16'd2939;
      108057:data<=-16'd2435;
      108058:data<=-16'd2613;
      108059:data<=-16'd2411;
      108060:data<=-16'd3011;
      108061:data<=-16'd4696;
      108062:data<=-16'd3861;
      108063:data<=-16'd1319;
      108064:data<=-16'd494;
      108065:data<=-16'd478;
      108066:data<=16'd55;
      108067:data<=16'd24;
      108068:data<=-16'd781;
      108069:data<=-16'd813;
      108070:data<=-16'd312;
      108071:data<=-16'd426;
      108072:data<=-16'd121;
      108073:data<=-16'd546;
      108074:data<=-16'd2911;
      108075:data<=-16'd3833;
      108076:data<=-16'd3112;
      108077:data<=-16'd3101;
      108078:data<=-16'd2828;
      108079:data<=-16'd2585;
      108080:data<=-16'd2728;
      108081:data<=-16'd2103;
      108082:data<=-16'd1838;
      108083:data<=-16'd2522;
      108084:data<=-16'd2946;
      108085:data<=-16'd2538;
      108086:data<=-16'd2340;
      108087:data<=-16'd3635;
      108088:data<=-16'd4698;
      108089:data<=-16'd4676;
      108090:data<=-16'd4575;
      108091:data<=-16'd3685;
      108092:data<=-16'd3644;
      108093:data<=-16'd4325;
      108094:data<=-16'd3348;
      108095:data<=-16'd5774;
      108096:data<=-16'd11684;
      108097:data<=-16'd12819;
      108098:data<=-16'd11233;
      108099:data<=-16'd11442;
      108100:data<=-16'd11509;
      108101:data<=-16'd12333;
      108102:data<=-16'd13204;
      108103:data<=-16'd11963;
      108104:data<=-16'd11294;
      108105:data<=-16'd10874;
      108106:data<=-16'd9360;
      108107:data<=-16'd10520;
      108108:data<=-16'd13790;
      108109:data<=-16'd14175;
      108110:data<=-16'd12530;
      108111:data<=-16'd11887;
      108112:data<=-16'd11496;
      108113:data<=-16'd11477;
      108114:data<=-16'd12628;
      108115:data<=-16'd12989;
      108116:data<=-16'd12240;
      108117:data<=-16'd11911;
      108118:data<=-16'd11415;
      108119:data<=-16'd10357;
      108120:data<=-16'd9577;
      108121:data<=-16'd9230;
      108122:data<=-16'd8742;
      108123:data<=-16'd7929;
      108124:data<=-16'd7486;
      108125:data<=-16'd7269;
      108126:data<=-16'd7345;
      108127:data<=-16'd8633;
      108128:data<=-16'd9354;
      108129:data<=-16'd8402;
      108130:data<=-16'd7658;
      108131:data<=-16'd7285;
      108132:data<=-16'd7094;
      108133:data<=-16'd6963;
      108134:data<=-16'd5941;
      108135:data<=-16'd5353;
      108136:data<=-16'd5297;
      108137:data<=-16'd4446;
      108138:data<=-16'd3968;
      108139:data<=-16'd3845;
      108140:data<=-16'd4352;
      108141:data<=-16'd6108;
      108142:data<=-16'd5873;
      108143:data<=-16'd4379;
      108144:data<=-16'd4840;
      108145:data<=-16'd4120;
      108146:data<=-16'd2823;
      108147:data<=-16'd4112;
      108148:data<=-16'd1610;
      108149:data<=16'd5379;
      108150:data<=16'd6946;
      108151:data<=16'd5509;
      108152:data<=16'd8675;
      108153:data<=16'd10534;
      108154:data<=16'd7987;
      108155:data<=16'd6909;
      108156:data<=16'd6960;
      108157:data<=16'd6373;
      108158:data<=16'd6862;
      108159:data<=16'd7172;
      108160:data<=16'd6485;
      108161:data<=16'd6122;
      108162:data<=16'd6370;
      108163:data<=16'd6669;
      108164:data<=16'd6275;
      108165:data<=16'd5958;
      108166:data<=16'd5313;
      108167:data<=16'd3363;
      108168:data<=16'd3049;
      108169:data<=16'd4081;
      108170:data<=16'd3466;
      108171:data<=16'd3363;
      108172:data<=16'd4052;
      108173:data<=16'd3659;
      108174:data<=16'd3735;
      108175:data<=16'd4137;
      108176:data<=16'd4020;
      108177:data<=16'd4244;
      108178:data<=16'd4379;
      108179:data<=16'd3633;
      108180:data<=16'd1994;
      108181:data<=16'd1010;
      108182:data<=16'd1598;
      108183:data<=16'd1862;
      108184:data<=16'd1415;
      108185:data<=16'd1192;
      108186:data<=16'd1325;
      108187:data<=16'd1885;
      108188:data<=16'd1991;
      108189:data<=16'd1697;
      108190:data<=16'd1400;
      108191:data<=16'd1257;
      108192:data<=16'd1871;
      108193:data<=16'd917;
      108194:data<=-16'd713;
      108195:data<=16'd129;
      108196:data<=-16'd790;
      108197:data<=-16'd3638;
      108198:data<=-16'd4137;
      108199:data<=-16'd4021;
      108200:data<=-16'd3195;
      108201:data<=-16'd4143;
      108202:data<=-16'd9682;
      108203:data<=-16'd11806;
      108204:data<=-16'd9993;
      108205:data<=-16'd9959;
      108206:data<=-16'd8909;
      108207:data<=-16'd8023;
      108208:data<=-16'd8646;
      108209:data<=-16'd7617;
      108210:data<=-16'd6972;
      108211:data<=-16'd6695;
      108212:data<=-16'd6078;
      108213:data<=-16'd6548;
      108214:data<=-16'd5624;
      108215:data<=-16'd4417;
      108216:data<=-16'd4322;
      108217:data<=-16'd3568;
      108218:data<=-16'd4050;
      108219:data<=-16'd3879;
      108220:data<=-16'd1483;
      108221:data<=-16'd989;
      108222:data<=-16'd1131;
      108223:data<=-16'd362;
      108224:data<=-16'd297;
      108225:data<=-16'd150;
      108226:data<=-16'd33;
      108227:data<=16'd449;
      108228:data<=16'd960;
      108229:data<=16'd587;
      108230:data<=16'd1303;
      108231:data<=16'd1415;
      108232:data<=16'd886;
      108233:data<=16'd2995;
      108234:data<=16'd4291;
      108235:data<=16'd4050;
      108236:data<=16'd4728;
      108237:data<=16'd4323;
      108238:data<=16'd4109;
      108239:data<=16'd4375;
      108240:data<=16'd4074;
      108241:data<=16'd6335;
      108242:data<=16'd8824;
      108243:data<=16'd8812;
      108244:data<=16'd8943;
      108245:data<=16'd9037;
      108246:data<=16'd9309;
      108247:data<=16'd10216;
      108248:data<=16'd10372;
      108249:data<=16'd10241;
      108250:data<=16'd9464;
      108251:data<=16'd8912;
      108252:data<=16'd8892;
      108253:data<=16'd7629;
      108254:data<=16'd9656;
      108255:data<=16'd15377;
      108256:data<=16'd17027;
      108257:data<=16'd15575;
      108258:data<=16'd15264;
      108259:data<=16'd15452;
      108260:data<=16'd16260;
      108261:data<=16'd16475;
      108262:data<=16'd15540;
      108263:data<=16'd15409;
      108264:data<=16'd15314;
      108265:data<=16'd14360;
      108266:data<=16'd13614;
      108267:data<=16'd13115;
      108268:data<=16'd12314;
      108269:data<=16'd11949;
      108270:data<=16'd12190;
      108271:data<=16'd11391;
      108272:data<=16'd11050;
      108273:data<=16'd12769;
      108274:data<=16'd13195;
      108275:data<=16'd12439;
      108276:data<=16'd12345;
      108277:data<=16'd11311;
      108278:data<=16'd10898;
      108279:data<=16'd11136;
      108280:data<=16'd9802;
      108281:data<=16'd9357;
      108282:data<=16'd9439;
      108283:data<=16'd8707;
      108284:data<=16'd9060;
      108285:data<=16'd8029;
      108286:data<=16'd5474;
      108287:data<=16'd5354;
      108288:data<=16'd5827;
      108289:data<=16'd5075;
      108290:data<=16'd4579;
      108291:data<=16'd4441;
      108292:data<=16'd4676;
      108293:data<=16'd4801;
      108294:data<=16'd4466;
      108295:data<=16'd4196;
      108296:data<=16'd3826;
      108297:data<=16'd3930;
      108298:data<=16'd4170;
      108299:data<=16'd3965;
      108300:data<=16'd5016;
      108301:data<=16'd6141;
      108302:data<=16'd5474;
      108303:data<=16'd5010;
      108304:data<=16'd4514;
      108305:data<=16'd3738;
      108306:data<=16'd4798;
      108307:data<=16'd3744;
      108308:data<=-16'd2149;
      108309:data<=-16'd5771;
      108310:data<=-16'd4767;
      108311:data<=-16'd4270;
      108312:data<=-16'd3677;
      108313:data<=-16'd1639;
      108314:data<=-16'd1284;
      108315:data<=-16'd1915;
      108316:data<=-16'd1354;
      108317:data<=-16'd1101;
      108318:data<=-16'd1451;
      108319:data<=-16'd1281;
      108320:data<=-16'd1102;
      108321:data<=-16'd1140;
      108322:data<=-16'd879;
      108323:data<=-16'd817;
      108324:data<=-16'd1163;
      108325:data<=-16'd720;
      108326:data<=16'd732;
      108327:data<=16'd1939;
      108328:data<=16'd1724;
      108329:data<=16'd638;
      108330:data<=16'd1841;
      108331:data<=16'd4934;
      108332:data<=16'd5495;
      108333:data<=16'd4684;
      108334:data<=16'd4930;
      108335:data<=16'd4645;
      108336:data<=16'd4683;
      108337:data<=16'd4913;
      108338:data<=16'd3795;
      108339:data<=16'd4094;
      108340:data<=16'd5864;
      108341:data<=16'd6244;
      108342:data<=16'd5736;
      108343:data<=16'd5116;
      108344:data<=16'd4713;
      108345:data<=16'd4520;
      108346:data<=16'd4108;
      108347:data<=16'd3971;
      108348:data<=16'd3629;
      108349:data<=16'd3492;
      108350:data<=16'd3858;
      108351:data<=16'd3297;
      108352:data<=16'd3706;
      108353:data<=16'd5133;
      108354:data<=16'd4758;
      108355:data<=16'd4525;
      108356:data<=16'd4607;
      108357:data<=16'd3568;
      108358:data<=16'd3501;
      108359:data<=16'd3445;
      108360:data<=16'd3685;
      108361:data<=16'd7373;
      108362:data<=16'd11177;
      108363:data<=16'd11300;
      108364:data<=16'd10119;
      108365:data<=16'd10536;
      108366:data<=16'd11577;
      108367:data<=16'd10907;
      108368:data<=16'd9996;
      108369:data<=16'd10193;
      108370:data<=16'd9700;
      108371:data<=16'd8725;
      108372:data<=16'd8225;
      108373:data<=16'd8119;
      108374:data<=16'd7294;
      108375:data<=16'd4138;
      108376:data<=16'd1353;
      108377:data<=16'd1102;
      108378:data<=16'd1853;
      108379:data<=16'd3645;
      108380:data<=16'd4599;
      108381:data<=16'd3563;
      108382:data<=16'd3488;
      108383:data<=16'd3727;
      108384:data<=16'd3242;
      108385:data<=16'd2943;
      108386:data<=16'd1996;
      108387:data<=16'd1386;
      108388:data<=16'd1506;
      108389:data<=16'd1190;
      108390:data<=16'd1011;
      108391:data<=16'd848;
      108392:data<=16'd1560;
      108393:data<=16'd2987;
      108394:data<=16'd2669;
      108395:data<=16'd2106;
      108396:data<=16'd2202;
      108397:data<=16'd1760;
      108398:data<=16'd1780;
      108399:data<=16'd1280;
      108400:data<=16'd123;
      108401:data<=16'd202;
      108402:data<=16'd502;
      108403:data<=16'd400;
      108404:data<=16'd59;
      108405:data<=-16'd12;
      108406:data<=16'd1296;
      108407:data<=16'd2080;
      108408:data<=16'd1601;
      108409:data<=16'd1416;
      108410:data<=16'd1111;
      108411:data<=16'd575;
      108412:data<=16'd719;
      108413:data<=16'd1207;
      108414:data<=-16'd1879;
      108415:data<=-16'd8478;
      108416:data<=-16'd9867;
      108417:data<=-16'd7561;
      108418:data<=-16'd8810;
      108419:data<=-16'd7714;
      108420:data<=-16'd3750;
      108421:data<=-16'd3372;
      108422:data<=-16'd3535;
      108423:data<=-16'd3427;
      108424:data<=-16'd4373;
      108425:data<=-16'd4270;
      108426:data<=-16'd4181;
      108427:data<=-16'd3730;
      108428:data<=-16'd3551;
      108429:data<=-16'd5098;
      108430:data<=-16'd4892;
      108431:data<=-16'd4300;
      108432:data<=-16'd5448;
      108433:data<=-16'd5726;
      108434:data<=-16'd6216;
      108435:data<=-16'd6614;
      108436:data<=-16'd5938;
      108437:data<=-16'd6055;
      108438:data<=-16'd5705;
      108439:data<=-16'd5391;
      108440:data<=-16'd5849;
      108441:data<=-16'd5360;
      108442:data<=-16'd5770;
      108443:data<=-16'd6464;
      108444:data<=-16'd6058;
      108445:data<=-16'd6768;
      108446:data<=-16'd7342;
      108447:data<=-16'd7426;
      108448:data<=-16'd8129;
      108449:data<=-16'd7944;
      108450:data<=-16'd7541;
      108451:data<=-16'd7160;
      108452:data<=-16'd6811;
      108453:data<=-16'd7216;
      108454:data<=-16'd6455;
      108455:data<=-16'd5865;
      108456:data<=-16'd6525;
      108457:data<=-16'd6065;
      108458:data<=-16'd6234;
      108459:data<=-16'd7450;
      108460:data<=-16'd7924;
      108461:data<=-16'd8119;
      108462:data<=-16'd7644;
      108463:data<=-16'd8064;
      108464:data<=-16'd9473;
      108465:data<=-16'd10207;
      108466:data<=-16'd11405;
      108467:data<=-16'd8740;
      108468:data<=-16'd2199;
      108469:data<=-16'd705;
      108470:data<=-16'd1953;
      108471:data<=-16'd1815;
      108472:data<=-16'd3213;
      108473:data<=-16'd3594;
      108474:data<=-16'd2858;
      108475:data<=-16'd3386;
      108476:data<=-16'd2834;
      108477:data<=-16'd2444;
      108478:data<=-16'd2975;
      108479:data<=-16'd2692;
      108480:data<=-16'd2702;
      108481:data<=-16'd2634;
      108482:data<=-16'd2663;
      108483:data<=-16'd3200;
      108484:data<=-16'd2817;
      108485:data<=-16'd3427;
      108486:data<=-16'd4960;
      108487:data<=-16'd4837;
      108488:data<=-16'd4411;
      108489:data<=-16'd4126;
      108490:data<=-16'd3635;
      108491:data<=-16'd3806;
      108492:data<=-16'd3803;
      108493:data<=-16'd3665;
      108494:data<=-16'd3695;
      108495:data<=-16'd3448;
      108496:data<=-16'd3338;
      108497:data<=-16'd2933;
      108498:data<=-16'd3165;
      108499:data<=-16'd4790;
      108500:data<=-16'd4784;
      108501:data<=-16'd2971;
      108502:data<=-16'd2525;
      108503:data<=-16'd3083;
      108504:data<=-16'd2685;
      108505:data<=-16'd2000;
      108506:data<=-16'd2475;
      108507:data<=-16'd2951;
      108508:data<=-16'd1911;
      108509:data<=-16'd361;
      108510:data<=16'd488;
      108511:data<=-16'd358;
      108512:data<=-16'd2237;
      108513:data<=-16'd2353;
      108514:data<=-16'd1836;
      108515:data<=-16'd2422;
      108516:data<=-16'd2171;
      108517:data<=-16'd2130;
      108518:data<=-16'd2588;
      108519:data<=-16'd1303;
      108520:data<=-16'd3027;
      108521:data<=-16'd9215;
      108522:data<=-16'd11139;
      108523:data<=-16'd8845;
      108524:data<=-16'd9539;
      108525:data<=-16'd11456;
      108526:data<=-16'd11591;
      108527:data<=-16'd11253;
      108528:data<=-16'd10440;
      108529:data<=-16'd10058;
      108530:data<=-16'd10334;
      108531:data<=-16'd9512;
      108532:data<=-16'd8818;
      108533:data<=-16'd8881;
      108534:data<=-16'd8275;
      108535:data<=-16'd7586;
      108536:data<=-16'd6998;
      108537:data<=-16'd6734;
      108538:data<=-16'd7837;
      108539:data<=-16'd8863;
      108540:data<=-16'd8655;
      108541:data<=-16'd8094;
      108542:data<=-16'd7699;
      108543:data<=-16'd7341;
      108544:data<=-16'd6639;
      108545:data<=-16'd6313;
      108546:data<=-16'd6429;
      108547:data<=-16'd5485;
      108548:data<=-16'd4552;
      108549:data<=-16'd4866;
      108550:data<=-16'd5325;
      108551:data<=-16'd5880;
      108552:data<=-16'd6440;
      108553:data<=-16'd6913;
      108554:data<=-16'd7881;
      108555:data<=-16'd8056;
      108556:data<=-16'd7081;
      108557:data<=-16'd6687;
      108558:data<=-16'd6851;
      108559:data<=-16'd6413;
      108560:data<=-16'd5517;
      108561:data<=-16'd4971;
      108562:data<=-16'd4499;
      108563:data<=-16'd4193;
      108564:data<=-16'd4986;
      108565:data<=-16'd5927;
      108566:data<=-16'd6225;
      108567:data<=-16'd6131;
      108568:data<=-16'd5611;
      108569:data<=-16'd5482;
      108570:data<=-16'd4616;
      108571:data<=-16'd3427;
      108572:data<=-16'd4686;
      108573:data<=-16'd3186;
      108574:data<=16'd2995;
      108575:data<=16'd5442;
      108576:data<=16'd4643;
      108577:data<=16'd4639;
      108578:data<=16'd2996;
      108579:data<=16'd1848;
      108580:data<=16'd2666;
      108581:data<=16'd2710;
      108582:data<=16'd2684;
      108583:data<=16'd2760;
      108584:data<=16'd2722;
      108585:data<=16'd2987;
      108586:data<=16'd2557;
      108587:data<=16'd2400;
      108588:data<=16'd2491;
      108589:data<=16'd2290;
      108590:data<=16'd3063;
      108591:data<=16'd2532;
      108592:data<=16'd326;
      108593:data<=16'd64;
      108594:data<=16'd1017;
      108595:data<=16'd1251;
      108596:data<=16'd1052;
      108597:data<=16'd1157;
      108598:data<=16'd2244;
      108599:data<=16'd3260;
      108600:data<=16'd3551;
      108601:data<=16'd3403;
      108602:data<=16'd3107;
      108603:data<=16'd3589;
      108604:data<=16'd3175;
      108605:data<=16'd1165;
      108606:data<=16'd306;
      108607:data<=16'd519;
      108608:data<=16'd916;
      108609:data<=16'd1374;
      108610:data<=16'd1146;
      108611:data<=16'd1234;
      108612:data<=16'd1222;
      108613:data<=16'd925;
      108614:data<=16'd1653;
      108615:data<=16'd1524;
      108616:data<=16'd908;
      108617:data<=16'd954;
      108618:data<=-16'd291;
      108619:data<=-16'd776;
      108620:data<=-16'd65;
      108621:data<=-16'd314;
      108622:data<=16'd563;
      108623:data<=16'd907;
      108624:data<=-16'd144;
      108625:data<=16'd1095;
      108626:data<=16'd334;
      108627:data<=-16'd4837;
      108628:data<=-16'd7749;
      108629:data<=-16'd7462;
      108630:data<=-16'd7092;
      108631:data<=-16'd6314;
      108632:data<=-16'd5242;
      108633:data<=-16'd5125;
      108634:data<=-16'd5647;
      108635:data<=-16'd5294;
      108636:data<=-16'd4696;
      108637:data<=-16'd4643;
      108638:data<=-16'd3877;
      108639:data<=-16'd3513;
      108640:data<=-16'd3785;
      108641:data<=-16'd2917;
      108642:data<=-16'd3107;
      108643:data<=-16'd4443;
      108644:data<=-16'd3604;
      108645:data<=-16'd1827;
      108646:data<=-16'd1334;
      108647:data<=-16'd1381;
      108648:data<=-16'd831;
      108649:data<=-16'd155;
      108650:data<=-16'd543;
      108651:data<=-16'd528;
      108652:data<=16'd303;
      108653:data<=-16'd76;
      108654:data<=-16'd344;
      108655:data<=16'd226;
      108656:data<=16'd165;
      108657:data<=16'd789;
      108658:data<=16'd2305;
      108659:data<=16'd2921;
      108660:data<=16'd2854;
      108661:data<=16'd3148;
      108662:data<=16'd3747;
      108663:data<=16'd3507;
      108664:data<=16'd2934;
      108665:data<=16'd3254;
      108666:data<=16'd3221;
      108667:data<=16'd3001;
      108668:data<=16'd3336;
      108669:data<=16'd2992;
      108670:data<=16'd3268;
      108671:data<=16'd4813;
      108672:data<=16'd5413;
      108673:data<=16'd5385;
      108674:data<=16'd5454;
      108675:data<=16'd5172;
      108676:data<=16'd5153;
      108677:data<=16'd5128;
      108678:data<=16'd4331;
      108679:data<=16'd4605;
      108680:data<=16'd8664;
      108681:data<=16'd13262;
      108682:data<=16'd12871;
      108683:data<=16'd11312;
      108684:data<=16'd12880;
      108685:data<=16'd13576;
      108686:data<=16'd13289;
      108687:data<=16'd14518;
      108688:data<=16'd14947;
      108689:data<=16'd14167;
      108690:data<=16'd13482;
      108691:data<=16'd13129;
      108692:data<=16'd13117;
      108693:data<=16'd12240;
      108694:data<=16'd11558;
      108695:data<=16'd11737;
      108696:data<=16'd10739;
      108697:data<=16'd10527;
      108698:data<=16'd11964;
      108699:data<=16'd11885;
      108700:data<=16'd11197;
      108701:data<=16'd10995;
      108702:data<=16'd10126;
      108703:data<=16'd9688;
      108704:data<=16'd9667;
      108705:data<=16'd9088;
      108706:data<=16'd8639;
      108707:data<=16'd8331;
      108708:data<=16'd7911;
      108709:data<=16'd7776;
      108710:data<=16'd8454;
      108711:data<=16'd9462;
      108712:data<=16'd9216;
      108713:data<=16'd8490;
      108714:data<=16'd8511;
      108715:data<=16'd7947;
      108716:data<=16'd7042;
      108717:data<=16'd6933;
      108718:data<=16'd6736;
      108719:data<=16'd6367;
      108720:data<=16'd6258;
      108721:data<=16'd5747;
      108722:data<=16'd5248;
      108723:data<=16'd5902;
      108724:data<=16'd6777;
      108725:data<=16'd6787;
      108726:data<=16'd7063;
      108727:data<=16'd7198;
      108728:data<=16'd6316;
      108729:data<=16'd6222;
      108730:data<=16'd5888;
      108731:data<=16'd4287;
      108732:data<=16'd3662;
      108733:data<=16'd737;
      108734:data<=-16'd5265;
      108735:data<=-16'd6993;
      108736:data<=-16'd5554;
      108737:data<=-16'd5184;
      108738:data<=-16'd3359;
      108739:data<=-16'd2106;
      108740:data<=-16'd3066;
      108741:data<=-16'd2646;
      108742:data<=-16'd2223;
      108743:data<=-16'd2872;
      108744:data<=-16'd2716;
      108745:data<=-16'd2781;
      108746:data<=-16'd2689;
      108747:data<=-16'd1839;
      108748:data<=-16'd1759;
      108749:data<=-16'd1953;
      108750:data<=-16'd1504;
      108751:data<=-16'd402;
      108752:data<=16'd446;
      108753:data<=16'd120;
      108754:data<=16'd174;
      108755:data<=16'd344;
      108756:data<=-16'd393;
      108757:data<=-16'd42;
      108758:data<=16'd587;
      108759:data<=16'd59;
      108760:data<=-16'd27;
      108761:data<=-16'd109;
      108762:data<=-16'd399;
      108763:data<=16'd334;
      108764:data<=16'd1319;
      108765:data<=16'd1823;
      108766:data<=16'd1718;
      108767:data<=16'd1541;
      108768:data<=16'd1804;
      108769:data<=16'd1394;
      108770:data<=16'd958;
      108771:data<=16'd1336;
      108772:data<=16'd1292;
      108773:data<=16'd1237;
      108774:data<=16'd1310;
      108775:data<=16'd990;
      108776:data<=16'd1817;
      108777:data<=16'd3956;
      108778:data<=16'd5269;
      108779:data<=16'd4667;
      108780:data<=16'd4109;
      108781:data<=16'd4631;
      108782:data<=16'd3917;
      108783:data<=16'd3627;
      108784:data<=16'd4470;
      108785:data<=16'd2716;
      108786:data<=16'd4000;
      108787:data<=16'd10812;
      108788:data<=16'd12340;
      108789:data<=16'd9735;
      108790:data<=16'd10868;
      108791:data<=16'd11638;
      108792:data<=16'd10549;
      108793:data<=16'd10366;
      108794:data<=16'd9841;
      108795:data<=16'd9124;
      108796:data<=16'd8621;
      108797:data<=16'd8264;
      108798:data<=16'd8025;
      108799:data<=16'd6966;
      108800:data<=16'd6675;
      108801:data<=16'd6784;
      108802:data<=16'd5588;
      108803:data<=16'd5796;
      108804:data<=16'd6983;
      108805:data<=16'd6837;
      108806:data<=16'd6924;
      108807:data<=16'd6648;
      108808:data<=16'd5447;
      108809:data<=16'd5107;
      108810:data<=16'd5046;
      108811:data<=16'd4619;
      108812:data<=16'd4194;
      108813:data<=16'd3795;
      108814:data<=16'd3494;
      108815:data<=16'd3268;
      108816:data<=16'd3862;
      108817:data<=16'd4426;
      108818:data<=16'd3996;
      108819:data<=16'd4372;
      108820:data<=16'd4190;
      108821:data<=16'd1974;
      108822:data<=16'd869;
      108823:data<=16'd901;
      108824:data<=16'd537;
      108825:data<=16'd503;
      108826:data<=-16'd30;
      108827:data<=-16'd974;
      108828:data<=-16'd1092;
      108829:data<=-16'd435;
      108830:data<=16'd509;
      108831:data<=16'd526;
      108832:data<=16'd487;
      108833:data<=16'd1077;
      108834:data<=16'd631;
      108835:data<=16'd596;
      108836:data<=16'd663;
      108837:data<=-16'd462;
      108838:data<=16'd253;
      108839:data<=-16'd1222;
      108840:data<=-16'd7709;
      108841:data<=-16'd10132;
      108842:data<=-16'd8537;
      108843:data<=-16'd9050;
      108844:data<=-16'd8843;
      108845:data<=-16'd8373;
      108846:data<=-16'd9239;
      108847:data<=-16'd8684;
      108848:data<=-16'd8085;
      108849:data<=-16'd7808;
      108850:data<=-16'd7057;
      108851:data<=-16'd7486;
      108852:data<=-16'd7413;
      108853:data<=-16'd6778;
      108854:data<=-16'd7101;
      108855:data<=-16'd6611;
      108856:data<=-16'd6670;
      108857:data<=-16'd8182;
      108858:data<=-16'd8508;
      108859:data<=-16'd8329;
      108860:data<=-16'd8633;
      108861:data<=-16'd8561;
      108862:data<=-16'd8067;
      108863:data<=-16'd7718;
      108864:data<=-16'd8081;
      108865:data<=-16'd7212;
      108866:data<=-16'd5072;
      108867:data<=-16'd4830;
      108868:data<=-16'd4966;
      108869:data<=-16'd4675;
      108870:data<=-16'd6043;
      108871:data<=-16'd6630;
      108872:data<=-16'd5950;
      108873:data<=-16'd6247;
      108874:data<=-16'd6282;
      108875:data<=-16'd5974;
      108876:data<=-16'd6065;
      108877:data<=-16'd5829;
      108878:data<=-16'd5506;
      108879:data<=-16'd5372;
      108880:data<=-16'd5523;
      108881:data<=-16'd5397;
      108882:data<=-16'd5174;
      108883:data<=-16'd6229;
      108884:data<=-16'd7122;
      108885:data<=-16'd7215;
      108886:data<=-16'd7360;
      108887:data<=-16'd6675;
      108888:data<=-16'd6552;
      108889:data<=-16'd6693;
      108890:data<=-16'd5695;
      108891:data<=-16'd5949;
      108892:data<=-16'd4146;
      108893:data<=16'd1333;
      108894:data<=16'd3140;
      108895:data<=16'd2229;
      108896:data<=16'd2375;
      108897:data<=16'd954;
      108898:data<=-16'd33;
      108899:data<=16'd281;
      108900:data<=-16'd449;
      108901:data<=-16'd162;
      108902:data<=16'd393;
      108903:data<=-16'd312;
      108904:data<=-16'd147;
      108905:data<=16'd33;
      108906:data<=-16'd632;
      108907:data<=-16'd761;
      108908:data<=-16'd778;
      108909:data<=-16'd1718;
      108910:data<=-16'd3454;
      108911:data<=-16'd4535;
      108912:data<=-16'd4626;
      108913:data<=-16'd4907;
      108914:data<=-16'd4934;
      108915:data<=-16'd4579;
      108916:data<=-16'd4361;
      108917:data<=-16'd4029;
      108918:data<=-16'd4155;
      108919:data<=-16'd4358;
      108920:data<=-16'd3853;
      108921:data<=-16'd3515;
      108922:data<=-16'd3867;
      108923:data<=-16'd4968;
      108924:data<=-16'd5873;
      108925:data<=-16'd5536;
      108926:data<=-16'd5051;
      108927:data<=-16'd4874;
      108928:data<=-16'd4711;
      108929:data<=-16'd4692;
      108930:data<=-16'd4548;
      108931:data<=-16'd4657;
      108932:data<=-16'd4463;
      108933:data<=-16'd3836;
      108934:data<=-16'd4014;
      108935:data<=-16'd3756;
      108936:data<=-16'd3820;
      108937:data<=-16'd5735;
      108938:data<=-16'd5930;
      108939:data<=-16'd4532;
      108940:data<=-16'd4491;
      108941:data<=-16'd4300;
      108942:data<=-16'd4235;
      108943:data<=-16'd4363;
      108944:data<=-16'd3163;
      108945:data<=-16'd4407;
      108946:data<=-16'd9233;
      108947:data<=-16'd11966;
      108948:data<=-16'd11295;
      108949:data<=-16'd11385;
      108950:data<=-16'd12868;
      108951:data<=-16'd12628;
      108952:data<=-16'd11391;
      108953:data<=-16'd11336;
      108954:data<=-16'd10343;
      108955:data<=-16'd8372;
      108956:data<=-16'd7811;
      108957:data<=-16'd7447;
      108958:data<=-16'd6687;
      108959:data<=-16'd6557;
      108960:data<=-16'd6305;
      108961:data<=-16'd5738;
      108962:data<=-16'd5768;
      108963:data<=-16'd6448;
      108964:data<=-16'd6746;
      108965:data<=-16'd6452;
      108966:data<=-16'd6485;
      108967:data<=-16'd6267;
      108968:data<=-16'd5492;
      108969:data<=-16'd5078;
      108970:data<=-16'd4730;
      108971:data<=-16'd4511;
      108972:data<=-16'd4447;
      108973:data<=-16'd3947;
      108974:data<=-16'd3768;
      108975:data<=-16'd3902;
      108976:data<=-16'd4264;
      108977:data<=-16'd5157;
      108978:data<=-16'd4969;
      108979:data<=-16'd4185;
      108980:data<=-16'd4405;
      108981:data<=-16'd4032;
      108982:data<=-16'd2977;
      108983:data<=-16'd2877;
      108984:data<=-16'd3030;
      108985:data<=-16'd2682;
      108986:data<=-16'd2419;
      108987:data<=-16'd2217;
      108988:data<=-16'd1692;
      108989:data<=-16'd2067;
      108990:data<=-16'd3506;
      108991:data<=-16'd3598;
      108992:data<=-16'd2939;
      108993:data<=-16'd3146;
      108994:data<=-16'd2672;
      108995:data<=-16'd1856;
      108996:data<=-16'd1996;
      108997:data<=-16'd2231;
      108998:data<=-16'd1462;
      108999:data<=16'd1548;
      109000:data<=16'd4933;
      109001:data<=16'd5591;
      109002:data<=16'd4739;
      109003:data<=16'd3523;
      109004:data<=16'd2558;
      109005:data<=16'd3013;
      109006:data<=16'd3119;
      109007:data<=16'd2707;
      109008:data<=16'd3184;
      109009:data<=16'd3363;
      109010:data<=16'd3266;
      109011:data<=16'd3231;
      109012:data<=16'd2934;
      109013:data<=16'd3377;
      109014:data<=16'd3601;
      109015:data<=16'd2604;
      109016:data<=16'd1801;
      109017:data<=16'd1665;
      109018:data<=16'd1786;
      109019:data<=16'd1641;
      109020:data<=16'd1212;
      109021:data<=16'd1485;
      109022:data<=16'd2085;
      109023:data<=16'd2079;
      109024:data<=16'd1770;
      109025:data<=16'd1817;
      109026:data<=16'd2040;
      109027:data<=16'd1820;
      109028:data<=16'd1770;
      109029:data<=16'd1442;
      109030:data<=-16'd58;
      109031:data<=-16'd438;
      109032:data<=16'd271;
      109033:data<=-16'd155;
      109034:data<=-16'd156;
      109035:data<=16'd397;
      109036:data<=16'd114;
      109037:data<=16'd368;
      109038:data<=16'd789;
      109039:data<=16'd375;
      109040:data<=16'd535;
      109041:data<=16'd1189;
      109042:data<=16'd732;
      109043:data<=-16'd253;
      109044:data<=16'd623;
      109045:data<=16'd2352;
      109046:data<=16'd1996;
      109047:data<=16'd1556;
      109048:data<=16'd2417;
      109049:data<=16'd2011;
      109050:data<=16'd1882;
      109051:data<=16'd2931;
      109052:data<=16'd120;
      109053:data<=-16'd5595;
      109054:data<=-16'd7030;
      109055:data<=-16'd5225;
      109056:data<=-16'd5325;
      109057:data<=-16'd5517;
      109058:data<=-16'd4626;
      109059:data<=-16'd4778;
      109060:data<=-16'd4364;
      109061:data<=-16'd3442;
      109062:data<=-16'd3911;
      109063:data<=-16'd3771;
      109064:data<=-16'd2946;
      109065:data<=-16'd2561;
      109066:data<=-16'd1909;
      109067:data<=-16'd1964;
      109068:data<=-16'd1859;
      109069:data<=-16'd281;
      109070:data<=16'd773;
      109071:data<=16'd952;
      109072:data<=16'd1022;
      109073:data<=16'd1216;
      109074:data<=16'd1709;
      109075:data<=16'd1575;
      109076:data<=16'd1542;
      109077:data<=16'd1883;
      109078:data<=16'd1642;
      109079:data<=16'd2070;
      109080:data<=16'd2322;
      109081:data<=16'd1501;
      109082:data<=16'd2167;
      109083:data<=16'd4141;
      109084:data<=16'd5328;
      109085:data<=16'd4925;
      109086:data<=16'd4027;
      109087:data<=16'd4636;
      109088:data<=16'd4567;
      109089:data<=16'd2834;
      109090:data<=16'd2328;
      109091:data<=16'd2253;
      109092:data<=16'd1889;
      109093:data<=16'd2120;
      109094:data<=16'd2118;
      109095:data<=16'd2708;
      109096:data<=16'd3852;
      109097:data<=16'd4115;
      109098:data<=16'd3896;
      109099:data<=16'd3660;
      109100:data<=16'd3808;
      109101:data<=16'd3748;
      109102:data<=16'd3788;
      109103:data<=16'd4294;
      109104:data<=16'd3224;
      109105:data<=16'd5083;
      109106:data<=16'd11524;
      109107:data<=16'd13000;
      109108:data<=16'd11327;
      109109:data<=16'd12928;
      109110:data<=16'd12866;
      109111:data<=16'd11819;
      109112:data<=16'd12416;
      109113:data<=16'd11662;
      109114:data<=16'd11056;
      109115:data<=16'd10883;
      109116:data<=16'd10201;
      109117:data<=16'd10311;
      109118:data<=16'd9602;
      109119:data<=16'd8570;
      109120:data<=16'd8385;
      109121:data<=16'd8332;
      109122:data<=16'd9351;
      109123:data<=16'd9770;
      109124:data<=16'd8954;
      109125:data<=16'd8724;
      109126:data<=16'd8382;
      109127:data<=16'd8498;
      109128:data<=16'd8298;
      109129:data<=16'd7124;
      109130:data<=16'd7279;
      109131:data<=16'd6795;
      109132:data<=16'd6258;
      109133:data<=16'd8044;
      109134:data<=16'd8408;
      109135:data<=16'd8434;
      109136:data<=16'd9776;
      109137:data<=16'd9262;
      109138:data<=16'd8778;
      109139:data<=16'd8737;
      109140:data<=16'd7688;
      109141:data<=16'd7574;
      109142:data<=16'd7322;
      109143:data<=16'd6616;
      109144:data<=16'd6422;
      109145:data<=16'd5985;
      109146:data<=16'd5930;
      109147:data<=16'd5345;
      109148:data<=16'd5197;
      109149:data<=16'd6799;
      109150:data<=16'd6808;
      109151:data<=16'd6460;
      109152:data<=16'd6721;
      109153:data<=16'd5456;
      109154:data<=16'd5383;
      109155:data<=16'd5116;
      109156:data<=16'd3977;
      109157:data<=16'd5368;
      109158:data<=16'd3062;
      109159:data<=-16'd3648;
      109160:data<=-16'd5604;
      109161:data<=-16'd3914;
      109162:data<=-16'd2679;
      109163:data<=-16'd1876;
      109164:data<=-16'd1888;
      109165:data<=-16'd1670;
      109166:data<=-16'd1598;
      109167:data<=-16'd2032;
      109168:data<=-16'd2079;
      109169:data<=-16'd2179;
      109170:data<=-16'd1806;
      109171:data<=-16'd1917;
      109172:data<=-16'd2610;
      109173:data<=-16'd1983;
      109174:data<=-16'd1917;
      109175:data<=-16'd1337;
      109176:data<=16'd946;
      109177:data<=16'd118;
      109178:data<=-16'd2018;
      109179:data<=-16'd1554;
      109180:data<=-16'd1372;
      109181:data<=-16'd1735;
      109182:data<=-16'd1419;
      109183:data<=-16'd1369;
      109184:data<=-16'd1565;
      109185:data<=-16'd1807;
      109186:data<=-16'd1900;
      109187:data<=-16'd2314;
      109188:data<=-16'd1947;
      109189:data<=16'd582;
      109190:data<=16'd1773;
      109191:data<=16'd1054;
      109192:data<=16'd1442;
      109193:data<=16'd1759;
      109194:data<=16'd1829;
      109195:data<=16'd2191;
      109196:data<=16'd1530;
      109197:data<=16'd1031;
      109198:data<=16'd1118;
      109199:data<=16'd999;
      109200:data<=16'd989;
      109201:data<=16'd1095;
      109202:data<=16'd2232;
      109203:data<=16'd3122;
      109204:data<=16'd2123;
      109205:data<=16'd2173;
      109206:data<=16'd2804;
      109207:data<=16'd1654;
      109208:data<=16'd1694;
      109209:data<=16'd2416;
      109210:data<=16'd1037;
      109211:data<=16'd1844;
      109212:data<=16'd6244;
      109213:data<=16'd7987;
      109214:data<=16'd6915;
      109215:data<=16'd7705;
      109216:data<=16'd8514;
      109217:data<=16'd7673;
      109218:data<=16'd7602;
      109219:data<=16'd7392;
      109220:data<=16'd6388;
      109221:data<=16'd6566;
      109222:data<=16'd7661;
      109223:data<=16'd8428;
      109224:data<=16'd8069;
      109225:data<=16'd7251;
      109226:data<=16'd7151;
      109227:data<=16'd6648;
      109228:data<=16'd6569;
      109229:data<=16'd7846;
      109230:data<=16'd7797;
      109231:data<=16'd6837;
      109232:data<=16'd6686;
      109233:data<=16'd6184;
      109234:data<=16'd5726;
      109235:data<=16'd5876;
      109236:data<=16'd5612;
      109237:data<=16'd4905;
      109238:data<=16'd4604;
      109239:data<=16'd4748;
      109240:data<=16'd4426;
      109241:data<=16'd4676;
      109242:data<=16'd5953;
      109243:data<=16'd5583;
      109244:data<=16'd4467;
      109245:data<=16'd4678;
      109246:data<=16'd4397;
      109247:data<=16'd3588;
      109248:data<=16'd3386;
      109249:data<=16'd3306;
      109250:data<=16'd3040;
      109251:data<=16'd2617;
      109252:data<=16'd2676;
      109253:data<=16'd2560;
      109254:data<=16'd2129;
      109255:data<=16'd2995;
      109256:data<=16'd3386;
      109257:data<=16'd2860;
      109258:data<=16'd3113;
      109259:data<=16'd2523;
      109260:data<=16'd2082;
      109261:data<=16'd2475;
      109262:data<=16'd1651;
      109263:data<=16'd1563;
      109264:data<=16'd881;
      109265:data<=-16'd2883;
      109266:data<=-16'd5797;
      109267:data<=-16'd7183;
      109268:data<=-16'd7988;
      109269:data<=-16'd7307;
      109270:data<=-16'd7110;
      109271:data<=-16'd7235;
      109272:data<=-16'd6972;
      109273:data<=-16'd7315;
      109274:data<=-16'd7200;
      109275:data<=-16'd7127;
      109276:data<=-16'd7194;
      109277:data<=-16'd6625;
      109278:data<=-16'd6905;
      109279:data<=-16'd6836;
      109280:data<=-16'd6056;
      109281:data<=-16'd6705;
      109282:data<=-16'd7673;
      109283:data<=-16'd8143;
      109284:data<=-16'd7999;
      109285:data<=-16'd7353;
      109286:data<=-16'd7555;
      109287:data<=-16'd7438;
      109288:data<=-16'd7065;
      109289:data<=-16'd7157;
      109290:data<=-16'd6466;
      109291:data<=-16'd6746;
      109292:data<=-16'd7245;
      109293:data<=-16'd6117;
      109294:data<=-16'd6734;
      109295:data<=-16'd8184;
      109296:data<=-16'd8006;
      109297:data<=-16'd8109;
      109298:data<=-16'd8144;
      109299:data<=-16'd7802;
      109300:data<=-16'd7370;
      109301:data<=-16'd6555;
      109302:data<=-16'd6669;
      109303:data<=-16'd6652;
      109304:data<=-16'd6304;
      109305:data<=-16'd6684;
      109306:data<=-16'd6166;
      109307:data<=-16'd6379;
      109308:data<=-16'd7712;
      109309:data<=-16'd7439;
      109310:data<=-16'd7529;
      109311:data<=-16'd7447;
      109312:data<=-16'd5406;
      109313:data<=-16'd4789;
      109314:data<=-16'd5213;
      109315:data<=-16'd4740;
      109316:data<=-16'd4896;
      109317:data<=-16'd4610;
      109318:data<=-16'd1632;
      109319:data<=16'd2328;
      109320:data<=16'd3031;
      109321:data<=16'd707;
      109322:data<=-16'd455;
      109323:data<=-16'd472;
      109324:data<=-16'd438;
      109325:data<=-16'd302;
      109326:data<=-16'd996;
      109327:data<=-16'd855;
      109328:data<=-16'd44;
      109329:data<=-16'd660;
      109330:data<=-16'd945;
      109331:data<=-16'd866;
      109332:data<=-16'd1008;
      109333:data<=-16'd528;
      109334:data<=-16'd1371;
      109335:data<=-16'd3066;
      109336:data<=-16'd3539;
      109337:data<=-16'd3392;
      109338:data<=-16'd2823;
      109339:data<=-16'd2816;
      109340:data<=-16'd3315;
      109341:data<=-16'd2990;
      109342:data<=-16'd2895;
      109343:data<=-16'd2836;
      109344:data<=-16'd2535;
      109345:data<=-16'd2622;
      109346:data<=-16'd2314;
      109347:data<=-16'd2581;
      109348:data<=-16'd3313;
      109349:data<=-16'd3529;
      109350:data<=-16'd4232;
      109351:data<=-16'd4011;
      109352:data<=-16'd3331;
      109353:data<=-16'd3949;
      109354:data<=-16'd3821;
      109355:data<=-16'd4061;
      109356:data<=-16'd5357;
      109357:data<=-16'd5327;
      109358:data<=-16'd5201;
      109359:data<=-16'd5153;
      109360:data<=-16'd5124;
      109361:data<=-16'd6282;
      109362:data<=-16'd6536;
      109363:data<=-16'd6159;
      109364:data<=-16'd6249;
      109365:data<=-16'd6032;
      109366:data<=-16'd6050;
      109367:data<=-16'd4996;
      109368:data<=-16'd4347;
      109369:data<=-16'd5312;
      109370:data<=-16'd4194;
      109371:data<=-16'd5221;
      109372:data<=-16'd9879;
      109373:data<=-16'd10278;
      109374:data<=-16'd9627;
      109375:data<=-16'd11717;
      109376:data<=-16'd11436;
      109377:data<=-16'd10248;
      109378:data<=-16'd10305;
      109379:data<=-16'd9806;
      109380:data<=-16'd9157;
      109381:data<=-16'd8511;
      109382:data<=-16'd8479;
      109383:data<=-16'd8645;
      109384:data<=-16'd7834;
      109385:data<=-16'd7110;
      109386:data<=-16'd6032;
      109387:data<=-16'd5883;
      109388:data<=-16'd7870;
      109389:data<=-16'd8094;
      109390:data<=-16'd6821;
      109391:data<=-16'd6532;
      109392:data<=-16'd6037;
      109393:data<=-16'd6003;
      109394:data<=-16'd6235;
      109395:data<=-16'd5485;
      109396:data<=-16'd5007;
      109397:data<=-16'd4755;
      109398:data<=-16'd4546;
      109399:data<=-16'd4429;
      109400:data<=-16'd3826;
      109401:data<=-16'd3738;
      109402:data<=-16'd3627;
      109403:data<=-16'd2767;
      109404:data<=-16'd2705;
      109405:data<=-16'd2807;
      109406:data<=-16'd2191;
      109407:data<=-16'd1999;
      109408:data<=-16'd2014;
      109409:data<=-16'd1439;
      109410:data<=-16'd1043;
      109411:data<=-16'd1343;
      109412:data<=-16'd1054;
      109413:data<=-16'd620;
      109414:data<=-16'd1697;
      109415:data<=-16'd2241;
      109416:data<=-16'd1701;
      109417:data<=-16'd2196;
      109418:data<=-16'd2165;
      109419:data<=-16'd1365;
      109420:data<=-16'd1574;
      109421:data<=-16'd1428;
      109422:data<=-16'd1249;
      109423:data<=-16'd1689;
      109424:data<=16'd420;
      109425:data<=16'd4854;
      109426:data<=16'd6761;
      109427:data<=16'd5136;
      109428:data<=16'd3758;
      109429:data<=16'd3900;
      109430:data<=16'd3817;
      109431:data<=16'd3480;
      109432:data<=16'd3172;
      109433:data<=16'd3043;
      109434:data<=16'd3576;
      109435:data<=16'd3486;
      109436:data<=16'd2908;
      109437:data<=16'd3162;
      109438:data<=16'd3530;
      109439:data<=16'd3833;
      109440:data<=16'd3453;
      109441:data<=16'd1733;
      109442:data<=16'd749;
      109443:data<=16'd1155;
      109444:data<=16'd1409;
      109445:data<=16'd441;
      109446:data<=-16'd1177;
      109447:data<=-16'd1333;
      109448:data<=-16'd644;
      109449:data<=-16'd531;
      109450:data<=-16'd262;
      109451:data<=-16'd273;
      109452:data<=-16'd226;
      109453:data<=-16'd91;
      109454:data<=-16'd1319;
      109455:data<=-16'd1970;
      109456:data<=-16'd1530;
      109457:data<=-16'd1630;
      109458:data<=-16'd990;
      109459:data<=-16'd415;
      109460:data<=-16'd930;
      109461:data<=-16'd993;
      109462:data<=-16'd886;
      109463:data<=-16'd394;
      109464:data<=16'd179;
      109465:data<=-16'd262;
      109466:data<=-16'd268;
      109467:data<=-16'd582;
      109468:data<=-16'd1903;
      109469:data<=-16'd1804;
      109470:data<=-16'd1060;
      109471:data<=-16'd1149;
      109472:data<=-16'd980;
      109473:data<=-16'd500;
      109474:data<=-16'd658;
      109475:data<=-16'd834;
      109476:data<=16'd259;
      109477:data<=-16'd792;
      109478:data<=-16'd5629;
      109479:data<=-16'd7365;
      109480:data<=-16'd5589;
      109481:data<=-16'd5644;
      109482:data<=-16'd5421;
      109483:data<=-16'd4508;
      109484:data<=-16'd4663;
      109485:data<=-16'd4068;
      109486:data<=-16'd3645;
      109487:data<=-16'd3460;
      109488:data<=-16'd2701;
      109489:data<=-16'd2658;
      109490:data<=-16'd1457;
      109491:data<=16'd359;
      109492:data<=16'd281;
      109493:data<=16'd691;
      109494:data<=16'd1996;
      109495:data<=16'd2687;
      109496:data<=16'd3037;
      109497:data<=16'd2924;
      109498:data<=16'd3250;
      109499:data<=16'd3550;
      109500:data<=16'd3068;
      109501:data<=16'd3275;
      109502:data<=16'd3272;
      109503:data<=16'd2807;
      109504:data<=16'd2972;
      109505:data<=16'd2770;
      109506:data<=16'd3212;
      109507:data<=16'd4587;
      109508:data<=16'd5072;
      109509:data<=16'd5275;
      109510:data<=16'd5325;
      109511:data<=16'd5165;
      109512:data<=16'd5225;
      109513:data<=16'd4675;
      109514:data<=16'd4399;
      109515:data<=16'd4572;
      109516:data<=16'd4185;
      109517:data<=16'd4032;
      109518:data<=16'd3750;
      109519:data<=16'd3680;
      109520:data<=16'd4934;
      109521:data<=16'd5985;
      109522:data<=16'd6123;
      109523:data<=16'd5601;
      109524:data<=16'd5257;
      109525:data<=16'd5789;
      109526:data<=16'd5265;
      109527:data<=16'd4816;
      109528:data<=16'd5441;
      109529:data<=16'd4452;
      109530:data<=16'd5333;
      109531:data<=16'd9603;
      109532:data<=16'd11138;
      109533:data<=16'd10918;
      109534:data<=16'd11635;
      109535:data<=16'd10407;
      109536:data<=16'd8663;
      109537:data<=16'd8739;
      109538:data<=16'd8680;
      109539:data<=16'd7840;
      109540:data<=16'd7357;
      109541:data<=16'd7514;
      109542:data<=16'd7400;
      109543:data<=16'd6805;
      109544:data<=16'd6560;
      109545:data<=16'd6475;
      109546:data<=16'd6752;
      109547:data<=16'd7636;
      109548:data<=16'd7935;
      109549:data<=16'd7564;
      109550:data<=16'd7098;
      109551:data<=16'd6402;
      109552:data<=16'd5736;
      109553:data<=16'd5492;
      109554:data<=16'd5645;
      109555:data<=16'd5527;
      109556:data<=16'd5080;
      109557:data<=16'd5056;
      109558:data<=16'd4971;
      109559:data<=16'd4989;
      109560:data<=16'd5923;
      109561:data<=16'd6455;
      109562:data<=16'd6008;
      109563:data<=16'd5620;
      109564:data<=16'd5432;
      109565:data<=16'd5172;
      109566:data<=16'd4695;
      109567:data<=16'd4520;
      109568:data<=16'd4819;
      109569:data<=16'd4555;
      109570:data<=16'd4052;
      109571:data<=16'd3689;
      109572:data<=16'd3143;
      109573:data<=16'd3838;
      109574:data<=16'd5265;
      109575:data<=16'd5092;
      109576:data<=16'd4599;
      109577:data<=16'd4895;
      109578:data<=16'd4593;
      109579:data<=16'd4645;
      109580:data<=16'd5761;
      109581:data<=16'd6102;
      109582:data<=16'd5874;
      109583:data<=16'd4874;
      109584:data<=16'd1011;
      109585:data<=-16'd2406;
      109586:data<=-16'd1312;
      109587:data<=16'd816;
      109588:data<=16'd866;
      109589:data<=16'd350;
      109590:data<=16'd124;
      109591:data<=16'd305;
      109592:data<=16'd579;
      109593:data<=16'd461;
      109594:data<=16'd334;
      109595:data<=16'd49;
      109596:data<=16'd32;
      109597:data<=16'd472;
      109598:data<=16'd194;
      109599:data<=16'd152;
      109600:data<=16'd1175;
      109601:data<=16'd2018;
      109602:data<=16'd2511;
      109603:data<=16'd2379;
      109604:data<=16'd1689;
      109605:data<=16'd1630;
      109606:data<=16'd1704;
      109607:data<=16'd1542;
      109608:data<=16'd1466;
      109609:data<=16'd1090;
      109610:data<=16'd814;
      109611:data<=16'd667;
      109612:data<=16'd564;
      109613:data<=16'd1230;
      109614:data<=16'd2000;
      109615:data<=16'd2325;
      109616:data<=16'd2596;
      109617:data<=16'd2425;
      109618:data<=16'd1858;
      109619:data<=16'd1689;
      109620:data<=16'd2053;
      109621:data<=16'd1902;
      109622:data<=16'd1169;
      109623:data<=16'd1049;
      109624:data<=16'd80;
      109625:data<=-16'd1779;
      109626:data<=-16'd1087;
      109627:data<=16'd605;
      109628:data<=16'd387;
      109629:data<=-16'd18;
      109630:data<=-16'd17;
      109631:data<=16'd6;
      109632:data<=16'd32;
      109633:data<=-16'd332;
      109634:data<=-16'd138;
      109635:data<=-16'd262;
      109636:data<=-16'd496;
      109637:data<=16'd2311;
      109638:data<=16'd5623;
      109639:data<=16'd6332;
      109640:data<=16'd6813;
      109641:data<=16'd7157;
      109642:data<=16'd6516;
      109643:data<=16'd6097;
      109644:data<=16'd5729;
      109645:data<=16'd5180;
      109646:data<=16'd4646;
      109647:data<=16'd4314;
      109648:data<=16'd4252;
      109649:data<=16'd3973;
      109650:data<=16'd4064;
      109651:data<=16'd4027;
      109652:data<=16'd3360;
      109653:data<=16'd4149;
      109654:data<=16'd5198;
      109655:data<=16'd4416;
      109656:data<=16'd3617;
      109657:data<=16'd3033;
      109658:data<=16'd2532;
      109659:data<=16'd2898;
      109660:data<=16'd2643;
      109661:data<=16'd1882;
      109662:data<=16'd1926;
      109663:data<=16'd2240;
      109664:data<=16'd2199;
      109665:data<=16'd1568;
      109666:data<=16'd1783;
      109667:data<=16'd3065;
      109668:data<=16'd3156;
      109669:data<=16'd3341;
      109670:data<=16'd4531;
      109671:data<=16'd4423;
      109672:data<=16'd3745;
      109673:data<=16'd3523;
      109674:data<=16'd3216;
      109675:data<=16'd3198;
      109676:data<=16'd3065;
      109677:data<=16'd2808;
      109678:data<=16'd2493;
      109679:data<=16'd2332;
      109680:data<=16'd3483;
      109681:data<=16'd3856;
      109682:data<=16'd2893;
      109683:data<=16'd3146;
      109684:data<=16'd2585;
      109685:data<=16'd1397;
      109686:data<=16'd2261;
      109687:data<=16'd2184;
      109688:data<=16'd1582;
      109689:data<=16'd2284;
      109690:data<=-16'd321;
      109691:data<=-16'd4958;
      109692:data<=-16'd5859;
      109693:data<=-16'd4872;
      109694:data<=-16'd5045;
      109695:data<=-16'd5429;
      109696:data<=-16'd5366;
      109697:data<=-16'd5292;
      109698:data<=-16'd5162;
      109699:data<=-16'd4911;
      109700:data<=-16'd5215;
      109701:data<=-16'd5404;
      109702:data<=-16'd4743;
      109703:data<=-16'd4784;
      109704:data<=-16'd5219;
      109705:data<=-16'd5012;
      109706:data<=-16'd5667;
      109707:data<=-16'd6616;
      109708:data<=-16'd6369;
      109709:data<=-16'd6123;
      109710:data<=-16'd6261;
      109711:data<=-16'd5908;
      109712:data<=-16'd5448;
      109713:data<=-16'd6031;
      109714:data<=-16'd7326;
      109715:data<=-16'd7783;
      109716:data<=-16'd7691;
      109717:data<=-16'd7450;
      109718:data<=-16'd6768;
      109719:data<=-16'd7438;
      109720:data<=-16'd9110;
      109721:data<=-16'd8945;
      109722:data<=-16'd8009;
      109723:data<=-16'd8061;
      109724:data<=-16'd8066;
      109725:data<=-16'd7665;
      109726:data<=-16'd7262;
      109727:data<=-16'd6951;
      109728:data<=-16'd6892;
      109729:data<=-16'd6960;
      109730:data<=-16'd6590;
      109731:data<=-16'd5694;
      109732:data<=-16'd6078;
      109733:data<=-16'd8067;
      109734:data<=-16'd8467;
      109735:data<=-16'd7380;
      109736:data<=-16'd7621;
      109737:data<=-16'd7665;
      109738:data<=-16'd6663;
      109739:data<=-16'd6871;
      109740:data<=-16'd6957;
      109741:data<=-16'd6181;
      109742:data<=-16'd6472;
      109743:data<=-16'd4605;
      109744:data<=16'd143;
      109745:data<=16'd1016;
      109746:data<=-16'd1256;
      109747:data<=-16'd1348;
      109748:data<=-16'd1307;
      109749:data<=-16'd1844;
      109750:data<=-16'd1151;
      109751:data<=-16'd1140;
      109752:data<=-16'd1580;
      109753:data<=-16'd1239;
      109754:data<=-16'd1184;
      109755:data<=-16'd1152;
      109756:data<=-16'd1266;
      109757:data<=-16'd1500;
      109758:data<=-16'd807;
      109759:data<=-16'd444;
      109760:data<=-16'd920;
      109761:data<=-16'd1237;
      109762:data<=-16'd1613;
      109763:data<=-16'd1771;
      109764:data<=-16'd1503;
      109765:data<=-16'd1122;
      109766:data<=-16'd920;
      109767:data<=-16'd1369;
      109768:data<=-16'd1460;
      109769:data<=-16'd928;
      109770:data<=-16'd772;
      109771:data<=-16'd740;
      109772:data<=-16'd1757;
      109773:data<=-16'd3680;
      109774:data<=-16'd3991;
      109775:data<=-16'd3515;
      109776:data<=-16'd3659;
      109777:data<=-16'd3441;
      109778:data<=-16'd2990;
      109779:data<=-16'd2896;
      109780:data<=-16'd3137;
      109781:data<=-16'd3109;
      109782:data<=-16'd2420;
      109783:data<=-16'd2070;
      109784:data<=-16'd2049;
      109785:data<=-16'd2413;
      109786:data<=-16'd3865;
      109787:data<=-16'd4681;
      109788:data<=-16'd4029;
      109789:data<=-16'd3406;
      109790:data<=-16'd3468;
      109791:data<=-16'd3862;
      109792:data<=-16'd3739;
      109793:data<=-16'd3624;
      109794:data<=-16'd3463;
      109795:data<=-16'd2305;
      109796:data<=-16'd3767;
      109797:data<=-16'd8147;
      109798:data<=-16'd9627;
      109799:data<=-16'd9579;
      109800:data<=-16'd10966;
      109801:data<=-16'd10681;
      109802:data<=-16'd9430;
      109803:data<=-16'd10028;
      109804:data<=-16'd11091;
      109805:data<=-16'd10974;
      109806:data<=-16'd10084;
      109807:data<=-16'd9644;
      109808:data<=-16'd9238;
      109809:data<=-16'd8408;
      109810:data<=-16'd8231;
      109811:data<=-16'd8029;
      109812:data<=-16'd7871;
      109813:data<=-16'd8721;
      109814:data<=-16'd8805;
      109815:data<=-16'd8207;
      109816:data<=-16'd8034;
      109817:data<=-16'd7163;
      109818:data<=-16'd6426;
      109819:data<=-16'd6649;
      109820:data<=-16'd6555;
      109821:data<=-16'd6111;
      109822:data<=-16'd5867;
      109823:data<=-16'd5595;
      109824:data<=-16'd4905;
      109825:data<=-16'd4772;
      109826:data<=-16'd5829;
      109827:data<=-16'd5817;
      109828:data<=-16'd5033;
      109829:data<=-16'd5450;
      109830:data<=-16'd5148;
      109831:data<=-16'd4199;
      109832:data<=-16'd4229;
      109833:data<=-16'd3748;
      109834:data<=-16'd3262;
      109835:data<=-16'd3630;
      109836:data<=-16'd3072;
      109837:data<=-16'd2027;
      109838:data<=-16'd2205;
      109839:data<=-16'd3310;
      109840:data<=-16'd3861;
      109841:data<=-16'd3450;
      109842:data<=-16'd3295;
      109843:data<=-16'd3149;
      109844:data<=-16'd2505;
      109845:data<=-16'd2241;
      109846:data<=-16'd1906;
      109847:data<=-16'd1747;
      109848:data<=-16'd1695;
      109849:data<=16'd1356;
      109850:data<=16'd6138;
      109851:data<=16'd7524;
      109852:data<=16'd6082;
      109853:data<=16'd5066;
      109854:data<=16'd4686;
      109855:data<=16'd4720;
      109856:data<=16'd5139;
      109857:data<=16'd5128;
      109858:data<=16'd4783;
      109859:data<=16'd4660;
      109860:data<=16'd4679;
      109861:data<=16'd4813;
      109862:data<=16'd4532;
      109863:data<=16'd3882;
      109864:data<=16'd4037;
      109865:data<=16'd4034;
      109866:data<=16'd2892;
      109867:data<=16'd2268;
      109868:data<=16'd2221;
      109869:data<=16'd1964;
      109870:data<=16'd2293;
      109871:data<=16'd2878;
      109872:data<=16'd3042;
      109873:data<=16'd3008;
      109874:data<=16'd2870;
      109875:data<=16'd2914;
      109876:data<=16'd3109;
      109877:data<=16'd3004;
      109878:data<=16'd2193;
      109879:data<=16'd943;
      109880:data<=16'd475;
      109881:data<=16'd647;
      109882:data<=16'd702;
      109883:data<=16'd846;
      109884:data<=16'd883;
      109885:data<=16'd1139;
      109886:data<=16'd1475;
      109887:data<=16'd1105;
      109888:data<=16'd1168;
      109889:data<=16'd1539;
      109890:data<=16'd1325;
      109891:data<=16'd1108;
      109892:data<=-16'd340;
      109893:data<=-16'd2432;
      109894:data<=-16'd2516;
      109895:data<=-16'd1847;
      109896:data<=-16'd1824;
      109897:data<=-16'd1820;
      109898:data<=-16'd1532;
      109899:data<=-16'd1139;
      109900:data<=-16'd1266;
      109901:data<=-16'd840;
      109902:data<=-16'd1037;
      109903:data<=-16'd4643;
      109904:data<=-16'd7248;
      109905:data<=-16'd6379;
      109906:data<=-16'd6102;
      109907:data<=-16'd6026;
      109908:data<=-16'd5388;
      109909:data<=-16'd5239;
      109910:data<=-16'd4589;
      109911:data<=-16'd4370;
      109912:data<=-16'd4053;
      109913:data<=-16'd2783;
      109914:data<=-16'd2792;
      109915:data<=-16'd2817;
      109916:data<=-16'd2378;
      109917:data<=-16'd2931;
      109918:data<=-16'd1926;
      109919:data<=16'd80;
      109920:data<=16'd479;
      109921:data<=16'd511;
      109922:data<=16'd728;
      109923:data<=16'd1115;
      109924:data<=16'd1427;
      109925:data<=16'd1245;
      109926:data<=16'd1588;
      109927:data<=16'd1791;
      109928:data<=16'd1710;
      109929:data<=16'd1903;
      109930:data<=16'd1322;
      109931:data<=16'd1844;
      109932:data<=16'd3864;
      109933:data<=16'd4419;
      109934:data<=16'd4428;
      109935:data<=16'd4655;
      109936:data<=16'd4387;
      109937:data<=16'd5077;
      109938:data<=16'd6299;
      109939:data<=16'd6613;
      109940:data<=16'd6263;
      109941:data<=16'd6021;
      109942:data<=16'd6156;
      109943:data<=16'd5838;
      109944:data<=16'd6105;
      109945:data<=16'd7544;
      109946:data<=16'd7834;
      109947:data<=16'd7538;
      109948:data<=16'd7600;
      109949:data<=16'd7274;
      109950:data<=16'd7574;
      109951:data<=16'd7579;
      109952:data<=16'd6898;
      109953:data<=16'd7153;
      109954:data<=16'd6772;
      109955:data<=16'd6816;
      109956:data<=16'd9920;
      109957:data<=16'd12878;
      109958:data<=16'd13788;
      109959:data<=16'd14258;
      109960:data<=16'd14242;
      109961:data<=16'd13650;
      109962:data<=16'd13135;
      109963:data<=16'd12894;
      109964:data<=16'd12513;
      109965:data<=16'd11937;
      109966:data<=16'd11691;
      109967:data<=16'd11165;
      109968:data<=16'd10464;
      109969:data<=16'd10157;
      109970:data<=16'd9471;
      109971:data<=16'd9633;
      109972:data<=16'd11069;
      109973:data<=16'd11035;
      109974:data<=16'd10103;
      109975:data<=16'd10251;
      109976:data<=16'd10111;
      109977:data<=16'd9489;
      109978:data<=16'd9594;
      109979:data<=16'd9283;
      109980:data<=16'd8361;
      109981:data<=16'd8490;
      109982:data<=16'd7887;
      109983:data<=16'd5500;
      109984:data<=16'd5369;
      109985:data<=16'd7344;
      109986:data<=16'd7368;
      109987:data<=16'd6314;
      109988:data<=16'd5902;
      109989:data<=16'd5753;
      109990:data<=16'd5824;
      109991:data<=16'd5733;
      109992:data<=16'd5459;
      109993:data<=16'd4817;
      109994:data<=16'd4121;
      109995:data<=16'd4334;
      109996:data<=16'd4111;
      109997:data<=16'd3729;
      109998:data<=16'd4843;
      109999:data<=16'd5633;
      110000:data<=16'd5342;
      110001:data<=16'd5039;
      110002:data<=16'd4934;
      110003:data<=16'd4930;
      110004:data<=16'd4259;
      110005:data<=16'd3888;
      110006:data<=16'd3856;
      110007:data<=16'd3186;
      110008:data<=16'd3732;
      110009:data<=16'd1933;
      110010:data<=-16'd3695;
      110011:data<=-16'd4231;
      110012:data<=-16'd986;
      110013:data<=-16'd1128;
      110014:data<=-16'd1304;
      110015:data<=-16'd832;
      110016:data<=-16'd1513;
      110017:data<=-16'd1334;
      110018:data<=-16'd1225;
      110019:data<=-16'd1401;
      110020:data<=-16'd1254;
      110021:data<=-16'd1488;
      110022:data<=-16'd1592;
      110023:data<=-16'd2149;
      110024:data<=-16'd1606;
      110025:data<=16'd538;
      110026:data<=16'd643;
      110027:data<=16'd854;
      110028:data<=16'd2591;
      110029:data<=16'd2299;
      110030:data<=16'd1680;
      110031:data<=16'd1895;
      110032:data<=16'd1580;
      110033:data<=16'd1688;
      110034:data<=16'd1283;
      110035:data<=16'd337;
      110036:data<=16'd235;
      110037:data<=16'd699;
      110038:data<=16'd1941;
      110039:data<=16'd2604;
      110040:data<=16'd2047;
      110041:data<=16'd1882;
      110042:data<=16'd1844;
      110043:data<=16'd2023;
      110044:data<=16'd2121;
      110045:data<=16'd1553;
      110046:data<=16'd1535;
      110047:data<=16'd1218;
      110048:data<=16'd795;
      110049:data<=16'd1259;
      110050:data<=16'd1083;
      110051:data<=16'd1654;
      110052:data<=16'd2902;
      110053:data<=16'd2514;
      110054:data<=16'd2273;
      110055:data<=16'd1973;
      110056:data<=16'd1353;
      110057:data<=16'd1786;
      110058:data<=16'd1230;
      110059:data<=16'd866;
      110060:data<=16'd1140;
      110061:data<=-16'd30;
      110062:data<=16'd1926;
      110063:data<=16'd6411;
      110064:data<=16'd7488;
      110065:data<=16'd7621;
      110066:data<=16'd8234;
      110067:data<=16'd7699;
      110068:data<=16'd7322;
      110069:data<=16'd6745;
      110070:data<=16'd6132;
      110071:data<=16'd5843;
      110072:data<=16'd4557;
      110073:data<=16'd3257;
      110074:data<=16'd2543;
      110075:data<=16'd2262;
      110076:data<=16'd2629;
      110077:data<=16'd2714;
      110078:data<=16'd3051;
      110079:data<=16'd3512;
      110080:data<=16'd3125;
      110081:data<=16'd2993;
      110082:data<=16'd2645;
      110083:data<=16'd1927;
      110084:data<=16'd2000;
      110085:data<=16'd1742;
      110086:data<=16'd1434;
      110087:data<=16'd1677;
      110088:data<=16'd1154;
      110089:data<=16'd720;
      110090:data<=16'd1412;
      110091:data<=16'd2514;
      110092:data<=16'd2914;
      110093:data<=16'd2005;
      110094:data<=16'd1491;
      110095:data<=16'd1764;
      110096:data<=16'd1184;
      110097:data<=16'd537;
      110098:data<=16'd406;
      110099:data<=16'd180;
      110100:data<=16'd258;
      110101:data<=16'd343;
      110102:data<=16'd5;
      110103:data<=-16'd214;
      110104:data<=16'd443;
      110105:data<=16'd1689;
      110106:data<=16'd1710;
      110107:data<=16'd845;
      110108:data<=16'd778;
      110109:data<=16'd531;
      110110:data<=16'd164;
      110111:data<=16'd578;
      110112:data<=-16'd42;
      110113:data<=-16'd776;
      110114:data<=16'd282;
      110115:data<=-16'd1125;
      110116:data<=-16'd5597;
      110117:data<=-16'd6583;
      110118:data<=-16'd5027;
      110119:data<=-16'd5400;
      110120:data<=-16'd5359;
      110121:data<=-16'd4955;
      110122:data<=-16'd5867;
      110123:data<=-16'd5679;
      110124:data<=-16'd5333;
      110125:data<=-16'd5829;
      110126:data<=-16'd5312;
      110127:data<=-16'd5192;
      110128:data<=-16'd5371;
      110129:data<=-16'd4619;
      110130:data<=-16'd5059;
      110131:data<=-16'd6457;
      110132:data<=-16'd7168;
      110133:data<=-16'd7071;
      110134:data<=-16'd6323;
      110135:data<=-16'd6384;
      110136:data<=-16'd7109;
      110137:data<=-16'd7195;
      110138:data<=-16'd6936;
      110139:data<=-16'd6384;
      110140:data<=-16'd6370;
      110141:data<=-16'd6646;
      110142:data<=-16'd5824;
      110143:data<=-16'd5867;
      110144:data<=-16'd7124;
      110145:data<=-16'd7482;
      110146:data<=-16'd7521;
      110147:data<=-16'd7561;
      110148:data<=-16'd7228;
      110149:data<=-16'd7050;
      110150:data<=-16'd7142;
      110151:data<=-16'd7232;
      110152:data<=-16'd6649;
      110153:data<=-16'd6267;
      110154:data<=-16'd6672;
      110155:data<=-16'd6340;
      110156:data<=-16'd5993;
      110157:data<=-16'd6376;
      110158:data<=-16'd6987;
      110159:data<=-16'd7794;
      110160:data<=-16'd7442;
      110161:data<=-16'd7611;
      110162:data<=-16'd9148;
      110163:data<=-16'd8549;
      110164:data<=-16'd7968;
      110165:data<=-16'd8425;
      110166:data<=-16'd7421;
      110167:data<=-16'd7905;
      110168:data<=-16'd6839;
      110169:data<=-16'd1547;
      110170:data<=-16'd317;
      110171:data<=-16'd2397;
      110172:data<=-16'd2252;
      110173:data<=-16'd2560;
      110174:data<=-16'd2886;
      110175:data<=-16'd2152;
      110176:data<=-16'd2137;
      110177:data<=-16'd2147;
      110178:data<=-16'd2253;
      110179:data<=-16'd2409;
      110180:data<=-16'd2479;
      110181:data<=-16'd2560;
      110182:data<=-16'd1660;
      110183:data<=-16'd2138;
      110184:data<=-16'd4135;
      110185:data<=-16'd4338;
      110186:data<=-16'd4120;
      110187:data<=-16'd3909;
      110188:data<=-16'd3062;
      110189:data<=-16'd3374;
      110190:data<=-16'd3592;
      110191:data<=-16'd3218;
      110192:data<=-16'd3231;
      110193:data<=-16'd2857;
      110194:data<=-16'd2864;
      110195:data<=-16'd2823;
      110196:data<=-16'd2520;
      110197:data<=-16'd3707;
      110198:data<=-16'd4736;
      110199:data<=-16'd4646;
      110200:data<=-16'd4451;
      110201:data<=-16'd4047;
      110202:data<=-16'd4212;
      110203:data<=-16'd4249;
      110204:data<=-16'd3987;
      110205:data<=-16'd4185;
      110206:data<=-16'd2740;
      110207:data<=-16'd1110;
      110208:data<=-16'd1386;
      110209:data<=-16'd1277;
      110210:data<=-16'd1764;
      110211:data<=-16'd3190;
      110212:data<=-16'd3198;
      110213:data<=-16'd3148;
      110214:data<=-16'd3328;
      110215:data<=-16'd2896;
      110216:data<=-16'd2804;
      110217:data<=-16'd2702;
      110218:data<=-16'd2848;
      110219:data<=-16'd3049;
      110220:data<=-16'd2249;
      110221:data<=-16'd2692;
      110222:data<=-16'd5815;
      110223:data<=-16'd9209;
      110224:data<=-16'd10480;
      110225:data<=-16'd10047;
      110226:data<=-16'd9902;
      110227:data<=-16'd9743;
      110228:data<=-16'd9081;
      110229:data<=-16'd8965;
      110230:data<=-16'd8648;
      110231:data<=-16'd7985;
      110232:data<=-16'd7908;
      110233:data<=-16'd7559;
      110234:data<=-16'd6596;
      110235:data<=-16'd5800;
      110236:data<=-16'd6105;
      110237:data<=-16'd7351;
      110238:data<=-16'd7733;
      110239:data<=-16'd7260;
      110240:data<=-16'd6846;
      110241:data<=-16'd6555;
      110242:data<=-16'd6693;
      110243:data<=-16'd6376;
      110244:data<=-16'd5764;
      110245:data<=-16'd5844;
      110246:data<=-16'd5341;
      110247:data<=-16'd4745;
      110248:data<=-16'd4830;
      110249:data<=-16'd4366;
      110250:data<=-16'd4937;
      110251:data<=-16'd7033;
      110252:data<=-16'd7697;
      110253:data<=-16'd6849;
      110254:data<=-16'd6329;
      110255:data<=-16'd6267;
      110256:data<=-16'd5873;
      110257:data<=-16'd5256;
      110258:data<=-16'd5116;
      110259:data<=-16'd4848;
      110260:data<=-16'd4387;
      110261:data<=-16'd4220;
      110262:data<=-16'd3703;
      110263:data<=-16'd3691;
      110264:data<=-16'd4651;
      110265:data<=-16'd4758;
      110266:data<=-16'd3987;
      110267:data<=-16'd3706;
      110268:data<=-16'd3903;
      110269:data<=-16'd3604;
      110270:data<=-16'd3033;
      110271:data<=-16'd3124;
      110272:data<=-16'd2792;
      110273:data<=-16'd2296;
      110274:data<=-16'd2050;
      110275:data<=16'd1084;
      110276:data<=16'd4672;
      110277:data<=16'd3943;
      110278:data<=16'd2783;
      110279:data<=16'd3268;
      110280:data<=16'd2866;
      110281:data<=16'd2925;
      110282:data<=16'd3697;
      110283:data<=16'd3711;
      110284:data<=16'd3685;
      110285:data<=16'd3680;
      110286:data<=16'd3538;
      110287:data<=16'd3432;
      110288:data<=16'd3294;
      110289:data<=16'd3083;
      110290:data<=16'd2137;
      110291:data<=16'd1340;
      110292:data<=16'd1774;
      110293:data<=16'd2041;
      110294:data<=16'd1894;
      110295:data<=16'd2654;
      110296:data<=16'd4247;
      110297:data<=16'd5204;
      110298:data<=16'd4845;
      110299:data<=16'd4522;
      110300:data<=16'd4572;
      110301:data<=16'd4534;
      110302:data<=16'd4764;
      110303:data<=16'd3871;
      110304:data<=16'd2147;
      110305:data<=16'd1912;
      110306:data<=16'd2033;
      110307:data<=16'd2003;
      110308:data<=16'd2634;
      110309:data<=16'd2537;
      110310:data<=16'd2196;
      110311:data<=16'd2576;
      110312:data<=16'd2641;
      110313:data<=16'd2464;
      110314:data<=16'd2455;
      110315:data<=16'd2663;
      110316:data<=16'd2241;
      110317:data<=16'd546;
      110318:data<=16'd21;
      110319:data<=16'd820;
      110320:data<=16'd887;
      110321:data<=16'd1381;
      110322:data<=16'd1677;
      110323:data<=16'd963;
      110324:data<=16'd1380;
      110325:data<=16'd1500;
      110326:data<=16'd1052;
      110327:data<=16'd2044;
      110328:data<=16'd262;
      110329:data<=-16'd4666;
      110330:data<=-16'd5843;
      110331:data<=-16'd4220;
      110332:data<=-16'd4150;
      110333:data<=-16'd3864;
      110334:data<=-16'd3048;
      110335:data<=-16'd3054;
      110336:data<=-16'd2742;
      110337:data<=-16'd2520;
      110338:data<=-16'd2661;
      110339:data<=-16'd1870;
      110340:data<=-16'd1897;
      110341:data<=-16'd3503;
      110342:data<=-16'd3471;
      110343:data<=-16'd1638;
      110344:data<=-16'd587;
      110345:data<=-16'd347;
      110346:data<=-16'd264;
      110347:data<=-16'd419;
      110348:data<=-16'd315;
      110349:data<=16'd200;
      110350:data<=16'd549;
      110351:data<=16'd476;
      110352:data<=16'd450;
      110353:data<=16'd789;
      110354:data<=16'd886;
      110355:data<=16'd782;
      110356:data<=16'd1600;
      110357:data<=16'd2893;
      110358:data<=16'd3325;
      110359:data<=16'd3418;
      110360:data<=16'd3657;
      110361:data<=16'd3509;
      110362:data<=16'd3515;
      110363:data<=16'd3794;
      110364:data<=16'd3489;
      110365:data<=16'd3183;
      110366:data<=16'd3377;
      110367:data<=16'd3418;
      110368:data<=16'd3418;
      110369:data<=16'd4134;
      110370:data<=16'd5468;
      110371:data<=16'd6047;
      110372:data<=16'd5697;
      110373:data<=16'd5761;
      110374:data<=16'd5726;
      110375:data<=16'd5459;
      110376:data<=16'd5685;
      110377:data<=16'd5153;
      110378:data<=16'd4954;
      110379:data<=16'd5686;
      110380:data<=16'd4784;
      110381:data<=16'd6017;
      110382:data<=16'd11550;
      110383:data<=16'd13984;
      110384:data<=16'd12872;
      110385:data<=16'd13470;
      110386:data<=16'd14066;
      110387:data<=16'd13593;
      110388:data<=16'd13509;
      110389:data<=16'd13056;
      110390:data<=16'd12449;
      110391:data<=16'd12104;
      110392:data<=16'd11837;
      110393:data<=16'd11667;
      110394:data<=16'd10869;
      110395:data<=16'd10272;
      110396:data<=16'd10875;
      110397:data<=16'd11524;
      110398:data<=16'd11544;
      110399:data<=16'd10968;
      110400:data<=16'd10275;
      110401:data<=16'd10067;
      110402:data<=16'd9782;
      110403:data<=16'd9448;
      110404:data<=16'd9266;
      110405:data<=16'd8840;
      110406:data<=16'd8710;
      110407:data<=16'd8552;
      110408:data<=16'd7787;
      110409:data<=16'd7744;
      110410:data<=16'd8733;
      110411:data<=16'd9127;
      110412:data<=16'd8428;
      110413:data<=16'd7961;
      110414:data<=16'd7873;
      110415:data<=16'd7103;
      110416:data<=16'd6784;
      110417:data<=16'd7086;
      110418:data<=16'd6197;
      110419:data<=16'd5635;
      110420:data<=16'd5940;
      110421:data<=16'd5213;
      110422:data<=16'd5230;
      110423:data<=16'd6481;
      110424:data<=16'd6566;
      110425:data<=16'd6075;
      110426:data<=16'd5788;
      110427:data<=16'd5433;
      110428:data<=16'd5136;
      110429:data<=16'd4431;
      110430:data<=16'd3422;
      110431:data<=16'd2008;
      110432:data<=16'd1360;
      110433:data<=16'd2331;
      110434:data<=16'd209;
      110435:data<=-16'd4457;
      110436:data<=-16'd4431;
      110437:data<=-16'd2314;
      110438:data<=-16'd2810;
      110439:data<=-16'd2834;
      110440:data<=-16'd2264;
      110441:data<=-16'd2540;
      110442:data<=-16'd2537;
      110443:data<=-16'd2805;
      110444:data<=-16'd2998;
      110445:data<=-16'd2599;
      110446:data<=-16'd2566;
      110447:data<=-16'd2517;
      110448:data<=-16'd2409;
      110449:data<=-16'd1886;
      110450:data<=-16'd499;
      110451:data<=-16'd62;
      110452:data<=-16'd459;
      110453:data<=-16'd508;
      110454:data<=-16'd866;
      110455:data<=-16'd920;
      110456:data<=-16'd644;
      110457:data<=-16'd1140;
      110458:data<=-16'd1530;
      110459:data<=-16'd1292;
      110460:data<=-16'd1171;
      110461:data<=-16'd1309;
      110462:data<=-16'd890;
      110463:data<=16'd402;
      110464:data<=16'd926;
      110465:data<=16'd493;
      110466:data<=16'd466;
      110467:data<=16'd305;
      110468:data<=16'd177;
      110469:data<=16'd358;
      110470:data<=16'd6;
      110471:data<=16'd165;
      110472:data<=16'd455;
      110473:data<=-16'd338;
      110474:data<=-16'd38;
      110475:data<=16'd1973;
      110476:data<=16'd3639;
      110477:data<=16'd4040;
      110478:data<=16'd3556;
      110479:data<=16'd3372;
      110480:data<=16'd3163;
      110481:data<=16'd2473;
      110482:data<=16'd2426;
      110483:data<=16'd2399;
      110484:data<=16'd2400;
      110485:data<=16'd2725;
      110486:data<=16'd1750;
      110487:data<=16'd2531;
      110488:data<=16'd7090;
      110489:data<=16'd9831;
      110490:data<=16'd9556;
      110491:data<=16'd9364;
      110492:data<=16'd8680;
      110493:data<=16'd7902;
      110494:data<=16'd7662;
      110495:data<=16'd6965;
      110496:data<=16'd6601;
      110497:data<=16'd6454;
      110498:data<=16'd5838;
      110499:data<=16'd5638;
      110500:data<=16'd5187;
      110501:data<=16'd4253;
      110502:data<=16'd4651;
      110503:data<=16'd5871;
      110504:data<=16'd5797;
      110505:data<=16'd4805;
      110506:data<=16'd4679;
      110507:data<=16'd5031;
      110508:data<=16'd4476;
      110509:data<=16'd3767;
      110510:data<=16'd3495;
      110511:data<=16'd3028;
      110512:data<=16'd3039;
      110513:data<=16'd3243;
      110514:data<=16'd2496;
      110515:data<=16'd2450;
      110516:data<=16'd3601;
      110517:data<=16'd3940;
      110518:data<=16'd3692;
      110519:data<=16'd2934;
      110520:data<=16'd948;
      110521:data<=-16'd140;
      110522:data<=16'd368;
      110523:data<=16'd293;
      110524:data<=-16'd318;
      110525:data<=-16'd423;
      110526:data<=-16'd462;
      110527:data<=-16'd682;
      110528:data<=-16'd543;
      110529:data<=16'd88;
      110530:data<=16'd426;
      110531:data<=16'd378;
      110532:data<=16'd409;
      110533:data<=16'd112;
      110534:data<=-16'd428;
      110535:data<=-16'd699;
      110536:data<=-16'd643;
      110537:data<=-16'd596;
      110538:data<=-16'd1162;
      110539:data<=-16'd1287;
      110540:data<=-16'd1850;
      110541:data<=-16'd5711;
      110542:data<=-16'd8836;
      110543:data<=-16'd8040;
      110544:data<=-16'd7802;
      110545:data<=-16'd8044;
      110546:data<=-16'd7028;
      110547:data<=-16'd7201;
      110548:data<=-16'd7570;
      110549:data<=-16'd7318;
      110550:data<=-16'd7298;
      110551:data<=-16'd6736;
      110552:data<=-16'd6981;
      110553:data<=-16'd7330;
      110554:data<=-16'd6363;
      110555:data<=-16'd6857;
      110556:data<=-16'd7988;
      110557:data<=-16'd7908;
      110558:data<=-16'd8170;
      110559:data<=-16'd8217;
      110560:data<=-16'd7808;
      110561:data<=-16'd7427;
      110562:data<=-16'd7083;
      110563:data<=-16'd7530;
      110564:data<=-16'd6813;
      110565:data<=-16'd5018;
      110566:data<=-16'd4851;
      110567:data<=-16'd4816;
      110568:data<=-16'd4978;
      110569:data<=-16'd6260;
      110570:data<=-16'd6586;
      110571:data<=-16'd6737;
      110572:data<=-16'd7045;
      110573:data<=-16'd6458;
      110574:data<=-16'd6197;
      110575:data<=-16'd5917;
      110576:data<=-16'd5580;
      110577:data<=-16'd5745;
      110578:data<=-16'd5435;
      110579:data<=-16'd5197;
      110580:data<=-16'd4921;
      110581:data<=-16'd4954;
      110582:data<=-16'd6363;
      110583:data<=-16'd6758;
      110584:data<=-16'd6185;
      110585:data<=-16'd6166;
      110586:data<=-16'd5732;
      110587:data<=-16'd6008;
      110588:data<=-16'd6156;
      110589:data<=-16'd5095;
      110590:data<=-16'd5142;
      110591:data<=-16'd5107;
      110592:data<=-16'd5092;
      110593:data<=-16'd5322;
      110594:data<=-16'd1721;
      110595:data<=16'd1557;
      110596:data<=16'd65;
      110597:data<=-16'd701;
      110598:data<=-16'd146;
      110599:data<=-16'd846;
      110600:data<=-16'd983;
      110601:data<=-16'd684;
      110602:data<=-16'd670;
      110603:data<=-16'd596;
      110604:data<=-16'd470;
      110605:data<=-16'd429;
      110606:data<=-16'd1037;
      110607:data<=-16'd1071;
      110608:data<=-16'd1155;
      110609:data<=-16'd3535;
      110610:data<=-16'd5150;
      110611:data<=-16'd4540;
      110612:data<=-16'd4460;
      110613:data<=-16'd4443;
      110614:data<=-16'd4115;
      110615:data<=-16'd4320;
      110616:data<=-16'd4121;
      110617:data<=-16'd3659;
      110618:data<=-16'd3845;
      110619:data<=-16'd4209;
      110620:data<=-16'd3874;
      110621:data<=-16'd3765;
      110622:data<=-16'd5046;
      110623:data<=-16'd5662;
      110624:data<=-16'd5075;
      110625:data<=-16'd5160;
      110626:data<=-16'd4911;
      110627:data<=-16'd4387;
      110628:data<=-16'd4667;
      110629:data<=-16'd4197;
      110630:data<=-16'd3700;
      110631:data<=-16'd4463;
      110632:data<=-16'd4596;
      110633:data<=-16'd3820;
      110634:data<=-16'd3835;
      110635:data<=-16'd5049;
      110636:data<=-16'd6032;
      110637:data<=-16'd5601;
      110638:data<=-16'd5103;
      110639:data<=-16'd5133;
      110640:data<=-16'd4576;
      110641:data<=-16'd4165;
      110642:data<=-16'd4267;
      110643:data<=-16'd3971;
      110644:data<=-16'd4081;
      110645:data<=-16'd4237;
      110646:data<=-16'd3268;
      110647:data<=-16'd4792;
      110648:data<=-16'd10266;
      110649:data<=-16'd13151;
      110650:data<=-16'd11617;
      110651:data<=-16'd10645;
      110652:data<=-16'd10220;
      110653:data<=-16'd8810;
      110654:data<=-16'd7862;
      110655:data<=-16'd7156;
      110656:data<=-16'd6351;
      110657:data<=-16'd5973;
      110658:data<=-16'd6072;
      110659:data<=-16'd6166;
      110660:data<=-16'd5157;
      110661:data<=-16'd4825;
      110662:data<=-16'd6369;
      110663:data<=-16'd6652;
      110664:data<=-16'd5830;
      110665:data<=-16'd5762;
      110666:data<=-16'd5325;
      110667:data<=-16'd5048;
      110668:data<=-16'd5142;
      110669:data<=-16'd4532;
      110670:data<=-16'd4052;
      110671:data<=-16'd3956;
      110672:data<=-16'd3855;
      110673:data<=-16'd3692;
      110674:data<=-16'd3753;
      110675:data<=-16'd4525;
      110676:data<=-16'd4589;
      110677:data<=-16'd3915;
      110678:data<=-16'd4026;
      110679:data<=-16'd3785;
      110680:data<=-16'd2999;
      110681:data<=-16'd2658;
      110682:data<=-16'd2582;
      110683:data<=-16'd2699;
      110684:data<=-16'd2153;
      110685:data<=-16'd1600;
      110686:data<=-16'd1994;
      110687:data<=-16'd1971;
      110688:data<=-16'd2370;
      110689:data<=-16'd3092;
      110690:data<=-16'd2373;
      110691:data<=-16'd1985;
      110692:data<=-16'd2082;
      110693:data<=-16'd1442;
      110694:data<=-16'd934;
      110695:data<=-16'd714;
      110696:data<=-16'd887;
      110697:data<=-16'd321;
      110698:data<=-16'd79;
      110699:data<=-16'd2238;
      110700:data<=-16'd763;
      110701:data<=16'd4202;
      110702:data<=16'd4197;
      110703:data<=16'd2837;
      110704:data<=16'd3823;
      110705:data<=16'd3234;
      110706:data<=16'd2939;
      110707:data<=16'd3488;
      110708:data<=16'd3253;
      110709:data<=16'd3808;
      110710:data<=16'd3827;
      110711:data<=16'd3419;
      110712:data<=16'd4064;
      110713:data<=16'd4002;
      110714:data<=16'd3233;
      110715:data<=16'd2290;
      110716:data<=16'd1654;
      110717:data<=16'd2220;
      110718:data<=16'd2473;
      110719:data<=16'd2469;
      110720:data<=16'd2763;
      110721:data<=16'd2649;
      110722:data<=16'd2981;
      110723:data<=16'd3074;
      110724:data<=16'd2701;
      110725:data<=16'd3065;
      110726:data<=16'd2980;
      110727:data<=16'd2397;
      110728:data<=16'd1600;
      110729:data<=16'd549;
      110730:data<=16'd826;
      110731:data<=16'd1304;
      110732:data<=16'd1237;
      110733:data<=16'd1506;
      110734:data<=16'd1061;
      110735:data<=16'd1096;
      110736:data<=16'd1791;
      110737:data<=16'd1381;
      110738:data<=16'd1431;
      110739:data<=16'd1726;
      110740:data<=16'd1481;
      110741:data<=16'd1157;
      110742:data<=-16'd350;
      110743:data<=-16'd353;
      110744:data<=16'd1838;
      110745:data<=16'd2256;
      110746:data<=16'd2288;
      110747:data<=16'd2687;
      110748:data<=16'd2273;
      110749:data<=16'd2840;
      110750:data<=16'd2616;
      110751:data<=16'd1833;
      110752:data<=16'd3080;
      110753:data<=16'd1695;
      110754:data<=-16'd3022;
      110755:data<=-16'd4945;
      110756:data<=-16'd4087;
      110757:data<=-16'd3448;
      110758:data<=-16'd3081;
      110759:data<=-16'd2658;
      110760:data<=-16'd2393;
      110761:data<=-16'd2181;
      110762:data<=-16'd1756;
      110763:data<=-16'd1591;
      110764:data<=-16'd1635;
      110765:data<=-16'd1512;
      110766:data<=-16'd1591;
      110767:data<=-16'd872;
      110768:data<=16'd669;
      110769:data<=16'd1177;
      110770:data<=16'd1222;
      110771:data<=16'd1574;
      110772:data<=16'd1554;
      110773:data<=16'd1466;
      110774:data<=16'd1477;
      110775:data<=16'd1456;
      110776:data<=16'd1679;
      110777:data<=16'd2124;
      110778:data<=16'd2196;
      110779:data<=16'd1694;
      110780:data<=16'd2232;
      110781:data<=16'd3973;
      110782:data<=16'd4811;
      110783:data<=16'd4611;
      110784:data<=16'd4061;
      110785:data<=16'd3920;
      110786:data<=16'd4751;
      110787:data<=16'd4444;
      110788:data<=16'd2713;
      110789:data<=16'd1883;
      110790:data<=16'd2050;
      110791:data<=16'd2452;
      110792:data<=16'd2272;
      110793:data<=16'd1736;
      110794:data<=16'd2880;
      110795:data<=16'd4714;
      110796:data<=16'd4872;
      110797:data<=16'd4220;
      110798:data<=16'd4140;
      110799:data<=16'd4246;
      110800:data<=16'd4159;
      110801:data<=16'd4346;
      110802:data<=16'd4120;
      110803:data<=16'd3529;
      110804:data<=16'd4017;
      110805:data<=16'd3833;
      110806:data<=16'd4287;
      110807:data<=16'd9257;
      110808:data<=16'd13024;
      110809:data<=16'd12000;
      110810:data<=16'd11674;
      110811:data<=16'd11850;
      110812:data<=16'd10751;
      110813:data<=16'd10176;
      110814:data<=16'd9759;
      110815:data<=16'd9734;
      110816:data<=16'd9589;
      110817:data<=16'd8815;
      110818:data<=16'd8977;
      110819:data<=16'd8572;
      110820:data<=16'd8153;
      110821:data<=16'd9605;
      110822:data<=16'd9846;
      110823:data<=16'd9015;
      110824:data<=16'd9041;
      110825:data<=16'd8669;
      110826:data<=16'd8351;
      110827:data<=16'd8025;
      110828:data<=16'd7517;
      110829:data<=16'd7655;
      110830:data<=16'd7156;
      110831:data<=16'd6390;
      110832:data<=16'd6481;
      110833:data<=16'd7464;
      110834:data<=16'd9441;
      110835:data<=16'd9988;
      110836:data<=16'd9075;
      110837:data<=16'd9036;
      110838:data<=16'd8768;
      110839:data<=16'd8436;
      110840:data<=16'd8320;
      110841:data<=16'd7432;
      110842:data<=16'd7028;
      110843:data<=16'd6607;
      110844:data<=16'd6196;
      110845:data<=16'd6555;
      110846:data<=16'd5765;
      110847:data<=16'd5841;
      110848:data<=16'd7473;
      110849:data<=16'd6936;
      110850:data<=16'd6005;
      110851:data<=16'd5973;
      110852:data<=16'd5266;
      110853:data<=16'd5169;
      110854:data<=16'd4974;
      110855:data<=16'd4228;
      110856:data<=16'd4049;
      110857:data<=16'd3852;
      110858:data<=16'd4219;
      110859:data<=16'd2945;
      110860:data<=-16'd1189;
      110861:data<=-16'd2384;
      110862:data<=-16'd937;
      110863:data<=-16'd1574;
      110864:data<=-16'd2073;
      110865:data<=-16'd1504;
      110866:data<=-16'd1767;
      110867:data<=-16'd1780;
      110868:data<=-16'd1583;
      110869:data<=-16'd1874;
      110870:data<=-16'd1780;
      110871:data<=-16'd1870;
      110872:data<=-16'd2394;
      110873:data<=-16'd1798;
      110874:data<=-16'd572;
      110875:data<=-16'd167;
      110876:data<=-16'd187;
      110877:data<=-16'd1033;
      110878:data<=-16'd2663;
      110879:data<=-16'd3178;
      110880:data<=-16'd3043;
      110881:data<=-16'd3162;
      110882:data<=-16'd2958;
      110883:data<=-16'd3066;
      110884:data<=-16'd3203;
      110885:data<=-16'd2899;
      110886:data<=-16'd2736;
      110887:data<=-16'd1806;
      110888:data<=-16'd669;
      110889:data<=-16'd725;
      110890:data<=-16'd1013;
      110891:data<=-16'd1254;
      110892:data<=-16'd1360;
      110893:data<=-16'd1034;
      110894:data<=-16'd1219;
      110895:data<=-16'd1503;
      110896:data<=-16'd1275;
      110897:data<=-16'd1260;
      110898:data<=-16'd1759;
      110899:data<=-16'd2226;
      110900:data<=-16'd1303;
      110901:data<=16'd420;
      110902:data<=16'd726;
      110903:data<=16'd115;
      110904:data<=-16'd97;
      110905:data<=16'd52;
      110906:data<=16'd183;
      110907:data<=-16'd52;
      110908:data<=-16'd462;
      110909:data<=-16'd570;
      110910:data<=16'd83;
      110911:data<=-16'd14;
      110912:data<=-16'd943;
      110913:data<=16'd2394;
      110914:data<=16'd7832;
      110915:data<=16'd8266;
      110916:data<=16'd7319;
      110917:data<=16'd7400;
      110918:data<=16'd5826;
      110919:data<=16'd5433;
      110920:data<=16'd5601;
      110921:data<=16'd4770;
      110922:data<=16'd5792;
      110923:data<=16'd6546;
      110924:data<=16'd6125;
      110925:data<=16'd6314;
      110926:data<=16'd5950;
      110927:data<=16'd6343;
      110928:data<=16'd7019;
      110929:data<=16'd6272;
      110930:data<=16'd6143;
      110931:data<=16'd5783;
      110932:data<=16'd5137;
      110933:data<=16'd5454;
      110934:data<=16'd4764;
      110935:data<=16'd4282;
      110936:data<=16'd4366;
      110937:data<=16'd3500;
      110938:data<=16'd3479;
      110939:data<=16'd3239;
      110940:data<=16'd2880;
      110941:data<=16'd4394;
      110942:data<=16'd4714;
      110943:data<=16'd3935;
      110944:data<=16'd3891;
      110945:data<=16'd3015;
      110946:data<=16'd2581;
      110947:data<=16'd2887;
      110948:data<=16'd2460;
      110949:data<=16'd1967;
      110950:data<=16'd1519;
      110951:data<=16'd1503;
      110952:data<=16'd1489;
      110953:data<=16'd1535;
      110954:data<=16'd2960;
      110955:data<=16'd3162;
      110956:data<=16'd2111;
      110957:data<=16'd2267;
      110958:data<=16'd1824;
      110959:data<=16'd1568;
      110960:data<=16'd1706;
      110961:data<=16'd564;
      110962:data<=16'd728;
      110963:data<=16'd825;
      110964:data<=16'd108;
      110965:data<=16'd1007;
      110966:data<=-16'd1886;
      110967:data<=-16'd7862;
      110968:data<=-16'd8990;
      110969:data<=-16'd8341;
      110970:data<=-16'd9022;
      110971:data<=-16'd8449;
      110972:data<=-16'd7788;
      110973:data<=-16'd7815;
      110974:data<=-16'd7864;
      110975:data<=-16'd7767;
      110976:data<=-16'd7286;
      110977:data<=-16'd7213;
      110978:data<=-16'd7210;
      110979:data<=-16'd7520;
      110980:data<=-16'd8789;
      110981:data<=-16'd9133;
      110982:data<=-16'd8604;
      110983:data<=-16'd8349;
      110984:data<=-16'd8125;
      110985:data<=-16'd8351;
      110986:data<=-16'd8316;
      110987:data<=-16'd7984;
      110988:data<=-16'd8093;
      110989:data<=-16'd7577;
      110990:data<=-16'd7321;
      110991:data<=-16'd7595;
      110992:data<=-16'd6909;
      110993:data<=-16'd7307;
      110994:data<=-16'd8857;
      110995:data<=-16'd8733;
      110996:data<=-16'd8119;
      110997:data<=-16'd8090;
      110998:data<=-16'd7509;
      110999:data<=-16'd7139;
      111000:data<=-16'd7504;
      111001:data<=-16'd7178;
      111002:data<=-16'd6188;
      111003:data<=-16'd6272;
      111004:data<=-16'd6771;
      111005:data<=-16'd6241;
      111006:data<=-16'd6473;
      111007:data<=-16'd7700;
      111008:data<=-16'd7558;
      111009:data<=-16'd6993;
      111010:data<=-16'd7007;
      111011:data<=-16'd5818;
      111012:data<=-16'd4147;
      111013:data<=-16'd3802;
      111014:data<=-16'd3868;
      111015:data<=-16'd3683;
      111016:data<=-16'd3656;
      111017:data<=-16'd3833;
      111018:data<=-16'd4117;
      111019:data<=-16'd2822;
      111020:data<=16'd325;
      111021:data<=16'd1585;
      111022:data<=16'd673;
      111023:data<=16'd613;
      111024:data<=16'd767;
      111025:data<=16'd661;
      111026:data<=16'd930;
      111027:data<=16'd663;
      111028:data<=16'd493;
      111029:data<=16'd538;
      111030:data<=16'd308;
      111031:data<=16'd907;
      111032:data<=16'd849;
      111033:data<=-16'd720;
      111034:data<=-16'd1532;
      111035:data<=-16'd1712;
      111036:data<=-16'd1867;
      111037:data<=-16'd1689;
      111038:data<=-16'd1541;
      111039:data<=-16'd1093;
      111040:data<=-16'd967;
      111041:data<=-16'd1262;
      111042:data<=-16'd1086;
      111043:data<=-16'd1398;
      111044:data<=-16'd1463;
      111045:data<=-16'd693;
      111046:data<=-16'd1548;
      111047:data<=-16'd3304;
      111048:data<=-16'd3600;
      111049:data<=-16'd3054;
      111050:data<=-16'd2670;
      111051:data<=-16'd2593;
      111052:data<=-16'd2689;
      111053:data<=-16'd2884;
      111054:data<=-16'd2775;
      111055:data<=-16'd2722;
      111056:data<=-16'd3988;
      111057:data<=-16'd4623;
      111058:data<=-16'd3714;
      111059:data<=-16'd4334;
      111060:data<=-16'd5852;
      111061:data<=-16'd6305;
      111062:data<=-16'd6094;
      111063:data<=-16'd5213;
      111064:data<=-16'd4998;
      111065:data<=-16'd5297;
      111066:data<=-16'd4930;
      111067:data<=-16'd4889;
      111068:data<=-16'd4299;
      111069:data<=-16'd4065;
      111070:data<=-16'd4702;
      111071:data<=-16'd3227;
      111072:data<=-16'd4558;
      111073:data<=-16'd10730;
      111074:data<=-16'd12675;
      111075:data<=-16'd10903;
      111076:data<=-16'd10895;
      111077:data<=-16'd10627;
      111078:data<=-16'd9903;
      111079:data<=-16'd9458;
      111080:data<=-16'd8818;
      111081:data<=-16'd8624;
      111082:data<=-16'd8076;
      111083:data<=-16'd7577;
      111084:data<=-16'd7257;
      111085:data<=-16'd6642;
      111086:data<=-16'd7611;
      111087:data<=-16'd8639;
      111088:data<=-16'd7803;
      111089:data<=-16'd7260;
      111090:data<=-16'd7163;
      111091:data<=-16'd6862;
      111092:data<=-16'd6451;
      111093:data<=-16'd5771;
      111094:data<=-16'd5585;
      111095:data<=-16'd5304;
      111096:data<=-16'd4811;
      111097:data<=-16'd4525;
      111098:data<=-16'd3780;
      111099:data<=-16'd4297;
      111100:data<=-16'd5184;
      111101:data<=-16'd3685;
      111102:data<=-16'd2573;
      111103:data<=-16'd2690;
      111104:data<=-16'd2147;
      111105:data<=-16'd1994;
      111106:data<=-16'd1770;
      111107:data<=-16'd1061;
      111108:data<=-16'd981;
      111109:data<=-16'd1090;
      111110:data<=-16'd986;
      111111:data<=-16'd326;
      111112:data<=-16'd334;
      111113:data<=-16'd2100;
      111114:data<=-16'd2763;
      111115:data<=-16'd1968;
      111116:data<=-16'd1709;
      111117:data<=-16'd1253;
      111118:data<=-16'd749;
      111119:data<=-16'd506;
      111120:data<=-16'd206;
      111121:data<=-16'd147;
      111122:data<=16'd469;
      111123:data<=16'd619;
      111124:data<=-16'd61;
      111125:data<=16'd1560;
      111126:data<=16'd4463;
      111127:data<=16'd5356;
      111128:data<=16'd5086;
      111129:data<=16'd4949;
      111130:data<=16'd4796;
      111131:data<=16'd4666;
      111132:data<=16'd4889;
      111133:data<=16'd5207;
      111134:data<=16'd5089;
      111135:data<=16'd5100;
      111136:data<=16'd5086;
      111137:data<=16'd4808;
      111138:data<=16'd4971;
      111139:data<=16'd4290;
      111140:data<=16'd2619;
      111141:data<=16'd2085;
      111142:data<=16'd2367;
      111143:data<=16'd2476;
      111144:data<=16'd2056;
      111145:data<=16'd1019;
      111146:data<=16'd616;
      111147:data<=16'd792;
      111148:data<=16'd825;
      111149:data<=16'd848;
      111150:data<=16'd798;
      111151:data<=16'd1204;
      111152:data<=16'd926;
      111153:data<=-16'd886;
      111154:data<=-16'd1456;
      111155:data<=-16'd717;
      111156:data<=-16'd738;
      111157:data<=-16'd848;
      111158:data<=-16'd746;
      111159:data<=-16'd484;
      111160:data<=-16'd5;
      111161:data<=-16'd59;
      111162:data<=-16'd271;
      111163:data<=-16'd129;
      111164:data<=16'd297;
      111165:data<=16'd112;
      111166:data<=-16'd1343;
      111167:data<=-16'd1961;
      111168:data<=-16'd1504;
      111169:data<=-16'd1586;
      111170:data<=-16'd1163;
      111171:data<=-16'd832;
      111172:data<=-16'd1397;
      111173:data<=-16'd1213;
      111174:data<=-16'd866;
      111175:data<=-16'd805;
      111176:data<=-16'd255;
      111177:data<=16'd200;
      111178:data<=-16'd511;
      111179:data<=-16'd3670;
      111180:data<=-16'd6623;
      111181:data<=-16'd6103;
      111182:data<=-16'd5345;
      111183:data<=-16'd5389;
      111184:data<=-16'd4513;
      111185:data<=-16'd4529;
      111186:data<=-16'd4494;
      111187:data<=-16'd3626;
      111188:data<=-16'd3750;
      111189:data<=-16'd2784;
      111190:data<=-16'd829;
      111191:data<=-16'd411;
      111192:data<=16'd355;
      111193:data<=16'd1753;
      111194:data<=16'd2043;
      111195:data<=16'd2153;
      111196:data<=16'd2311;
      111197:data<=16'd1947;
      111198:data<=16'd1933;
      111199:data<=16'd2575;
      111200:data<=16'd2784;
      111201:data<=16'd2544;
      111202:data<=16'd2887;
      111203:data<=16'd3019;
      111204:data<=16'd2705;
      111205:data<=16'd3513;
      111206:data<=16'd4801;
      111207:data<=16'd5307;
      111208:data<=16'd5197;
      111209:data<=16'd4758;
      111210:data<=16'd4683;
      111211:data<=16'd4749;
      111212:data<=16'd4687;
      111213:data<=16'd4943;
      111214:data<=16'd4802;
      111215:data<=16'd4614;
      111216:data<=16'd4713;
      111217:data<=16'd4435;
      111218:data<=16'd5336;
      111219:data<=16'd6745;
      111220:data<=16'd6488;
      111221:data<=16'd6387;
      111222:data<=16'd6716;
      111223:data<=16'd6343;
      111224:data<=16'd6270;
      111225:data<=16'd6150;
      111226:data<=16'd6015;
      111227:data<=16'd6105;
      111228:data<=16'd5788;
      111229:data<=16'd6099;
      111230:data<=16'd5874;
      111231:data<=16'd5468;
      111232:data<=16'd9260;
      111233:data<=16'd13518;
      111234:data<=16'd12637;
      111235:data<=16'd10833;
      111236:data<=16'd10654;
      111237:data<=16'd10009;
      111238:data<=16'd9636;
      111239:data<=16'd9662;
      111240:data<=16'd8907;
      111241:data<=16'd8229;
      111242:data<=16'd8483;
      111243:data<=16'd8516;
      111244:data<=16'd7618;
      111245:data<=16'd7861;
      111246:data<=16'd9362;
      111247:data<=16'd9230;
      111248:data<=16'd8273;
      111249:data<=16'd8226;
      111250:data<=16'd7888;
      111251:data<=16'd7594;
      111252:data<=16'd7659;
      111253:data<=16'd7100;
      111254:data<=16'd6713;
      111255:data<=16'd6660;
      111256:data<=16'd6531;
      111257:data<=16'd6978;
      111258:data<=16'd7758;
      111259:data<=16'd8918;
      111260:data<=16'd9962;
      111261:data<=16'd9404;
      111262:data<=16'd8560;
      111263:data<=16'd8205;
      111264:data<=16'd7224;
      111265:data<=16'd6966;
      111266:data<=16'd7426;
      111267:data<=16'd6855;
      111268:data<=16'd6355;
      111269:data<=16'd6169;
      111270:data<=16'd5438;
      111271:data<=16'd5448;
      111272:data<=16'd6394;
      111273:data<=16'd6780;
      111274:data<=16'd6316;
      111275:data<=16'd6018;
      111276:data<=16'd6032;
      111277:data<=16'd5241;
      111278:data<=16'd4511;
      111279:data<=16'd4810;
      111280:data<=16'd4593;
      111281:data<=16'd4003;
      111282:data<=16'd3554;
      111283:data<=16'd2781;
      111284:data<=16'd3001;
      111285:data<=16'd2969;
      111286:data<=16'd1136;
      111287:data<=16'd503;
      111288:data<=16'd948;
      111289:data<=16'd420;
      111290:data<=16'd461;
      111291:data<=16'd743;
      111292:data<=16'd312;
      111293:data<=16'd230;
      111294:data<=16'd130;
      111295:data<=-16'd86;
      111296:data<=-16'd285;
      111297:data<=-16'd802;
      111298:data<=-16'd281;
      111299:data<=16'd1148;
      111300:data<=16'd1588;
      111301:data<=16'd1209;
      111302:data<=16'd1014;
      111303:data<=16'd1025;
      111304:data<=16'd693;
      111305:data<=16'd293;
      111306:data<=16'd359;
      111307:data<=16'd76;
      111308:data<=-16'd274;
      111309:data<=-16'd138;
      111310:data<=-16'd356;
      111311:data<=16'd140;
      111312:data<=16'd1591;
      111313:data<=16'd1807;
      111314:data<=16'd1240;
      111315:data<=16'd1040;
      111316:data<=16'd820;
      111317:data<=16'd704;
      111318:data<=16'd594;
      111319:data<=16'd578;
      111320:data<=16'd570;
      111321:data<=16'd127;
      111322:data<=-16'd41;
      111323:data<=-16'd152;
      111324:data<=-16'd400;
      111325:data<=16'd321;
      111326:data<=16'd1168;
      111327:data<=16'd1368;
      111328:data<=16'd1368;
      111329:data<=16'd990;
      111330:data<=16'd826;
      111331:data<=16'd799;
      111332:data<=16'd614;
      111333:data<=16'd723;
      111334:data<=16'd202;
      111335:data<=-16'd17;
      111336:data<=16'd226;
      111337:data<=-16'd920;
      111338:data<=16'd722;
      111339:data<=16'd5524;
      111340:data<=16'd6125;
      111341:data<=16'd4538;
      111342:data<=16'd5040;
      111343:data<=16'd4419;
      111344:data<=16'd3498;
      111345:data<=16'd3795;
      111346:data<=16'd3192;
      111347:data<=16'd2725;
      111348:data<=16'd2778;
      111349:data<=16'd2229;
      111350:data<=16'd2021;
      111351:data<=16'd2573;
      111352:data<=16'd3686;
      111353:data<=16'd4184;
      111354:data<=16'd3256;
      111355:data<=16'd2717;
      111356:data<=16'd2696;
      111357:data<=16'd2253;
      111358:data<=16'd2120;
      111359:data<=16'd1992;
      111360:data<=16'd1688;
      111361:data<=16'd1680;
      111362:data<=16'd1404;
      111363:data<=16'd866;
      111364:data<=16'd958;
      111365:data<=16'd1983;
      111366:data<=16'd2596;
      111367:data<=16'd2062;
      111368:data<=16'd1932;
      111369:data<=16'd2041;
      111370:data<=16'd1712;
      111371:data<=16'd1757;
      111372:data<=16'd1158;
      111373:data<=16'd265;
      111374:data<=16'd444;
      111375:data<=16'd187;
      111376:data<=-16'd187;
      111377:data<=16'd217;
      111378:data<=16'd472;
      111379:data<=16'd1108;
      111380:data<=16'd1374;
      111381:data<=16'd875;
      111382:data<=16'd1104;
      111383:data<=16'd732;
      111384:data<=-16'd99;
      111385:data<=16'd168;
      111386:data<=-16'd26;
      111387:data<=-16'd672;
      111388:data<=-16'd1155;
      111389:data<=-16'd1463;
      111390:data<=-16'd693;
      111391:data<=-16'd1713;
      111392:data<=-16'd5186;
      111393:data<=-16'd6252;
      111394:data<=-16'd5406;
      111395:data<=-16'd5551;
      111396:data<=-16'd5550;
      111397:data<=-16'd5318;
      111398:data<=-16'd5409;
      111399:data<=-16'd5244;
      111400:data<=-16'd5274;
      111401:data<=-16'd5618;
      111402:data<=-16'd5406;
      111403:data<=-16'd4980;
      111404:data<=-16'd5650;
      111405:data<=-16'd6787;
      111406:data<=-16'd7074;
      111407:data<=-16'd7112;
      111408:data<=-16'd6857;
      111409:data<=-16'd6132;
      111410:data<=-16'd6099;
      111411:data<=-16'd6326;
      111412:data<=-16'd6346;
      111413:data<=-16'd6522;
      111414:data<=-16'd6302;
      111415:data<=-16'd6188;
      111416:data<=-16'd6405;
      111417:data<=-16'd6354;
      111418:data<=-16'd6834;
      111419:data<=-16'd7503;
      111420:data<=-16'd7515;
      111421:data<=-16'd7567;
      111422:data<=-16'd7485;
      111423:data<=-16'd6937;
      111424:data<=-16'd6505;
      111425:data<=-16'd6546;
      111426:data<=-16'd6587;
      111427:data<=-16'd5896;
      111428:data<=-16'd5568;
      111429:data<=-16'd5883;
      111430:data<=-16'd5430;
      111431:data<=-16'd5773;
      111432:data<=-16'd7347;
      111433:data<=-16'd7353;
      111434:data<=-16'd6619;
      111435:data<=-16'd6702;
      111436:data<=-16'd6123;
      111437:data<=-16'd5200;
      111438:data<=-16'd5277;
      111439:data<=-16'd5580;
      111440:data<=-16'd5257;
      111441:data<=-16'd4739;
      111442:data<=-16'd4620;
      111443:data<=-16'd4746;
      111444:data<=-16'd4196;
      111445:data<=-16'd2746;
      111446:data<=-16'd1864;
      111447:data<=-16'd1879;
      111448:data<=-16'd1653;
      111449:data<=-16'd1709;
      111450:data<=-16'd1888;
      111451:data<=-16'd1425;
      111452:data<=-16'd1527;
      111453:data<=-16'd1509;
      111454:data<=-16'd963;
      111455:data<=-16'd1457;
      111456:data<=-16'd1445;
      111457:data<=-16'd1284;
      111458:data<=-16'd2933;
      111459:data<=-16'd3580;
      111460:data<=-16'd3022;
      111461:data<=-16'd3386;
      111462:data<=-16'd3287;
      111463:data<=-16'd2852;
      111464:data<=-16'd2787;
      111465:data<=-16'd2602;
      111466:data<=-16'd2623;
      111467:data<=-16'd2331;
      111468:data<=-16'd2068;
      111469:data<=-16'd2194;
      111470:data<=-16'd2256;
      111471:data<=-16'd3380;
      111472:data<=-16'd4297;
      111473:data<=-16'd3803;
      111474:data<=-16'd3850;
      111475:data<=-16'd3723;
      111476:data<=-16'd2942;
      111477:data<=-16'd2779;
      111478:data<=-16'd2732;
      111479:data<=-16'd3075;
      111480:data<=-16'd3243;
      111481:data<=-16'd2640;
      111482:data<=-16'd2575;
      111483:data<=-16'd2419;
      111484:data<=-16'd2795;
      111485:data<=-16'd4240;
      111486:data<=-16'd4323;
      111487:data<=-16'd4217;
      111488:data<=-16'd4684;
      111489:data<=-16'd3990;
      111490:data<=-16'd3755;
      111491:data<=-16'd4055;
      111492:data<=-16'd3667;
      111493:data<=-16'd3617;
      111494:data<=-16'd3548;
      111495:data<=-16'd2901;
      111496:data<=-16'd2103;
      111497:data<=-16'd3292;
      111498:data<=-16'd7611;
      111499:data<=-16'd10093;
      111500:data<=-16'd9103;
      111501:data<=-16'd8454;
      111502:data<=-16'd7874;
      111503:data<=-16'd7288;
      111504:data<=-16'd7530;
      111505:data<=-16'd7169;
      111506:data<=-16'd6858;
      111507:data<=-16'd6730;
      111508:data<=-16'd5952;
      111509:data<=-16'd5550;
      111510:data<=-16'd5805;
      111511:data<=-16'd6739;
      111512:data<=-16'd7300;
      111513:data<=-16'd6511;
      111514:data<=-16'd6043;
      111515:data<=-16'd5630;
      111516:data<=-16'd4930;
      111517:data<=-16'd5184;
      111518:data<=-16'd5165;
      111519:data<=-16'd4625;
      111520:data<=-16'd4319;
      111521:data<=-16'd3824;
      111522:data<=-16'd3709;
      111523:data<=-16'd3751;
      111524:data<=-16'd4114;
      111525:data<=-16'd5048;
      111526:data<=-16'd4986;
      111527:data<=-16'd4816;
      111528:data<=-16'd4969;
      111529:data<=-16'd4134;
      111530:data<=-16'd3682;
      111531:data<=-16'd3577;
      111532:data<=-16'd3102;
      111533:data<=-16'd3057;
      111534:data<=-16'd2717;
      111535:data<=-16'd2425;
      111536:data<=-16'd2361;
      111537:data<=-16'd2249;
      111538:data<=-16'd3541;
      111539:data<=-16'd4205;
      111540:data<=-16'd3112;
      111541:data<=-16'd3074;
      111542:data<=-16'd2919;
      111543:data<=-16'd1812;
      111544:data<=-16'd1574;
      111545:data<=-16'd1395;
      111546:data<=-16'd1196;
      111547:data<=-16'd1257;
      111548:data<=-16'd617;
      111549:data<=-16'd294;
      111550:data<=-16'd855;
      111551:data<=-16'd570;
      111552:data<=16'd1359;
      111553:data<=16'd2711;
      111554:data<=16'd2184;
      111555:data<=16'd2129;
      111556:data<=16'd2634;
      111557:data<=16'd2355;
      111558:data<=16'd2705;
      111559:data<=16'd3115;
      111560:data<=16'd2587;
      111561:data<=16'd2617;
      111562:data<=16'd3099;
      111563:data<=16'd2867;
      111564:data<=16'd1641;
      111565:data<=16'd578;
      111566:data<=16'd725;
      111567:data<=16'd807;
      111568:data<=16'd831;
      111569:data<=16'd1293;
      111570:data<=16'd1248;
      111571:data<=16'd1450;
      111572:data<=16'd1880;
      111573:data<=16'd1902;
      111574:data<=16'd2126;
      111575:data<=16'd1961;
      111576:data<=16'd1754;
      111577:data<=16'd1340;
      111578:data<=-16'd173;
      111579:data<=-16'd385;
      111580:data<=16'd475;
      111581:data<=16'd344;
      111582:data<=16'd540;
      111583:data<=16'd804;
      111584:data<=16'd629;
      111585:data<=16'd772;
      111586:data<=16'd769;
      111587:data<=16'd1043;
      111588:data<=16'd1378;
      111589:data<=16'd1389;
      111590:data<=16'd1008;
      111591:data<=-16'd459;
      111592:data<=-16'd758;
      111593:data<=-16'd15;
      111594:data<=-16'd710;
      111595:data<=-16'd719;
      111596:data<=-16'd356;
      111597:data<=-16'd647;
      111598:data<=16'd99;
      111599:data<=16'd79;
      111600:data<=-16'd18;
      111601:data<=16'd679;
      111602:data<=16'd143;
      111603:data<=16'd707;
      111604:data<=16'd249;
      111605:data<=-16'd3228;
      111606:data<=-16'd3620;
      111607:data<=-16'd2608;
      111608:data<=-16'd3257;
      111609:data<=-16'd2469;
      111610:data<=-16'd1994;
      111611:data<=-16'd1847;
      111612:data<=-16'd1017;
      111613:data<=-16'd1577;
      111614:data<=-16'd1428;
      111615:data<=-16'd814;
      111616:data<=-16'd646;
      111617:data<=16'd1115;
      111618:data<=16'd1770;
      111619:data<=16'd1354;
      111620:data<=16'd2106;
      111621:data<=16'd2033;
      111622:data<=16'd2041;
      111623:data<=16'd2308;
      111624:data<=16'd1876;
      111625:data<=16'd2375;
      111626:data<=16'd2391;
      111627:data<=16'd2033;
      111628:data<=16'd2610;
      111629:data<=16'd2607;
      111630:data<=16'd3469;
      111631:data<=16'd4925;
      111632:data<=16'd4824;
      111633:data<=16'd4666;
      111634:data<=16'd4498;
      111635:data<=16'd4370;
      111636:data<=16'd4645;
      111637:data<=16'd4237;
      111638:data<=16'd4373;
      111639:data<=16'd4622;
      111640:data<=16'd4297;
      111641:data<=16'd4476;
      111642:data<=16'd3847;
      111643:data<=16'd4246;
      111644:data<=16'd6516;
      111645:data<=16'd6576;
      111646:data<=16'd5820;
      111647:data<=16'd6058;
      111648:data<=16'd5796;
      111649:data<=16'd5902;
      111650:data<=16'd5715;
      111651:data<=16'd5328;
      111652:data<=16'd5755;
      111653:data<=16'd5507;
      111654:data<=16'd5604;
      111655:data<=16'd5618;
      111656:data<=16'd4843;
      111657:data<=16'd7336;
      111658:data<=16'd11157;
      111659:data<=16'd11571;
      111660:data<=16'd10756;
      111661:data<=16'd10343;
      111662:data<=16'd9878;
      111663:data<=16'd9777;
      111664:data<=16'd9691;
      111665:data<=16'd9461;
      111666:data<=16'd9154;
      111667:data<=16'd8906;
      111668:data<=16'd8589;
      111669:data<=16'd8296;
      111670:data<=16'd9010;
      111671:data<=16'd9685;
      111672:data<=16'd9374;
      111673:data<=16'd9095;
      111674:data<=16'd8511;
      111675:data<=16'd7906;
      111676:data<=16'd7911;
      111677:data<=16'd7685;
      111678:data<=16'd7465;
      111679:data<=16'd7269;
      111680:data<=16'd6857;
      111681:data<=16'd6549;
      111682:data<=16'd6203;
      111683:data<=16'd6860;
      111684:data<=16'd8113;
      111685:data<=16'd8017;
      111686:data<=16'd7532;
      111687:data<=16'd7426;
      111688:data<=16'd7183;
      111689:data<=16'd6862;
      111690:data<=16'd6153;
      111691:data<=16'd5638;
      111692:data<=16'd5650;
      111693:data<=16'd5580;
      111694:data<=16'd5359;
      111695:data<=16'd4880;
      111696:data<=16'd5318;
      111697:data<=16'd6721;
      111698:data<=16'd6771;
      111699:data<=16'd5967;
      111700:data<=16'd5612;
      111701:data<=16'd5292;
      111702:data<=16'd4934;
      111703:data<=16'd4353;
      111704:data<=16'd3955;
      111705:data<=16'd3745;
      111706:data<=16'd3415;
      111707:data<=16'd3466;
      111708:data<=16'd3301;
      111709:data<=16'd3718;
      111710:data<=16'd4194;
      111711:data<=16'd1859;
      111712:data<=16'd130;
      111713:data<=16'd848;
      111714:data<=16'd320;
      111715:data<=-16'd15;
      111716:data<=16'd329;
      111717:data<=-16'd238;
      111718:data<=-16'd129;
      111719:data<=-16'd426;
      111720:data<=-16'd793;
      111721:data<=-16'd61;
      111722:data<=-16'd449;
      111723:data<=-16'd129;
      111724:data<=16'd1337;
      111725:data<=16'd1281;
      111726:data<=16'd1171;
      111727:data<=16'd958;
      111728:data<=16'd494;
      111729:data<=16'd826;
      111730:data<=16'd400;
      111731:data<=16'd206;
      111732:data<=16'd353;
      111733:data<=-16'd378;
      111734:data<=-16'd256;
      111735:data<=-16'd344;
      111736:data<=-16'd149;
      111737:data<=16'd1783;
      111738:data<=16'd1815;
      111739:data<=16'd873;
      111740:data<=16'd1140;
      111741:data<=16'd560;
      111742:data<=16'd183;
      111743:data<=16'd346;
      111744:data<=16'd249;
      111745:data<=16'd388;
      111746:data<=-16'd241;
      111747:data<=-16'd619;
      111748:data<=-16'd529;
      111749:data<=-16'd362;
      111750:data<=16'd1471;
      111751:data<=16'd1992;
      111752:data<=16'd778;
      111753:data<=16'd1207;
      111754:data<=16'd1125;
      111755:data<=16'd678;
      111756:data<=16'd1163;
      111757:data<=16'd564;
      111758:data<=16'd183;
      111759:data<=16'd114;
      111760:data<=-16'd206;
      111761:data<=16'd36;
      111762:data<=-16'd487;
      111763:data<=16'd1098;
      111764:data<=16'd5107;
      111765:data<=16'd5818;
      111766:data<=16'd4857;
      111767:data<=16'd4811;
      111768:data<=16'd4384;
      111769:data<=16'd4417;
      111770:data<=16'd3900;
      111771:data<=16'd2971;
      111772:data<=16'd3163;
      111773:data<=16'd3030;
      111774:data<=16'd2911;
      111775:data<=16'd2831;
      111776:data<=16'd2543;
      111777:data<=16'd3676;
      111778:data<=16'd4340;
      111779:data<=16'd3577;
      111780:data<=16'd3113;
      111781:data<=16'd2544;
      111782:data<=16'd2220;
      111783:data<=16'd2250;
      111784:data<=16'd1956;
      111785:data<=16'd1727;
      111786:data<=16'd1310;
      111787:data<=16'd1216;
      111788:data<=16'd1268;
      111789:data<=16'd1142;
      111790:data<=16'd2179;
      111791:data<=16'd2737;
      111792:data<=16'd2265;
      111793:data<=16'd2431;
      111794:data<=16'd1770;
      111795:data<=16'd1118;
      111796:data<=16'd1495;
      111797:data<=16'd980;
      111798:data<=16'd711;
      111799:data<=16'd869;
      111800:data<=16'd271;
      111801:data<=16'd132;
      111802:data<=16'd637;
      111803:data<=16'd1721;
      111804:data<=16'd2258;
      111805:data<=16'd1374;
      111806:data<=16'd1206;
      111807:data<=16'd1139;
      111808:data<=16'd614;
      111809:data<=16'd751;
      111810:data<=-16'd80;
      111811:data<=-16'd600;
      111812:data<=16'd73;
      111813:data<=-16'd745;
      111814:data<=-16'd1242;
      111815:data<=-16'd438;
      111816:data<=-16'd1158;
      111817:data<=-16'd3498;
      111818:data<=-16'd5647;
      111819:data<=-16'd5927;
      111820:data<=-16'd5462;
      111821:data<=-16'd5624;
      111822:data<=-16'd5124;
      111823:data<=-16'd5369;
      111824:data<=-16'd6202;
      111825:data<=-16'd5491;
      111826:data<=-16'd5453;
      111827:data<=-16'd5682;
      111828:data<=-16'd5045;
      111829:data<=-16'd5935;
      111830:data<=-16'd7115;
      111831:data<=-16'd7306;
      111832:data<=-16'd7251;
      111833:data<=-16'd6827;
      111834:data<=-16'd6907;
      111835:data<=-16'd6596;
      111836:data<=-16'd6040;
      111837:data<=-16'd6813;
      111838:data<=-16'd6821;
      111839:data<=-16'd6378;
      111840:data<=-16'd6387;
      111841:data<=-16'd5579;
      111842:data<=-16'd6390;
      111843:data<=-16'd8138;
      111844:data<=-16'd7877;
      111845:data<=-16'd7606;
      111846:data<=-16'd7539;
      111847:data<=-16'd7054;
      111848:data<=-16'd7086;
      111849:data<=-16'd6953;
      111850:data<=-16'd6928;
      111851:data<=-16'd6763;
      111852:data<=-16'd6208;
      111853:data<=-16'd6273;
      111854:data<=-16'd5937;
      111855:data<=-16'd6035;
      111856:data<=-16'd7454;
      111857:data<=-16'd7811;
      111858:data<=-16'd7498;
      111859:data<=-16'd7357;
      111860:data<=-16'd6871;
      111861:data<=-16'd6746;
      111862:data<=-16'd6602;
      111863:data<=-16'd6496;
      111864:data<=-16'd6267;
      111865:data<=-16'd5497;
      111866:data<=-16'd5691;
      111867:data<=-16'd5715;
      111868:data<=-16'd5397;
      111869:data<=-16'd6323;
      111870:data<=-16'd5259;
      111871:data<=-16'd2679;
      111872:data<=-16'd2367;
      111873:data<=-16'd2399;
      111874:data<=-16'd2029;
      111875:data<=-16'd2149;
      111876:data<=-16'd2009;
      111877:data<=-16'd2188;
      111878:data<=-16'd2159;
      111879:data<=-16'd1811;
      111880:data<=-16'd1886;
      111881:data<=-16'd1598;
      111882:data<=-16'd2187;
      111883:data<=-16'd3606;
      111884:data<=-16'd3645;
      111885:data<=-16'd3395;
      111886:data<=-16'd3539;
      111887:data<=-16'd3297;
      111888:data<=-16'd3058;
      111889:data<=-16'd2861;
      111890:data<=-16'd2833;
      111891:data<=-16'd2772;
      111892:data<=-16'd2573;
      111893:data<=-16'd2549;
      111894:data<=-16'd2149;
      111895:data<=-16'd2479;
      111896:data<=-16'd3941;
      111897:data<=-16'd4364;
      111898:data<=-16'd3982;
      111899:data<=-16'd3664;
      111900:data<=-16'd3386;
      111901:data<=-16'd3592;
      111902:data<=-16'd3328;
      111903:data<=-16'd2848;
      111904:data<=-16'd3080;
      111905:data<=-16'd2999;
      111906:data<=-16'd2855;
      111907:data<=-16'd2778;
      111908:data<=-16'd2590;
      111909:data<=-16'd3526;
      111910:data<=-16'd4400;
      111911:data<=-16'd4046;
      111912:data<=-16'd3800;
      111913:data<=-16'd3685;
      111914:data<=-16'd3513;
      111915:data<=-16'd3548;
      111916:data<=-16'd3339;
      111917:data<=-16'd3115;
      111918:data<=-16'd2921;
      111919:data<=-16'd2758;
      111920:data<=-16'd2980;
      111921:data<=-16'd2751;
      111922:data<=-16'd2576;
      111923:data<=-16'd4905;
      111924:data<=-16'd8310;
      111925:data<=-16'd8810;
      111926:data<=-16'd7664;
      111927:data<=-16'd7553;
      111928:data<=-16'd7103;
      111929:data<=-16'd6614;
      111930:data<=-16'd6905;
      111931:data<=-16'd6184;
      111932:data<=-16'd5565;
      111933:data<=-16'd5762;
      111934:data<=-16'd5142;
      111935:data<=-16'd5327;
      111936:data<=-16'd6549;
      111937:data<=-16'd6639;
      111938:data<=-16'd6122;
      111939:data<=-16'd5756;
      111940:data<=-16'd5560;
      111941:data<=-16'd5131;
      111942:data<=-16'd4384;
      111943:data<=-16'd4443;
      111944:data<=-16'd4316;
      111945:data<=-16'd3700;
      111946:data<=-16'd3647;
      111947:data<=-16'd2890;
      111948:data<=-16'd2904;
      111949:data<=-16'd4716;
      111950:data<=-16'd4945;
      111951:data<=-16'd4190;
      111952:data<=-16'd4152;
      111953:data<=-16'd3701;
      111954:data<=-16'd3413;
      111955:data<=-16'd3234;
      111956:data<=-16'd2722;
      111957:data<=-16'd2422;
      111958:data<=-16'd2055;
      111959:data<=-16'd1967;
      111960:data<=-16'd1668;
      111961:data<=-16'd1204;
      111962:data<=-16'd2158;
      111963:data<=-16'd3178;
      111964:data<=-16'd3300;
      111965:data<=-16'd2996;
      111966:data<=-16'd1942;
      111967:data<=-16'd1612;
      111968:data<=-16'd1765;
      111969:data<=-16'd1216;
      111970:data<=-16'd1031;
      111971:data<=-16'd619;
      111972:data<=-16'd281;
      111973:data<=-16'd246;
      111974:data<=16'd505;
      111975:data<=-16'd456;
      111976:data<=-16'd1149;
      111977:data<=16'd1618;
      111978:data<=16'd2919;
      111979:data<=16'd2514;
      111980:data<=16'd3392;
      111981:data<=16'd3104;
      111982:data<=16'd2729;
      111983:data<=16'd3468;
      111984:data<=16'd3336;
      111985:data<=16'd3407;
      111986:data<=16'd3788;
      111987:data<=16'd3724;
      111988:data<=16'd3278;
      111989:data<=16'd1850;
      111990:data<=16'd1268;
      111991:data<=16'd1824;
      111992:data<=16'd1715;
      111993:data<=16'd1807;
      111994:data<=16'd1882;
      111995:data<=16'd1615;
      111996:data<=16'd2067;
      111997:data<=16'd2375;
      111998:data<=16'd2385;
      111999:data<=16'd2572;
      112000:data<=16'd2590;
      112001:data<=16'd2238;
      112002:data<=16'd992;
      112003:data<=16'd253;
      112004:data<=16'd757;
      112005:data<=16'd657;
      112006:data<=16'd560;
      112007:data<=16'd983;
      112008:data<=16'd1075;
      112009:data<=16'd1381;
      112010:data<=16'd1412;
      112011:data<=16'd1284;
      112012:data<=16'd1545;
      112013:data<=16'd1450;
      112014:data<=16'd1579;
      112015:data<=16'd1002;
      112016:data<=-16'd526;
      112017:data<=-16'd367;
      112018:data<=16'd135;
      112019:data<=-16'd55;
      112020:data<=16'd438;
      112021:data<=16'd252;
      112022:data<=16'd171;
      112023:data<=16'd858;
      112024:data<=16'd637;
      112025:data<=16'd878;
      112026:data<=16'd1051;
      112027:data<=16'd731;
      112028:data<=16'd1915;
      112029:data<=16'd1107;
      112030:data<=-16'd2221;
      112031:data<=-16'd2996;
      112032:data<=-16'd2272;
      112033:data<=-16'd2121;
      112034:data<=-16'd1921;
      112035:data<=-16'd2088;
      112036:data<=-16'd1867;
      112037:data<=-16'd1448;
      112038:data<=-16'd1284;
      112039:data<=-16'd655;
      112040:data<=-16'd660;
      112041:data<=-16'd376;
      112042:data<=16'd1262;
      112043:data<=16'd1886;
      112044:data<=16'd1807;
      112045:data<=16'd1980;
      112046:data<=16'd1744;
      112047:data<=16'd2038;
      112048:data<=16'd2190;
      112049:data<=16'd1703;
      112050:data<=16'd2065;
      112051:data<=16'd2441;
      112052:data<=16'd2414;
      112053:data<=16'd2623;
      112054:data<=16'd2775;
      112055:data<=16'd3721;
      112056:data<=16'd4845;
      112057:data<=16'd4793;
      112058:data<=16'd4757;
      112059:data<=16'd4737;
      112060:data<=16'd4240;
      112061:data<=16'd4225;
      112062:data<=16'd4473;
      112063:data<=16'd4478;
      112064:data<=16'd4244;
      112065:data<=16'd4076;
      112066:data<=16'd4294;
      112067:data<=16'd4223;
      112068:data<=16'd4696;
      112069:data<=16'd6087;
      112070:data<=16'd6119;
      112071:data<=16'd5647;
      112072:data<=16'd6131;
      112073:data<=16'd5792;
      112074:data<=16'd5283;
      112075:data<=16'd5698;
      112076:data<=16'd5735;
      112077:data<=16'd5426;
      112078:data<=16'd5086;
      112079:data<=16'd4919;
      112080:data<=16'd5089;
      112081:data<=16'd5266;
      112082:data<=16'd7248;
      112083:data<=16'd10320;
      112084:data<=16'd10818;
      112085:data<=16'd10357;
      112086:data<=16'd10740;
      112087:data<=16'd10194;
      112088:data<=16'd9711;
      112089:data<=16'd9811;
      112090:data<=16'd9320;
      112091:data<=16'd9098;
      112092:data<=16'd8728;
      112093:data<=16'd7856;
      112094:data<=16'd8279;
      112095:data<=16'd9518;
      112096:data<=16'd9799;
      112097:data<=16'd9236;
      112098:data<=16'd8828;
      112099:data<=16'd8715;
      112100:data<=16'd8169;
      112101:data<=16'd7697;
      112102:data<=16'd7677;
      112103:data<=16'd7150;
      112104:data<=16'd6816;
      112105:data<=16'd7057;
      112106:data<=16'd6543;
      112107:data<=16'd6078;
      112108:data<=16'd6781;
      112109:data<=16'd7582;
      112110:data<=16'd7642;
      112111:data<=16'd7095;
      112112:data<=16'd6388;
      112113:data<=16'd5927;
      112114:data<=16'd5799;
      112115:data<=16'd5794;
      112116:data<=16'd5404;
      112117:data<=16'd4937;
      112118:data<=16'd4945;
      112119:data<=16'd4834;
      112120:data<=16'd4482;
      112121:data<=16'd4696;
      112122:data<=16'd5653;
      112123:data<=16'd6366;
      112124:data<=16'd5952;
      112125:data<=16'd5289;
      112126:data<=16'd4887;
      112127:data<=16'd4256;
      112128:data<=16'd4203;
      112129:data<=16'd4385;
      112130:data<=16'd3824;
      112131:data<=16'd3632;
      112132:data<=16'd3210;
      112133:data<=16'd2331;
      112134:data<=16'd3550;
      112135:data<=16'd4842;
      112136:data<=16'd2769;
      112137:data<=16'd300;
      112138:data<=16'd15;
      112139:data<=16'd92;
      112140:data<=-16'd265;
      112141:data<=-16'd412;
      112142:data<=-16'd444;
      112143:data<=-16'd619;
      112144:data<=-16'd860;
      112145:data<=-16'd1145;
      112146:data<=-16'd1265;
      112147:data<=-16'd464;
      112148:data<=16'd1022;
      112149:data<=16'd1548;
      112150:data<=16'd870;
      112151:data<=16'd405;
      112152:data<=16'd519;
      112153:data<=16'd564;
      112154:data<=16'd434;
      112155:data<=16'd243;
      112156:data<=16'd85;
      112157:data<=16'd176;
      112158:data<=16'd135;
      112159:data<=-16'd325;
      112160:data<=-16'd218;
      112161:data<=16'd831;
      112162:data<=16'd1657;
      112163:data<=16'd1806;
      112164:data<=16'd1765;
      112165:data<=16'd1579;
      112166:data<=16'd1259;
      112167:data<=16'd954;
      112168:data<=16'd522;
      112169:data<=16'd165;
      112170:data<=16'd358;
      112171:data<=16'd719;
      112172:data<=16'd452;
      112173:data<=-16'd56;
      112174:data<=16'd429;
      112175:data<=16'd1715;
      112176:data<=16'd2229;
      112177:data<=16'd1864;
      112178:data<=16'd1626;
      112179:data<=16'd1375;
      112180:data<=16'd1101;
      112181:data<=16'd1122;
      112182:data<=16'd925;
      112183:data<=16'd749;
      112184:data<=16'd843;
      112185:data<=16'd564;
      112186:data<=16'd438;
      112187:data<=16'd796;
      112188:data<=16'd1748;
      112189:data<=16'd4290;
      112190:data<=16'd6479;
      112191:data<=16'd6111;
      112192:data<=16'd5336;
      112193:data<=16'd5247;
      112194:data<=16'd4962;
      112195:data<=16'd4942;
      112196:data<=16'd4731;
      112197:data<=16'd4087;
      112198:data<=16'd3800;
      112199:data<=16'd3424;
      112200:data<=16'd3471;
      112201:data<=16'd4499;
      112202:data<=16'd4957;
      112203:data<=16'd4511;
      112204:data<=16'd3930;
      112205:data<=16'd3479;
      112206:data<=16'd3368;
      112207:data<=16'd3027;
      112208:data<=16'd2535;
      112209:data<=16'd2420;
      112210:data<=16'd2006;
      112211:data<=16'd1607;
      112212:data<=16'd1460;
      112213:data<=16'd1021;
      112214:data<=16'd1601;
      112215:data<=16'd3027;
      112216:data<=16'd3037;
      112217:data<=16'd2027;
      112218:data<=16'd1460;
      112219:data<=16'd1497;
      112220:data<=16'd1624;
      112221:data<=16'd1221;
      112222:data<=16'd714;
      112223:data<=16'd491;
      112224:data<=16'd440;
      112225:data<=16'd470;
      112226:data<=-16'd12;
      112227:data<=16'd38;
      112228:data<=16'd1350;
      112229:data<=16'd1818;
      112230:data<=16'd1354;
      112231:data<=16'd1017;
      112232:data<=16'd432;
      112233:data<=16'd347;
      112234:data<=16'd426;
      112235:data<=-16'd176;
      112236:data<=-16'd614;
      112237:data<=-16'd937;
      112238:data<=-16'd939;
      112239:data<=-16'd983;
      112240:data<=-16'd1500;
      112241:data<=-16'd1005;
      112242:data<=-16'd2140;
      112243:data<=-16'd5841;
      112244:data<=-16'd6604;
      112245:data<=-16'd5814;
      112246:data<=-16'd6639;
      112247:data<=-16'd6287;
      112248:data<=-16'd5999;
      112249:data<=-16'd6592;
      112250:data<=-16'd6159;
      112251:data<=-16'd6347;
      112252:data<=-16'd6534;
      112253:data<=-16'd6269;
      112254:data<=-16'd7294;
      112255:data<=-16'd7821;
      112256:data<=-16'd7741;
      112257:data<=-16'd7946;
      112258:data<=-16'd7606;
      112259:data<=-16'd7777;
      112260:data<=-16'd7703;
      112261:data<=-16'd7233;
      112262:data<=-16'd7711;
      112263:data<=-16'd7141;
      112264:data<=-16'd6583;
      112265:data<=-16'd7233;
      112266:data<=-16'd6683;
      112267:data<=-16'd7007;
      112268:data<=-16'd8499;
      112269:data<=-16'd8238;
      112270:data<=-16'd8000;
      112271:data<=-16'd8116;
      112272:data<=-16'd7561;
      112273:data<=-16'd7423;
      112274:data<=-16'd7357;
      112275:data<=-16'd7468;
      112276:data<=-16'd7491;
      112277:data<=-16'd6983;
      112278:data<=-16'd6909;
      112279:data<=-16'd6561;
      112280:data<=-16'd6927;
      112281:data<=-16'd8516;
      112282:data<=-16'd8420;
      112283:data<=-16'd7952;
      112284:data<=-16'd8216;
      112285:data<=-16'd7370;
      112286:data<=-16'd6954;
      112287:data<=-16'd7083;
      112288:data<=-16'd6751;
      112289:data<=-16'd6710;
      112290:data<=-16'd6357;
      112291:data<=-16'd6064;
      112292:data<=-16'd5583;
      112293:data<=-16'd5357;
      112294:data<=-16'd7333;
      112295:data<=-16'd6946;
      112296:data<=-16'd3004;
      112297:data<=-16'd1944;
      112298:data<=-16'd2689;
      112299:data<=-16'd2356;
      112300:data<=-16'd2491;
      112301:data<=-16'd2240;
      112302:data<=-16'd1968;
      112303:data<=-16'd2441;
      112304:data<=-16'd2335;
      112305:data<=-16'd1941;
      112306:data<=-16'd1748;
      112307:data<=-16'd2604;
      112308:data<=-16'd3993;
      112309:data<=-16'd3741;
      112310:data<=-16'd3289;
      112311:data<=-16'd3407;
      112312:data<=-16'd3124;
      112313:data<=-16'd3386;
      112314:data<=-16'd3266;
      112315:data<=-16'd2575;
      112316:data<=-16'd2773;
      112317:data<=-16'd2845;
      112318:data<=-16'd2547;
      112319:data<=-16'd2329;
      112320:data<=-16'd2572;
      112321:data<=-16'd3859;
      112322:data<=-16'd4267;
      112323:data<=-16'd3841;
      112324:data<=-16'd4020;
      112325:data<=-16'd3504;
      112326:data<=-16'd3127;
      112327:data<=-16'd3529;
      112328:data<=-16'd3174;
      112329:data<=-16'd2833;
      112330:data<=-16'd2726;
      112331:data<=-16'd2487;
      112332:data<=-16'd2619;
      112333:data<=-16'd2849;
      112334:data<=-16'd3735;
      112335:data<=-16'd4411;
      112336:data<=-16'd3808;
      112337:data<=-16'd3751;
      112338:data<=-16'd3811;
      112339:data<=-16'd3256;
      112340:data<=-16'd3184;
      112341:data<=-16'd2719;
      112342:data<=-16'd2523;
      112343:data<=-16'd3159;
      112344:data<=-16'd2628;
      112345:data<=-16'd2143;
      112346:data<=-16'd2833;
      112347:data<=-16'd3553;
      112348:data<=-16'd5357;
      112349:data<=-16'd7759;
      112350:data<=-16'd8345;
      112351:data<=-16'd7821;
      112352:data<=-16'd7645;
      112353:data<=-16'd7313;
      112354:data<=-16'd6610;
      112355:data<=-16'd6370;
      112356:data<=-16'd6473;
      112357:data<=-16'd6100;
      112358:data<=-16'd5424;
      112359:data<=-16'd5089;
      112360:data<=-16'd5739;
      112361:data<=-16'd6805;
      112362:data<=-16'd6604;
      112363:data<=-16'd5708;
      112364:data<=-16'd5403;
      112365:data<=-16'd5090;
      112366:data<=-16'd4678;
      112367:data<=-16'd4422;
      112368:data<=-16'd3897;
      112369:data<=-16'd3347;
      112370:data<=-16'd3388;
      112371:data<=-16'd3529;
      112372:data<=-16'd2989;
      112373:data<=-16'd3031;
      112374:data<=-16'd4337;
      112375:data<=-16'd4746;
      112376:data<=-16'd4068;
      112377:data<=-16'd3586;
      112378:data<=-16'd2893;
      112379:data<=-16'd2561;
      112380:data<=-16'd2826;
      112381:data<=-16'd2411;
      112382:data<=-16'd1712;
      112383:data<=-16'd1657;
      112384:data<=-16'd1735;
      112385:data<=-16'd1409;
      112386:data<=-16'd1613;
      112387:data<=-16'd2784;
      112388:data<=-16'd3146;
      112389:data<=-16'd2673;
      112390:data<=-16'd2572;
      112391:data<=-16'd2053;
      112392:data<=-16'd1424;
      112393:data<=-16'd1383;
      112394:data<=-16'd1336;
      112395:data<=-16'd1207;
      112396:data<=-16'd778;
      112397:data<=-16'd475;
      112398:data<=-16'd270;
      112399:data<=-16'd83;
      112400:data<=-16'd1541;
      112401:data<=-16'd1659;
      112402:data<=16'd1774;
      112403:data<=16'd3421;
      112404:data<=16'd2930;
      112405:data<=16'd3342;
      112406:data<=16'd3200;
      112407:data<=16'd3306;
      112408:data<=16'd3927;
      112409:data<=16'd3510;
      112410:data<=16'd3428;
      112411:data<=16'd3709;
      112412:data<=16'd3845;
      112413:data<=16'd3345;
      112414:data<=16'd1471;
      112415:data<=16'd996;
      112416:data<=16'd1903;
      112417:data<=16'd1858;
      112418:data<=16'd2137;
      112419:data<=16'd2308;
      112420:data<=16'd2033;
      112421:data<=16'd2400;
      112422:data<=16'd2167;
      112423:data<=16'd1855;
      112424:data<=16'd2226;
      112425:data<=16'd2461;
      112426:data<=16'd2299;
      112427:data<=16'd854;
      112428:data<=-16'd33;
      112429:data<=16'd776;
      112430:data<=16'd717;
      112431:data<=16'd807;
      112432:data<=16'd1412;
      112433:data<=16'd905;
      112434:data<=16'd1057;
      112435:data<=16'd1497;
      112436:data<=16'd1310;
      112437:data<=16'd1633;
      112438:data<=16'd1682;
      112439:data<=16'd1416;
      112440:data<=16'd717;
      112441:data<=-16'd185;
      112442:data<=16'd294;
      112443:data<=16'd382;
      112444:data<=16'd77;
      112445:data<=16'd754;
      112446:data<=16'd350;
      112447:data<=16'd162;
      112448:data<=16'd1042;
      112449:data<=16'd866;
      112450:data<=16'd933;
      112451:data<=16'd1045;
      112452:data<=16'd746;
      112453:data<=16'd1491;
      112454:data<=16'd1004;
      112455:data<=-16'd1189;
      112456:data<=-16'd2628;
      112457:data<=-16'd2928;
      112458:data<=-16'd2329;
      112459:data<=-16'd2015;
      112460:data<=-16'd1847;
      112461:data<=-16'd1257;
      112462:data<=-16'd1588;
      112463:data<=-16'd1348;
      112464:data<=-16'd487;
      112465:data<=-16'd926;
      112466:data<=-16'd300;
      112467:data<=16'd1324;
      112468:data<=16'd1744;
      112469:data<=16'd2000;
      112470:data<=16'd2103;
      112471:data<=16'd1985;
      112472:data<=16'd2073;
      112473:data<=16'd2187;
      112474:data<=16'd2760;
      112475:data<=16'd2798;
      112476:data<=16'd2544;
      112477:data<=16'd2875;
      112478:data<=16'd2604;
      112479:data<=16'd3228;
      112480:data<=16'd4927;
      112481:data<=16'd5060;
      112482:data<=16'd4792;
      112483:data<=16'd4971;
      112484:data<=16'd4954;
      112485:data<=16'd5009;
      112486:data<=16'd4623;
      112487:data<=16'd4551;
      112488:data<=16'd4795;
      112489:data<=16'd4444;
      112490:data<=16'd4372;
      112491:data<=16'd4103;
      112492:data<=16'd4408;
      112493:data<=16'd6128;
      112494:data<=16'd6467;
      112495:data<=16'd5858;
      112496:data<=16'd5958;
      112497:data<=16'd5883;
      112498:data<=16'd6079;
      112499:data<=16'd5946;
      112500:data<=16'd5213;
      112501:data<=16'd5140;
      112502:data<=16'd5213;
      112503:data<=16'd5468;
      112504:data<=16'd5429;
      112505:data<=16'd4966;
      112506:data<=16'd5717;
      112507:data<=16'd6781;
      112508:data<=16'd8511;
      112509:data<=16'd10991;
      112510:data<=16'd11006;
      112511:data<=16'd10240;
      112512:data<=16'd10263;
      112513:data<=16'd9298;
      112514:data<=16'd8945;
      112515:data<=16'd8989;
      112516:data<=16'd8619;
      112517:data<=16'd8765;
      112518:data<=16'd7962;
      112519:data<=16'd7921;
      112520:data<=16'd9582;
      112521:data<=16'd9588;
      112522:data<=16'd9036;
      112523:data<=16'd8919;
      112524:data<=16'd8108;
      112525:data<=16'd7706;
      112526:data<=16'd7342;
      112527:data<=16'd6972;
      112528:data<=16'd6828;
      112529:data<=16'd6179;
      112530:data<=16'd6056;
      112531:data<=16'd5755;
      112532:data<=16'd5680;
      112533:data<=16'd7338;
      112534:data<=16'd7629;
      112535:data<=16'd6799;
      112536:data<=16'd7062;
      112537:data<=16'd6394;
      112538:data<=16'd5568;
      112539:data<=16'd5495;
      112540:data<=16'd5087;
      112541:data<=16'd5109;
      112542:data<=16'd4869;
      112543:data<=16'd4364;
      112544:data<=16'd4337;
      112545:data<=16'd4244;
      112546:data<=16'd5328;
      112547:data<=16'd6287;
      112548:data<=16'd5547;
      112549:data<=16'd5345;
      112550:data<=16'd5093;
      112551:data<=16'd4428;
      112552:data<=16'd4400;
      112553:data<=16'd3656;
      112554:data<=16'd3192;
      112555:data<=16'd3457;
      112556:data<=16'd3171;
      112557:data<=16'd3074;
      112558:data<=16'd2438;
      112559:data<=16'd2836;
      112560:data<=16'd5313;
      112561:data<=16'd4097;
      112562:data<=-16'd3;
      112563:data<=-16'd852;
      112564:data<=-16'd356;
      112565:data<=-16'd751;
      112566:data<=-16'd879;
      112567:data<=-16'd1324;
      112568:data<=-16'd1674;
      112569:data<=-16'd1242;
      112570:data<=-16'd1155;
      112571:data<=-16'd1515;
      112572:data<=-16'd890;
      112573:data<=16'd652;
      112574:data<=16'd1242;
      112575:data<=16'd845;
      112576:data<=16'd616;
      112577:data<=16'd258;
      112578:data<=-16'd82;
      112579:data<=16'd8;
      112580:data<=-16'd121;
      112581:data<=-16'd476;
      112582:data<=-16'd511;
      112583:data<=-16'd516;
      112584:data<=-16'd726;
      112585:data<=-16'd115;
      112586:data<=16'd1201;
      112587:data<=16'd1389;
      112588:data<=16'd952;
      112589:data<=16'd1034;
      112590:data<=16'd816;
      112591:data<=16'd466;
      112592:data<=16'd334;
      112593:data<=16'd89;
      112594:data<=16'd8;
      112595:data<=-16'd124;
      112596:data<=-16'd347;
      112597:data<=-16'd534;
      112598:data<=-16'd399;
      112599:data<=16'd864;
      112600:data<=16'd1756;
      112601:data<=16'd1212;
      112602:data<=16'd920;
      112603:data<=16'd919;
      112604:data<=16'd749;
      112605:data<=16'd701;
      112606:data<=16'd193;
      112607:data<=-16'd220;
      112608:data<=-16'd18;
      112609:data<=-16'd21;
      112610:data<=-16'd467;
      112611:data<=-16'd546;
      112612:data<=16'd381;
      112613:data<=16'd1221;
      112614:data<=16'd2317;
      112615:data<=16'd4805;
      112616:data<=16'd5774;
      112617:data<=16'd4874;
      112618:data<=16'd4814;
      112619:data<=16'd4414;
      112620:data<=16'd3762;
      112621:data<=16'd3845;
      112622:data<=16'd3579;
      112623:data<=16'd3571;
      112624:data<=16'd3228;
      112625:data<=16'd2801;
      112626:data<=16'd4076;
      112627:data<=16'd4460;
      112628:data<=16'd3626;
      112629:data<=16'd3559;
      112630:data<=16'd2917;
      112631:data<=16'd2473;
      112632:data<=16'd2472;
      112633:data<=16'd1676;
      112634:data<=16'd1516;
      112635:data<=16'd1418;
      112636:data<=16'd946;
      112637:data<=16'd986;
      112638:data<=16'd725;
      112639:data<=16'd1359;
      112640:data<=16'd2432;
      112641:data<=16'd2093;
      112642:data<=16'd2068;
      112643:data<=16'd1882;
      112644:data<=16'd869;
      112645:data<=16'd708;
      112646:data<=16'd658;
      112647:data<=16'd614;
      112648:data<=16'd567;
      112649:data<=-16'd124;
      112650:data<=-16'd271;
      112651:data<=-16'd249;
      112652:data<=16'd253;
      112653:data<=16'd1412;
      112654:data<=16'd1043;
      112655:data<=16'd766;
      112656:data<=16'd1064;
      112657:data<=-16'd96;
      112658:data<=-16'd538;
      112659:data<=-16'd109;
      112660:data<=-16'd247;
      112661:data<=-16'd256;
      112662:data<=-16'd814;
      112663:data<=-16'd1201;
      112664:data<=-16'd1409;
      112665:data<=-16'd1970;
      112666:data<=-16'd1058;
      112667:data<=-16'd1844;
      112668:data<=-16'd5548;
      112669:data<=-16'd6834;
      112670:data<=-16'd6294;
      112671:data<=-16'd6200;
      112672:data<=-16'd6014;
      112673:data<=-16'd6680;
      112674:data<=-16'd6871;
      112675:data<=-16'd6335;
      112676:data<=-16'd6420;
      112677:data<=-16'd6037;
      112678:data<=-16'd6434;
      112679:data<=-16'd7827;
      112680:data<=-16'd7982;
      112681:data<=-16'd7817;
      112682:data<=-16'd7712;
      112683:data<=-16'd7418;
      112684:data<=-16'd7397;
      112685:data<=-16'd6980;
      112686:data<=-16'd6963;
      112687:data<=-16'd7279;
      112688:data<=-16'd6889;
      112689:data<=-16'd6702;
      112690:data<=-16'd6354;
      112691:data<=-16'd6310;
      112692:data<=-16'd7694;
      112693:data<=-16'd8505;
      112694:data<=-16'd8160;
      112695:data<=-16'd7720;
      112696:data<=-16'd7483;
      112697:data<=-16'd7696;
      112698:data<=-16'd7468;
      112699:data<=-16'd7054;
      112700:data<=-16'd7065;
      112701:data<=-16'd6725;
      112702:data<=-16'd6775;
      112703:data<=-16'd6798;
      112704:data<=-16'd6205;
      112705:data<=-16'd6983;
      112706:data<=-16'd8197;
      112707:data<=-16'd8070;
      112708:data<=-16'd7553;
      112709:data<=-16'd7043;
      112710:data<=-16'd6843;
      112711:data<=-16'd6673;
      112712:data<=-16'd6175;
      112713:data<=-16'd6159;
      112714:data<=-16'd5832;
      112715:data<=-16'd5448;
      112716:data<=-16'd5911;
      112717:data<=-16'd5404;
      112718:data<=-16'd5204;
      112719:data<=-16'd6940;
      112720:data<=-16'd6581;
      112721:data<=-16'd3365;
      112722:data<=-16'd1709;
      112723:data<=-16'd1900;
      112724:data<=-16'd1592;
      112725:data<=-16'd1439;
      112726:data<=-16'd1786;
      112727:data<=-16'd1368;
      112728:data<=-16'd1145;
      112729:data<=-16'd1574;
      112730:data<=-16'd1415;
      112731:data<=-16'd1879;
      112732:data<=-16'd3174;
      112733:data<=-16'd3359;
      112734:data<=-16'd3086;
      112735:data<=-16'd3133;
      112736:data<=-16'd2924;
      112737:data<=-16'd2608;
      112738:data<=-16'd2367;
      112739:data<=-16'd2387;
      112740:data<=-16'd2328;
      112741:data<=-16'd2047;
      112742:data<=-16'd2126;
      112743:data<=-16'd1924;
      112744:data<=-16'd1965;
      112745:data<=-16'd3245;
      112746:data<=-16'd3950;
      112747:data<=-16'd3544;
      112748:data<=-16'd3283;
      112749:data<=-16'd3193;
      112750:data<=-16'd3024;
      112751:data<=-16'd2555;
      112752:data<=-16'd2335;
      112753:data<=-16'd2569;
      112754:data<=-16'd2329;
      112755:data<=-16'd2212;
      112756:data<=-16'd2168;
      112757:data<=-16'd1623;
      112758:data<=-16'd2226;
      112759:data<=-16'd3607;
      112760:data<=-16'd3747;
      112761:data<=-16'd3122;
      112762:data<=-16'd2822;
      112763:data<=-16'd2889;
      112764:data<=-16'd2786;
      112765:data<=-16'd2689;
      112766:data<=-16'd2649;
      112767:data<=-16'd2073;
      112768:data<=-16'd2140;
      112769:data<=-16'd2504;
      112770:data<=-16'd1856;
      112771:data<=-16'd2460;
      112772:data<=-16'd3829;
      112773:data<=-16'd4314;
      112774:data<=-16'd6140;
      112775:data<=-16'd7715;
      112776:data<=-16'd7045;
      112777:data<=-16'd6875;
      112778:data<=-16'd7131;
      112779:data<=-16'd6495;
      112780:data<=-16'd5799;
      112781:data<=-16'd5397;
      112782:data<=-16'd5266;
      112783:data<=-16'd4839;
      112784:data<=-16'd4910;
      112785:data<=-16'd6120;
      112786:data<=-16'd6325;
      112787:data<=-16'd5765;
      112788:data<=-16'd5510;
      112789:data<=-16'd4777;
      112790:data<=-16'd4534;
      112791:data<=-16'd4575;
      112792:data<=-16'd3958;
      112793:data<=-16'd3667;
      112794:data<=-16'd3359;
      112795:data<=-16'd3025;
      112796:data<=-16'd2945;
      112797:data<=-16'd2699;
      112798:data<=-16'd3554;
      112799:data<=-16'd4549;
      112800:data<=-16'd3923;
      112801:data<=-16'd3415;
      112802:data<=-16'd3375;
      112803:data<=-16'd3069;
      112804:data<=-16'd2845;
      112805:data<=-16'd2366;
      112806:data<=-16'd1991;
      112807:data<=-16'd1868;
      112808:data<=-16'd1662;
      112809:data<=-16'd1430;
      112810:data<=-16'd758;
      112811:data<=-16'd1149;
      112812:data<=-16'd2957;
      112813:data<=-16'd3203;
      112814:data<=-16'd2258;
      112815:data<=-16'd1941;
      112816:data<=-16'd1729;
      112817:data<=-16'd1712;
      112818:data<=-16'd1463;
      112819:data<=-16'd761;
      112820:data<=-16'd702;
      112821:data<=-16'd813;
      112822:data<=-16'd472;
      112823:data<=16'd83;
      112824:data<=16'd79;
      112825:data<=-16'd1465;
      112826:data<=-16'd2231;
      112827:data<=16'd227;
      112828:data<=16'd3186;
      112829:data<=16'd3882;
      112830:data<=16'd3598;
      112831:data<=16'd3792;
      112832:data<=16'd3911;
      112833:data<=16'd3824;
      112834:data<=16'd4159;
      112835:data<=16'd4353;
      112836:data<=16'd4158;
      112837:data<=16'd3798;
      112838:data<=16'd2635;
      112839:data<=16'd1626;
      112840:data<=16'd1897;
      112841:data<=16'd2181;
      112842:data<=16'd2127;
      112843:data<=16'd2362;
      112844:data<=16'd2399;
      112845:data<=16'd2223;
      112846:data<=16'd2359;
      112847:data<=16'd2673;
      112848:data<=16'd2781;
      112849:data<=16'd2796;
      112850:data<=16'd2748;
      112851:data<=16'd1959;
      112852:data<=16'd878;
      112853:data<=16'd839;
      112854:data<=16'd1401;
      112855:data<=16'd1406;
      112856:data<=16'd1169;
      112857:data<=16'd1503;
      112858:data<=16'd1936;
      112859:data<=16'd1835;
      112860:data<=16'd1798;
      112861:data<=16'd1880;
      112862:data<=16'd1979;
      112863:data<=16'd2308;
      112864:data<=16'd1527;
      112865:data<=16'd73;
      112866:data<=16'd183;
      112867:data<=16'd781;
      112868:data<=16'd591;
      112869:data<=16'd441;
      112870:data<=16'd376;
      112871:data<=16'd484;
      112872:data<=16'd904;
      112873:data<=16'd1312;
      112874:data<=16'd1424;
      112875:data<=16'd1192;
      112876:data<=16'd1524;
      112877:data<=16'd1804;
      112878:data<=16'd1395;
      112879:data<=16'd1791;
      112880:data<=16'd940;
      112881:data<=-16'd1955;
      112882:data<=-16'd2455;
      112883:data<=-16'd1686;
      112884:data<=-16'd2296;
      112885:data<=-16'd1902;
      112886:data<=-16'd1324;
      112887:data<=-16'd1629;
      112888:data<=-16'd1122;
      112889:data<=-16'd748;
      112890:data<=-16'd314;
      112891:data<=16'd1163;
      112892:data<=16'd1971;
      112893:data<=16'd1911;
      112894:data<=16'd1918;
      112895:data<=16'd2217;
      112896:data<=16'd2722;
      112897:data<=16'd2640;
      112898:data<=16'd2494;
      112899:data<=16'd2795;
      112900:data<=16'd2861;
      112901:data<=16'd3093;
      112902:data<=16'd3051;
      112903:data<=16'd2547;
      112904:data<=16'd3512;
      112905:data<=16'd5321;
      112906:data<=16'd5717;
      112907:data<=16'd5174;
      112908:data<=16'd5037;
      112909:data<=16'd5300;
      112910:data<=16'd5257;
      112911:data<=16'd4983;
      112912:data<=16'd4942;
      112913:data<=16'd4968;
      112914:data<=16'd5095;
      112915:data<=16'd5049;
      112916:data<=16'd4708;
      112917:data<=16'd5285;
      112918:data<=16'd6586;
      112919:data<=16'd7086;
      112920:data<=16'd6777;
      112921:data<=16'd6495;
      112922:data<=16'd6487;
      112923:data<=16'd6308;
      112924:data<=16'd6164;
      112925:data<=16'd6311;
      112926:data<=16'd5824;
      112927:data<=16'd5597;
      112928:data<=16'd6103;
      112929:data<=16'd5510;
      112930:data<=16'd5607;
      112931:data<=16'd7178;
      112932:data<=16'd7166;
      112933:data<=16'd7975;
      112934:data<=16'd10957;
      112935:data<=16'd11402;
      112936:data<=16'd10346;
      112937:data<=16'd10645;
      112938:data<=16'd10260;
      112939:data<=16'd9608;
      112940:data<=16'd9729;
      112941:data<=16'd9317;
      112942:data<=16'd8693;
      112943:data<=16'd8548;
      112944:data<=16'd9230;
      112945:data<=16'd10223;
      112946:data<=16'd9737;
      112947:data<=16'd8715;
      112948:data<=16'd8608;
      112949:data<=16'd8290;
      112950:data<=16'd7721;
      112951:data<=16'd7544;
      112952:data<=16'd7341;
      112953:data<=16'd7169;
      112954:data<=16'd7101;
      112955:data<=16'd6658;
      112956:data<=16'd5949;
      112957:data<=16'd6460;
      112958:data<=16'd8031;
      112959:data<=16'd7761;
      112960:data<=16'd6385;
      112961:data<=16'd6584;
      112962:data<=16'd6619;
      112963:data<=16'd5850;
      112964:data<=16'd5862;
      112965:data<=16'd5547;
      112966:data<=16'd4866;
      112967:data<=16'd4995;
      112968:data<=16'd4939;
      112969:data<=16'd4490;
      112970:data<=16'd4749;
      112971:data<=16'd5720;
      112972:data<=16'd6141;
      112973:data<=16'd5459;
      112974:data<=16'd5018;
      112975:data<=16'd4916;
      112976:data<=16'd4273;
      112977:data<=16'd3952;
      112978:data<=16'd4008;
      112979:data<=16'd3785;
      112980:data<=16'd3482;
      112981:data<=16'd3068;
      112982:data<=16'd3022;
      112983:data<=16'd3388;
      112984:data<=16'd3990;
      112985:data<=16'd4925;
      112986:data<=16'd3750;
      112987:data<=16'd458;
      112988:data<=-16'd819;
      112989:data<=-16'd497;
      112990:data<=-16'd751;
      112991:data<=-16'd714;
      112992:data<=-16'd822;
      112993:data<=-16'd1315;
      112994:data<=-16'd1366;
      112995:data<=-16'd1447;
      112996:data<=-16'd1095;
      112997:data<=16'd29;
      112998:data<=16'd758;
      112999:data<=16'd643;
      113000:data<=16'd50;
      113001:data<=-16'd179;
      113002:data<=16'd61;
      113003:data<=-16'd92;
      113004:data<=-16'd405;
      113005:data<=-16'd660;
      113006:data<=-16'd949;
      113007:data<=-16'd970;
      113008:data<=-16'd1240;
      113009:data<=-16'd1401;
      113010:data<=-16'd423;
      113011:data<=16'd701;
      113012:data<=16'd905;
      113013:data<=16'd506;
      113014:data<=16'd220;
      113015:data<=16'd340;
      113016:data<=16'd258;
      113017:data<=-16'd126;
      113018:data<=-16'd500;
      113019:data<=-16'd793;
      113020:data<=-16'd484;
      113021:data<=-16'd409;
      113022:data<=-16'd1140;
      113023:data<=-16'd667;
      113024:data<=16'd817;
      113025:data<=16'd1152;
      113026:data<=16'd802;
      113027:data<=16'd488;
      113028:data<=16'd0;
      113029:data<=-16'd58;
      113030:data<=16'd241;
      113031:data<=-16'd153;
      113032:data<=-16'd996;
      113033:data<=-16'd916;
      113034:data<=-16'd496;
      113035:data<=-16'd1057;
      113036:data<=-16'd922;
      113037:data<=16'd256;
      113038:data<=16'd367;
      113039:data<=16'd1239;
      113040:data<=16'd3735;
      113041:data<=16'd4214;
      113042:data<=16'd3292;
      113043:data<=16'd3541;
      113044:data<=16'd3600;
      113045:data<=16'd3049;
      113046:data<=16'd2594;
      113047:data<=16'd2117;
      113048:data<=16'd1982;
      113049:data<=16'd1773;
      113050:data<=16'd1939;
      113051:data<=16'd3140;
      113052:data<=16'd3316;
      113053:data<=16'd2538;
      113054:data<=16'd2538;
      113055:data<=16'd2146;
      113056:data<=16'd1350;
      113057:data<=16'd1271;
      113058:data<=16'd1039;
      113059:data<=16'd711;
      113060:data<=16'd789;
      113061:data<=16'd496;
      113062:data<=-16'd86;
      113063:data<=16'd284;
      113064:data<=16'd1717;
      113065:data<=16'd2161;
      113066:data<=16'd1063;
      113067:data<=16'd544;
      113068:data<=16'd682;
      113069:data<=16'd431;
      113070:data<=16'd253;
      113071:data<=-16'd20;
      113072:data<=-16'd467;
      113073:data<=-16'd599;
      113074:data<=-16'd810;
      113075:data<=-16'd1234;
      113076:data<=-16'd1083;
      113077:data<=16'd140;
      113078:data<=16'd1013;
      113079:data<=16'd375;
      113080:data<=-16'd103;
      113081:data<=-16'd105;
      113082:data<=-16'd564;
      113083:data<=-16'd579;
      113084:data<=-16'd593;
      113085:data<=-16'd964;
      113086:data<=-16'd866;
      113087:data<=-16'd1146;
      113088:data<=-16'd1416;
      113089:data<=-16'd1366;
      113090:data<=-16'd1902;
      113091:data<=-16'd1779;
      113092:data<=-16'd2212;
      113093:data<=-16'd4833;
      113094:data<=-16'd6405;
      113095:data<=-16'd6375;
      113096:data<=-16'd6648;
      113097:data<=-16'd6593;
      113098:data<=-16'd6437;
      113099:data<=-16'd6663;
      113100:data<=-16'd6930;
      113101:data<=-16'd6760;
      113102:data<=-16'd5962;
      113103:data<=-16'd6575;
      113104:data<=-16'd8237;
      113105:data<=-16'd8258;
      113106:data<=-16'd7953;
      113107:data<=-16'd8131;
      113108:data<=-16'd7670;
      113109:data<=-16'd7521;
      113110:data<=-16'd7602;
      113111:data<=-16'd7224;
      113112:data<=-16'd7003;
      113113:data<=-16'd7065;
      113114:data<=-16'd7134;
      113115:data<=-16'd6777;
      113116:data<=-16'd6883;
      113117:data<=-16'd8032;
      113118:data<=-16'd8301;
      113119:data<=-16'd7953;
      113120:data<=-16'd8109;
      113121:data<=-16'd7752;
      113122:data<=-16'd7486;
      113123:data<=-16'd7530;
      113124:data<=-16'd7100;
      113125:data<=-16'd7080;
      113126:data<=-16'd7053;
      113127:data<=-16'd6593;
      113128:data<=-16'd6661;
      113129:data<=-16'd6986;
      113130:data<=-16'd7571;
      113131:data<=-16'd8185;
      113132:data<=-16'd8005;
      113133:data<=-16'd7803;
      113134:data<=-16'd7676;
      113135:data<=-16'd7122;
      113136:data<=-16'd6740;
      113137:data<=-16'd6584;
      113138:data<=-16'd6642;
      113139:data<=-16'd6851;
      113140:data<=-16'd6537;
      113141:data<=-16'd5984;
      113142:data<=-16'd5970;
      113143:data<=-16'd6640;
      113144:data<=-16'd7568;
      113145:data<=-16'd7558;
      113146:data<=-16'd5553;
      113147:data<=-16'd3016;
      113148:data<=-16'd2420;
      113149:data<=-16'd2494;
      113150:data<=-16'd1630;
      113151:data<=-16'd1697;
      113152:data<=-16'd2361;
      113153:data<=-16'd2096;
      113154:data<=-16'd1924;
      113155:data<=-16'd1738;
      113156:data<=-16'd2096;
      113157:data<=-16'd3829;
      113158:data<=-16'd4329;
      113159:data<=-16'd3422;
      113160:data<=-16'd3256;
      113161:data<=-16'd3134;
      113162:data<=-16'd2834;
      113163:data<=-16'd2886;
      113164:data<=-16'd2740;
      113165:data<=-16'd2523;
      113166:data<=-16'd2617;
      113167:data<=-16'd2679;
      113168:data<=-16'd2315;
      113169:data<=-16'd2591;
      113170:data<=-16'd4029;
      113171:data<=-16'd4552;
      113172:data<=-16'd4087;
      113173:data<=-16'd3950;
      113174:data<=-16'd3465;
      113175:data<=-16'd3203;
      113176:data<=-16'd3447;
      113177:data<=-16'd3046;
      113178:data<=-16'd2649;
      113179:data<=-16'd2528;
      113180:data<=-16'd2431;
      113181:data<=-16'd2547;
      113182:data<=-16'd2657;
      113183:data<=-16'd3427;
      113184:data<=-16'd4128;
      113185:data<=-16'd3679;
      113186:data<=-16'd3560;
      113187:data<=-16'd3621;
      113188:data<=-16'd3187;
      113189:data<=-16'd3057;
      113190:data<=-16'd2883;
      113191:data<=-16'd2667;
      113192:data<=-16'd2275;
      113193:data<=-16'd1788;
      113194:data<=-16'd2126;
      113195:data<=-16'd2152;
      113196:data<=-16'd2648;
      113197:data<=-16'd4231;
      113198:data<=-16'd3933;
      113199:data<=-16'd4331;
      113200:data<=-16'd7379;
      113201:data<=-16'd7906;
      113202:data<=-16'd6619;
      113203:data<=-16'd6742;
      113204:data<=-16'd6272;
      113205:data<=-16'd5580;
      113206:data<=-16'd5823;
      113207:data<=-16'd5515;
      113208:data<=-16'd4664;
      113209:data<=-16'd4740;
      113210:data<=-16'd6096;
      113211:data<=-16'd6652;
      113212:data<=-16'd5611;
      113213:data<=-16'd5054;
      113214:data<=-16'd5027;
      113215:data<=-16'd4737;
      113216:data<=-16'd4323;
      113217:data<=-16'd3439;
      113218:data<=-16'd3002;
      113219:data<=-16'd3186;
      113220:data<=-16'd2792;
      113221:data<=-16'd2270;
      113222:data<=-16'd2267;
      113223:data<=-16'd3075;
      113224:data<=-16'd4064;
      113225:data<=-16'd3706;
      113226:data<=-16'd2869;
      113227:data<=-16'd2588;
      113228:data<=-16'd2259;
      113229:data<=-16'd2061;
      113230:data<=-16'd1932;
      113231:data<=-16'd1557;
      113232:data<=-16'd1151;
      113233:data<=-16'd837;
      113234:data<=-16'd754;
      113235:data<=-16'd629;
      113236:data<=-16'd1064;
      113237:data<=-16'd2309;
      113238:data<=-16'd2460;
      113239:data<=-16'd1748;
      113240:data<=-16'd1538;
      113241:data<=-16'd1143;
      113242:data<=-16'd883;
      113243:data<=-16'd870;
      113244:data<=-16'd384;
      113245:data<=-16'd115;
      113246:data<=16'd96;
      113247:data<=16'd505;
      113248:data<=16'd406;
      113249:data<=16'd33;
      113250:data<=-16'd817;
      113251:data<=-16'd1469;
      113252:data<=16'd276;
      113253:data<=16'd3157;
      113254:data<=16'd4102;
      113255:data<=16'd3756;
      113256:data<=16'd4034;
      113257:data<=16'd4469;
      113258:data<=16'd4437;
      113259:data<=16'd4358;
      113260:data<=16'd4356;
      113261:data<=16'd4496;
      113262:data<=16'd3906;
      113263:data<=16'd2190;
      113264:data<=16'd1753;
      113265:data<=16'd2635;
      113266:data<=16'd2429;
      113267:data<=16'd2094;
      113268:data<=16'd2417;
      113269:data<=16'd2469;
      113270:data<=16'd2729;
      113271:data<=16'd2857;
      113272:data<=16'd2370;
      113273:data<=16'd2326;
      113274:data<=16'd2846;
      113275:data<=16'd2681;
      113276:data<=16'd1239;
      113277:data<=16'd253;
      113278:data<=16'd613;
      113279:data<=16'd716;
      113280:data<=16'd864;
      113281:data<=16'd1365;
      113282:data<=16'd1240;
      113283:data<=16'd1528;
      113284:data<=16'd2021;
      113285:data<=16'd1739;
      113286:data<=16'd1606;
      113287:data<=16'd1592;
      113288:data<=16'd1606;
      113289:data<=16'd1257;
      113290:data<=16'd99;
      113291:data<=-16'd89;
      113292:data<=16'd282;
      113293:data<=16'd100;
      113294:data<=16'd658;
      113295:data<=16'd1049;
      113296:data<=16'd760;
      113297:data<=16'd1034;
      113298:data<=16'd1248;
      113299:data<=16'd1228;
      113300:data<=16'd1224;
      113301:data<=16'd1293;
      113302:data<=16'd1545;
      113303:data<=16'd1480;
      113304:data<=16'd1891;
      113305:data<=16'd1268;
      113306:data<=-16'd1817;
      113307:data<=-16'd2843;
      113308:data<=-16'd1571;
      113309:data<=-16'd1642;
      113310:data<=-16'd1600;
      113311:data<=-16'd1246;
      113312:data<=-16'd1127;
      113313:data<=-16'd560;
      113314:data<=-16'd995;
      113315:data<=-16'd596;
      113316:data<=16'd1539;
      113317:data<=16'd2099;
      113318:data<=16'd2040;
      113319:data<=16'd2400;
      113320:data<=16'd1991;
      113321:data<=16'd2102;
      113322:data<=16'd2537;
      113323:data<=16'd2591;
      113324:data<=16'd3347;
      113325:data<=16'd4482;
      113326:data<=16'd4910;
      113327:data<=16'd4452;
      113328:data<=16'd4783;
      113329:data<=16'd6275;
      113330:data<=16'd6660;
      113331:data<=16'd6534;
      113332:data<=16'd6760;
      113333:data<=16'd6316;
      113334:data<=16'd6182;
      113335:data<=16'd6272;
      113336:data<=16'd5911;
      113337:data<=16'd5915;
      113338:data<=16'd5839;
      113339:data<=16'd5765;
      113340:data<=16'd5685;
      113341:data<=16'd5398;
      113342:data<=16'd6372;
      113343:data<=16'd7368;
      113344:data<=16'd7054;
      113345:data<=16'd6904;
      113346:data<=16'd6681;
      113347:data<=16'd6560;
      113348:data<=16'd6886;
      113349:data<=16'd6484;
      113350:data<=16'd6094;
      113351:data<=16'd6021;
      113352:data<=16'd5920;
      113353:data<=16'd5943;
      113354:data<=16'd5275;
      113355:data<=16'd5611;
      113356:data<=16'd7360;
      113357:data<=16'd7394;
      113358:data<=16'd7050;
      113359:data<=16'd8166;
      113360:data<=16'd8672;
      113361:data<=16'd8370;
      113362:data<=16'd8069;
      113363:data<=16'd7785;
      113364:data<=16'd7621;
      113365:data<=16'd7354;
      113366:data<=16'd7086;
      113367:data<=16'd6608;
      113368:data<=16'd6467;
      113369:data<=16'd7507;
      113370:data<=16'd8164;
      113371:data<=16'd7794;
      113372:data<=16'd7400;
      113373:data<=16'd6939;
      113374:data<=16'd6473;
      113375:data<=16'd6146;
      113376:data<=16'd6146;
      113377:data<=16'd6182;
      113378:data<=16'd5500;
      113379:data<=16'd5203;
      113380:data<=16'd5307;
      113381:data<=16'd4852;
      113382:data<=16'd5350;
      113383:data<=16'd6401;
      113384:data<=16'd6216;
      113385:data<=16'd5600;
      113386:data<=16'd5289;
      113387:data<=16'd5215;
      113388:data<=16'd5010;
      113389:data<=16'd4711;
      113390:data<=16'd4842;
      113391:data<=16'd4470;
      113392:data<=16'd3938;
      113393:data<=16'd3842;
      113394:data<=16'd3109;
      113395:data<=16'd3576;
      113396:data<=16'd5426;
      113397:data<=16'd5292;
      113398:data<=16'd4369;
      113399:data<=16'd4463;
      113400:data<=16'd4232;
      113401:data<=16'd3779;
      113402:data<=16'd3547;
      113403:data<=16'd3366;
      113404:data<=16'd3165;
      113405:data<=16'd2866;
      113406:data<=16'd2617;
      113407:data<=16'd2097;
      113408:data<=16'd2538;
      113409:data<=16'd4432;
      113410:data<=16'd4769;
      113411:data<=16'd3368;
      113412:data<=16'd2206;
      113413:data<=16'd1199;
      113414:data<=16'd839;
      113415:data<=16'd905;
      113416:data<=16'd576;
      113417:data<=16'd487;
      113418:data<=16'd546;
      113419:data<=16'd543;
      113420:data<=16'd390;
      113421:data<=16'd359;
      113422:data<=16'd1527;
      113423:data<=16'd2453;
      113424:data<=16'd2026;
      113425:data<=16'd1665;
      113426:data<=16'd1322;
      113427:data<=16'd1034;
      113428:data<=16'd1181;
      113429:data<=16'd1022;
      113430:data<=16'd834;
      113431:data<=16'd764;
      113432:data<=16'd710;
      113433:data<=16'd673;
      113434:data<=16'd411;
      113435:data<=16'd1187;
      113436:data<=16'd2366;
      113437:data<=16'd2153;
      113438:data<=16'd2067;
      113439:data<=16'd2108;
      113440:data<=16'd1257;
      113441:data<=16'd842;
      113442:data<=16'd691;
      113443:data<=16'd414;
      113444:data<=16'd334;
      113445:data<=16'd36;
      113446:data<=-16'd42;
      113447:data<=-16'd50;
      113448:data<=16'd223;
      113449:data<=16'd1410;
      113450:data<=16'd1807;
      113451:data<=16'd1495;
      113452:data<=16'd1641;
      113453:data<=16'd1098;
      113454:data<=16'd318;
      113455:data<=16'd196;
      113456:data<=16'd132;
      113457:data<=16'd67;
      113458:data<=-16'd226;
      113459:data<=-16'd488;
      113460:data<=-16'd452;
      113461:data<=-16'd162;
      113462:data<=16'd1002;
      113463:data<=16'd1656;
      113464:data<=16'd1207;
      113465:data<=16'd1871;
      113466:data<=16'd2880;
      113467:data<=16'd2673;
      113468:data<=16'd2290;
      113469:data<=16'd1888;
      113470:data<=16'd1278;
      113471:data<=16'd1016;
      113472:data<=16'd1005;
      113473:data<=16'd704;
      113474:data<=16'd506;
      113475:data<=16'd1551;
      113476:data<=16'd2641;
      113477:data<=16'd2209;
      113478:data<=16'd1657;
      113479:data<=16'd1560;
      113480:data<=16'd1177;
      113481:data<=16'd807;
      113482:data<=16'd500;
      113483:data<=16'd168;
      113484:data<=-16'd194;
      113485:data<=-16'd244;
      113486:data<=16'd35;
      113487:data<=-16'd417;
      113488:data<=-16'd329;
      113489:data<=16'd1121;
      113490:data<=16'd1260;
      113491:data<=16'd417;
      113492:data<=16'd409;
      113493:data<=16'd117;
      113494:data<=-16'd443;
      113495:data<=-16'd509;
      113496:data<=-16'd567;
      113497:data<=-16'd782;
      113498:data<=-16'd963;
      113499:data<=-16'd993;
      113500:data<=-16'd1254;
      113501:data<=-16'd1028;
      113502:data<=16'd227;
      113503:data<=16'd296;
      113504:data<=-16'd453;
      113505:data<=-16'd17;
      113506:data<=-16'd82;
      113507:data<=-16'd914;
      113508:data<=-16'd1133;
      113509:data<=-16'd1310;
      113510:data<=-16'd1281;
      113511:data<=-16'd1145;
      113512:data<=-16'd1585;
      113513:data<=-16'd1871;
      113514:data<=-16'd1732;
      113515:data<=-16'd1701;
      113516:data<=-16'd2012;
      113517:data<=-16'd2221;
      113518:data<=-16'd2605;
      113519:data<=-16'd4040;
      113520:data<=-16'd4878;
      113521:data<=-16'd4742;
      113522:data<=-16'd5301;
      113523:data<=-16'd5053;
      113524:data<=-16'd4335;
      113525:data<=-16'd4992;
      113526:data<=-16'd5031;
      113527:data<=-16'd4893;
      113528:data<=-16'd6000;
      113529:data<=-16'd6511;
      113530:data<=-16'd6560;
      113531:data<=-16'd6633;
      113532:data<=-16'd6273;
      113533:data<=-16'd6241;
      113534:data<=-16'd6260;
      113535:data<=-16'd6304;
      113536:data<=-16'd6504;
      113537:data<=-16'd6170;
      113538:data<=-16'd6056;
      113539:data<=-16'd5888;
      113540:data<=-16'd5344;
      113541:data<=-16'd6111;
      113542:data<=-16'd7350;
      113543:data<=-16'd7386;
      113544:data<=-16'd7048;
      113545:data<=-16'd7066;
      113546:data<=-16'd7109;
      113547:data<=-16'd6818;
      113548:data<=-16'd6760;
      113549:data<=-16'd6983;
      113550:data<=-16'd6687;
      113551:data<=-16'd6479;
      113552:data<=-16'd6094;
      113553:data<=-16'd5339;
      113554:data<=-16'd6159;
      113555:data<=-16'd7676;
      113556:data<=-16'd7894;
      113557:data<=-16'd7439;
      113558:data<=-16'd6852;
      113559:data<=-16'd6683;
      113560:data<=-16'd6804;
      113561:data<=-16'd6561;
      113562:data<=-16'd6546;
      113563:data<=-16'd6308;
      113564:data<=-16'd5912;
      113565:data<=-16'd5900;
      113566:data<=-16'd5245;
      113567:data<=-16'd5295;
      113568:data<=-16'd6786;
      113569:data<=-16'd7574;
      113570:data<=-16'd7626;
      113571:data<=-16'd6522;
      113572:data<=-16'd4379;
      113573:data<=-16'd3906;
      113574:data<=-16'd4338;
      113575:data<=-16'd4070;
      113576:data<=-16'd3871;
      113577:data<=-16'd3597;
      113578:data<=-16'd3500;
      113579:data<=-16'd3492;
      113580:data<=-16'd3397;
      113581:data<=-16'd4413;
      113582:data<=-16'd5266;
      113583:data<=-16'd4911;
      113584:data<=-16'd4927;
      113585:data<=-16'd4954;
      113586:data<=-16'd4452;
      113587:data<=-16'd4249;
      113588:data<=-16'd4299;
      113589:data<=-16'd4264;
      113590:data<=-16'd3838;
      113591:data<=-16'd3462;
      113592:data<=-16'd3428;
      113593:data<=-16'd3201;
      113594:data<=-16'd3865;
      113595:data<=-16'd5280;
      113596:data<=-16'd5285;
      113597:data<=-16'd4799;
      113598:data<=-16'd5039;
      113599:data<=-16'd4723;
      113600:data<=-16'd4064;
      113601:data<=-16'd3958;
      113602:data<=-16'd3676;
      113603:data<=-16'd3233;
      113604:data<=-16'd3422;
      113605:data<=-16'd3228;
      113606:data<=-16'd2317;
      113607:data<=-16'd2898;
      113608:data<=-16'd4684;
      113609:data<=-16'd5119;
      113610:data<=-16'd4520;
      113611:data<=-16'd4108;
      113612:data<=-16'd3914;
      113613:data<=-16'd3861;
      113614:data<=-16'd3609;
      113615:data<=-16'd3280;
      113616:data<=-16'd3016;
      113617:data<=-16'd2789;
      113618:data<=-16'd2886;
      113619:data<=-16'd2479;
      113620:data<=-16'd2220;
      113621:data<=-16'd3964;
      113622:data<=-16'd5344;
      113623:data<=-16'd4402;
      113624:data<=-16'd3950;
      113625:data<=-16'd4990;
      113626:data<=-16'd5495;
      113627:data<=-16'd5140;
      113628:data<=-16'd4836;
      113629:data<=-16'd4408;
      113630:data<=-16'd3682;
      113631:data<=-16'd3500;
      113632:data<=-16'd3613;
      113633:data<=-16'd3368;
      113634:data<=-16'd3897;
      113635:data<=-16'd5031;
      113636:data<=-16'd4983;
      113637:data<=-16'd4206;
      113638:data<=-16'd3802;
      113639:data<=-16'd3318;
      113640:data<=-16'd2675;
      113641:data<=-16'd2457;
      113642:data<=-16'd2355;
      113643:data<=-16'd1856;
      113644:data<=-16'd1589;
      113645:data<=-16'd1588;
      113646:data<=-16'd1180;
      113647:data<=-16'd1400;
      113648:data<=-16'd2544;
      113649:data<=-16'd2823;
      113650:data<=-16'd2240;
      113651:data<=-16'd1959;
      113652:data<=-16'd1736;
      113653:data<=-16'd1298;
      113654:data<=-16'd911;
      113655:data<=-16'd694;
      113656:data<=-16'd600;
      113657:data<=-16'd375;
      113658:data<=16'd147;
      113659:data<=16'd544;
      113660:data<=16'd41;
      113661:data<=-16'd1140;
      113662:data<=-16'd1695;
      113663:data<=-16'd1312;
      113664:data<=-16'd814;
      113665:data<=-16'd552;
      113666:data<=-16'd300;
      113667:data<=16'd55;
      113668:data<=16'd409;
      113669:data<=16'd570;
      113670:data<=16'd550;
      113671:data<=16'd937;
      113672:data<=16'd1663;
      113673:data<=16'd1377;
      113674:data<=16'd180;
      113675:data<=-16'd520;
      113676:data<=-16'd513;
      113677:data<=16'd478;
      113678:data<=16'd2096;
      113679:data<=16'd2707;
      113680:data<=16'd2679;
      113681:data<=16'd2922;
      113682:data<=16'd3072;
      113683:data<=16'd3171;
      113684:data<=16'd2930;
      113685:data<=16'd2899;
      113686:data<=16'd3700;
      113687:data<=16'd3154;
      113688:data<=16'd1398;
      113689:data<=16'd1187;
      113690:data<=16'd1574;
      113691:data<=16'd1292;
      113692:data<=16'd1492;
      113693:data<=16'd1985;
      113694:data<=16'd2049;
      113695:data<=16'd2120;
      113696:data<=16'd2423;
      113697:data<=16'd2470;
      113698:data<=16'd2396;
      113699:data<=16'd2726;
      113700:data<=16'd2200;
      113701:data<=16'd705;
      113702:data<=16'd597;
      113703:data<=16'd1151;
      113704:data<=16'd719;
      113705:data<=16'd811;
      113706:data<=16'd1521;
      113707:data<=16'd1624;
      113708:data<=16'd1656;
      113709:data<=16'd1792;
      113710:data<=16'd1729;
      113711:data<=16'd1838;
      113712:data<=16'd2223;
      113713:data<=16'd1932;
      113714:data<=16'd496;
      113715:data<=-16'd129;
      113716:data<=16'd676;
      113717:data<=16'd793;
      113718:data<=16'd469;
      113719:data<=16'd848;
      113720:data<=16'd1148;
      113721:data<=16'd1289;
      113722:data<=16'd1375;
      113723:data<=16'd1345;
      113724:data<=16'd1569;
      113725:data<=16'd1662;
      113726:data<=16'd1820;
      113727:data<=16'd2090;
      113728:data<=16'd1832;
      113729:data<=16'd2027;
      113730:data<=16'd2176;
      113731:data<=16'd738;
      113732:data<=-16'd343;
      113733:data<=16'd100;
      113734:data<=16'd582;
      113735:data<=16'd795;
      113736:data<=16'd907;
      113737:data<=16'd1021;
      113738:data<=16'd1137;
      113739:data<=16'd1102;
      113740:data<=16'd1944;
      113741:data<=16'd3278;
      113742:data<=16'd3410;
      113743:data<=16'd3169;
      113744:data<=16'd3513;
      113745:data<=16'd3767;
      113746:data<=16'd3894;
      113747:data<=16'd4037;
      113748:data<=16'd3938;
      113749:data<=16'd3814;
      113750:data<=16'd4065;
      113751:data<=16'd4115;
      113752:data<=16'd3504;
      113753:data<=16'd3943;
      113754:data<=16'd5642;
      113755:data<=16'd5927;
      113756:data<=16'd5087;
      113757:data<=16'd5071;
      113758:data<=16'd5194;
      113759:data<=16'd5115;
      113760:data<=16'd5259;
      113761:data<=16'd5075;
      113762:data<=16'd4784;
      113763:data<=16'd5001;
      113764:data<=16'd5113;
      113765:data<=16'd4640;
      113766:data<=16'd4693;
      113767:data<=16'd5839;
      113768:data<=16'd6557;
      113769:data<=16'd6387;
      113770:data<=16'd6332;
      113771:data<=16'd6203;
      113772:data<=16'd5823;
      113773:data<=16'd5714;
      113774:data<=16'd5880;
      113775:data<=16'd5887;
      113776:data<=16'd5351;
      113777:data<=16'd4984;
      113778:data<=16'd5134;
      113779:data<=16'd4890;
      113780:data<=16'd5127;
      113781:data<=16'd6396;
      113782:data<=16'd6599;
      113783:data<=16'd6061;
      113784:data<=16'd6875;
      113785:data<=16'd7843;
      113786:data<=16'd7588;
      113787:data<=16'd7526;
      113788:data<=16'd7782;
      113789:data<=16'd7078;
      113790:data<=16'd6464;
      113791:data<=16'd6391;
      113792:data<=16'd5820;
      113793:data<=16'd6361;
      113794:data<=16'd7962;
      113795:data<=16'd7694;
      113796:data<=16'd6751;
      113797:data<=16'd6893;
      113798:data<=16'd6687;
      113799:data<=16'd6185;
      113800:data<=16'd5988;
      113801:data<=16'd5843;
      113802:data<=16'd5820;
      113803:data<=16'd5459;
      113804:data<=16'd4908;
      113805:data<=16'd4673;
      113806:data<=16'd5025;
      113807:data<=16'd6199;
      113808:data<=16'd6522;
      113809:data<=16'd5650;
      113810:data<=16'd5568;
      113811:data<=16'd5682;
      113812:data<=16'd5271;
      113813:data<=16'd5195;
      113814:data<=16'd4901;
      113815:data<=16'd4366;
      113816:data<=16'd4300;
      113817:data<=16'd4237;
      113818:data<=16'd3768;
      113819:data<=16'd3532;
      113820:data<=16'd4476;
      113821:data<=16'd5504;
      113822:data<=16'd5100;
      113823:data<=16'd4452;
      113824:data<=16'd4270;
      113825:data<=16'd4049;
      113826:data<=16'd4026;
      113827:data<=16'd3797;
      113828:data<=16'd3230;
      113829:data<=16'd2995;
      113830:data<=16'd3058;
      113831:data<=16'd2833;
      113832:data<=16'd2349;
      113833:data<=16'd3131;
      113834:data<=16'd4592;
      113835:data<=16'd4487;
      113836:data<=16'd4121;
      113837:data<=16'd3550;
      113838:data<=16'd1450;
      113839:data<=16'd675;
      113840:data<=16'd1363;
      113841:data<=16'd987;
      113842:data<=16'd599;
      113843:data<=16'd459;
      113844:data<=16'd147;
      113845:data<=16'd196;
      113846:data<=16'd414;
      113847:data<=16'd1463;
      113848:data<=16'd2359;
      113849:data<=16'd1927;
      113850:data<=16'd1814;
      113851:data<=16'd1513;
      113852:data<=16'd785;
      113853:data<=16'd1115;
      113854:data<=16'd1092;
      113855:data<=16'd613;
      113856:data<=16'd708;
      113857:data<=16'd218;
      113858:data<=-16'd291;
      113859:data<=16'd296;
      113860:data<=16'd1562;
      113861:data<=16'd2446;
      113862:data<=16'd1835;
      113863:data<=16'd1230;
      113864:data<=16'd1545;
      113865:data<=16'd1290;
      113866:data<=16'd972;
      113867:data<=16'd763;
      113868:data<=16'd100;
      113869:data<=16'd127;
      113870:data<=16'd235;
      113871:data<=-16'd384;
      113872:data<=-16'd305;
      113873:data<=16'd755;
      113874:data<=16'd1635;
      113875:data<=16'd1627;
      113876:data<=16'd1213;
      113877:data<=16'd1054;
      113878:data<=16'd933;
      113879:data<=16'd854;
      113880:data<=16'd576;
      113881:data<=-16'd77;
      113882:data<=-16'd370;
      113883:data<=-16'd282;
      113884:data<=-16'd232;
      113885:data<=-16'd519;
      113886:data<=-16'd516;
      113887:data<=16'd855;
      113888:data<=16'd1545;
      113889:data<=16'd743;
      113890:data<=16'd1359;
      113891:data<=16'd2570;
      113892:data<=16'd2458;
      113893:data<=16'd2211;
      113894:data<=16'd1663;
      113895:data<=16'd920;
      113896:data<=16'd1013;
      113897:data<=16'd975;
      113898:data<=16'd555;
      113899:data<=16'd913;
      113900:data<=16'd2011;
      113901:data<=16'd2416;
      113902:data<=16'd1801;
      113903:data<=16'd1688;
      113904:data<=16'd1715;
      113905:data<=16'd966;
      113906:data<=16'd625;
      113907:data<=16'd532;
      113908:data<=16'd177;
      113909:data<=16'd200;
      113910:data<=-16'd71;
      113911:data<=-16'd682;
      113912:data<=-16'd302;
      113913:data<=16'd1017;
      113914:data<=16'd1626;
      113915:data<=16'd933;
      113916:data<=16'd647;
      113917:data<=16'd899;
      113918:data<=16'd426;
      113919:data<=16'd97;
      113920:data<=-16'd20;
      113921:data<=-16'd381;
      113922:data<=-16'd308;
      113923:data<=-16'd625;
      113924:data<=-16'd1301;
      113925:data<=-16'd1099;
      113926:data<=-16'd250;
      113927:data<=16'd654;
      113928:data<=16'd470;
      113929:data<=-16'd437;
      113930:data<=-16'd311;
      113931:data<=-16'd183;
      113932:data<=-16'd591;
      113933:data<=-16'd749;
      113934:data<=-16'd1228;
      113935:data<=-16'd1491;
      113936:data<=-16'd1303;
      113937:data<=-16'd1465;
      113938:data<=-16'd1724;
      113939:data<=-16'd2137;
      113940:data<=-16'd2314;
      113941:data<=-16'd2056;
      113942:data<=-16'd2246;
      113943:data<=-16'd2964;
      113944:data<=-16'd4287;
      113945:data<=-16'd5147;
      113946:data<=-16'd4869;
      113947:data<=-16'd5286;
      113948:data<=-16'd5661;
      113949:data<=-16'd5160;
      113950:data<=-16'd5130;
      113951:data<=-16'd4852;
      113952:data<=-16'd5394;
      113953:data<=-16'd7322;
      113954:data<=-16'd7470;
      113955:data<=-16'd6637;
      113956:data<=-16'd6678;
      113957:data<=-16'd6639;
      113958:data<=-16'd6836;
      113959:data<=-16'd6957;
      113960:data<=-16'd6701;
      113961:data<=-16'd6673;
      113962:data<=-16'd6616;
      113963:data<=-16'd6787;
      113964:data<=-16'd6510;
      113965:data<=-16'd6238;
      113966:data<=-16'd7656;
      113967:data<=-16'd8537;
      113968:data<=-16'd8181;
      113969:data<=-16'd8161;
      113970:data<=-16'd7602;
      113971:data<=-16'd7403;
      113972:data<=-16'd7944;
      113973:data<=-16'd7620;
      113974:data<=-16'd7213;
      113975:data<=-16'd6986;
      113976:data<=-16'd6940;
      113977:data<=-16'd7174;
      113978:data<=-16'd6705;
      113979:data<=-16'd7018;
      113980:data<=-16'd8129;
      113981:data<=-16'd8105;
      113982:data<=-16'd8026;
      113983:data<=-16'd7959;
      113984:data<=-16'd7421;
      113985:data<=-16'd7304;
      113986:data<=-16'd7244;
      113987:data<=-16'd7330;
      113988:data<=-16'd7138;
      113989:data<=-16'd6482;
      113990:data<=-16'd6555;
      113991:data<=-16'd6367;
      113992:data<=-16'd6464;
      113993:data<=-16'd7749;
      113994:data<=-16'd7814;
      113995:data<=-16'd7382;
      113996:data<=-16'd7219;
      113997:data<=-16'd5547;
      113998:data<=-16'd4138;
      113999:data<=-16'd4206;
      114000:data<=-16'd4451;
      114001:data<=-16'd4478;
      114002:data<=-16'd4178;
      114003:data<=-16'd4009;
      114004:data<=-16'd3629;
      114005:data<=-16'd3547;
      114006:data<=-16'd5128;
      114007:data<=-16'd5783;
      114008:data<=-16'd4868;
      114009:data<=-16'd4881;
      114010:data<=-16'd4934;
      114011:data<=-16'd4655;
      114012:data<=-16'd4608;
      114013:data<=-16'd4294;
      114014:data<=-16'd4317;
      114015:data<=-16'd4299;
      114016:data<=-16'd3968;
      114017:data<=-16'd3577;
      114018:data<=-16'd3137;
      114019:data<=-16'd4285;
      114020:data<=-16'd5636;
      114021:data<=-16'd5133;
      114022:data<=-16'd4848;
      114023:data<=-16'd4686;
      114024:data<=-16'd4134;
      114025:data<=-16'd4253;
      114026:data<=-16'd4009;
      114027:data<=-16'd3647;
      114028:data<=-16'd3495;
      114029:data<=-16'd3198;
      114030:data<=-16'd3322;
      114031:data<=-16'd2764;
      114032:data<=-16'd2893;
      114033:data<=-16'd4660;
      114034:data<=-16'd4666;
      114035:data<=-16'd4108;
      114036:data<=-16'd4411;
      114037:data<=-16'd3604;
      114038:data<=-16'd3456;
      114039:data<=-16'd3836;
      114040:data<=-16'd3071;
      114041:data<=-16'd2814;
      114042:data<=-16'd2872;
      114043:data<=-16'd2704;
      114044:data<=-16'd2552;
      114045:data<=-16'd2770;
      114046:data<=-16'd4411;
      114047:data<=-16'd4827;
      114048:data<=-16'd3542;
      114049:data<=-16'd4206;
      114050:data<=-16'd5309;
      114051:data<=-16'd5231;
      114052:data<=-16'd5218;
      114053:data<=-16'd4825;
      114054:data<=-16'd4651;
      114055:data<=-16'd4625;
      114056:data<=-16'd3833;
      114057:data<=-16'd3391;
      114058:data<=-16'd3826;
      114059:data<=-16'd4992;
      114060:data<=-16'd5480;
      114061:data<=-16'd4563;
      114062:data<=-16'd4428;
      114063:data<=-16'd4496;
      114064:data<=-16'd3748;
      114065:data<=-16'd3571;
      114066:data<=-16'd3153;
      114067:data<=-16'd2631;
      114068:data<=-16'd2840;
      114069:data<=-16'd2537;
      114070:data<=-16'd2021;
      114071:data<=-16'd1902;
      114072:data<=-16'd2505;
      114073:data<=-16'd3613;
      114074:data<=-16'd3369;
      114075:data<=-16'd2748;
      114076:data<=-16'd2799;
      114077:data<=-16'd2340;
      114078:data<=-16'd2191;
      114079:data<=-16'd2170;
      114080:data<=-16'd1528;
      114081:data<=-16'd1342;
      114082:data<=-16'd1300;
      114083:data<=-16'd1140;
      114084:data<=-16'd886;
      114085:data<=-16'd866;
      114086:data<=-16'd2099;
      114087:data<=-16'd2610;
      114088:data<=-16'd1811;
      114089:data<=-16'd1704;
      114090:data<=-16'd1407;
      114091:data<=-16'd998;
      114092:data<=-16'd1221;
      114093:data<=-16'd790;
      114094:data<=-16'd217;
      114095:data<=-16'd21;
      114096:data<=16'd271;
      114097:data<=16'd472;
      114098:data<=16'd194;
      114099:data<=-16'd957;
      114100:data<=-16'd1201;
      114101:data<=-16'd393;
      114102:data<=-16'd708;
      114103:data<=16'd80;
      114104:data<=16'd2111;
      114105:data<=16'd2190;
      114106:data<=16'd2102;
      114107:data<=16'd2610;
      114108:data<=16'd2409;
      114109:data<=16'd2666;
      114110:data<=16'd2971;
      114111:data<=16'd2551;
      114112:data<=16'd1704;
      114113:data<=16'd1011;
      114114:data<=16'd1456;
      114115:data<=16'd1503;
      114116:data<=16'd920;
      114117:data<=16'd1495;
      114118:data<=16'd1929;
      114119:data<=16'd1874;
      114120:data<=16'd2147;
      114121:data<=16'd2115;
      114122:data<=16'd2235;
      114123:data<=16'd2569;
      114124:data<=16'd2833;
      114125:data<=16'd2369;
      114126:data<=16'd640;
      114127:data<=16'd346;
      114128:data<=16'd1322;
      114129:data<=16'd963;
      114130:data<=16'd964;
      114131:data<=16'd1462;
      114132:data<=16'd1327;
      114133:data<=16'd1795;
      114134:data<=16'd2055;
      114135:data<=16'd1800;
      114136:data<=16'd2196;
      114137:data<=16'd2619;
      114138:data<=16'd2132;
      114139:data<=16'd679;
      114140:data<=16'd115;
      114141:data<=16'd749;
      114142:data<=16'd657;
      114143:data<=16'd1025;
      114144:data<=16'd1741;
      114145:data<=16'd1306;
      114146:data<=16'd1488;
      114147:data<=16'd1789;
      114148:data<=16'd1544;
      114149:data<=16'd2008;
      114150:data<=16'd1945;
      114151:data<=16'd1874;
      114152:data<=16'd2478;
      114153:data<=16'd2209;
      114154:data<=16'd2193;
      114155:data<=16'd2475;
      114156:data<=16'd1727;
      114157:data<=16'd899;
      114158:data<=16'd447;
      114159:data<=16'd620;
      114160:data<=16'd949;
      114161:data<=16'd920;
      114162:data<=16'd1580;
      114163:data<=16'd1836;
      114164:data<=16'd1718;
      114165:data<=16'd2992;
      114166:data<=16'd3940;
      114167:data<=16'd3983;
      114168:data<=16'd4114;
      114169:data<=16'd3845;
      114170:data<=16'd3827;
      114171:data<=16'd4064;
      114172:data<=16'd4168;
      114173:data<=16'd4278;
      114174:data<=16'd3836;
      114175:data<=16'd3876;
      114176:data<=16'd4106;
      114177:data<=16'd3536;
      114178:data<=16'd4375;
      114179:data<=16'd6003;
      114180:data<=16'd6214;
      114181:data<=16'd6155;
      114182:data<=16'd6170;
      114183:data<=16'd5906;
      114184:data<=16'd5726;
      114185:data<=16'd5764;
      114186:data<=16'd5873;
      114187:data<=16'd5374;
      114188:data<=16'd5178;
      114189:data<=16'd5342;
      114190:data<=16'd4686;
      114191:data<=16'd5353;
      114192:data<=16'd7048;
      114193:data<=16'd7033;
      114194:data<=16'd6777;
      114195:data<=16'd6836;
      114196:data<=16'd6426;
      114197:data<=16'd6313;
      114198:data<=16'd6164;
      114199:data<=16'd6181;
      114200:data<=16'd6335;
      114201:data<=16'd6006;
      114202:data<=16'd5827;
      114203:data<=16'd5503;
      114204:data<=16'd5770;
      114205:data<=16'd7177;
      114206:data<=16'd7576;
      114207:data<=16'd7078;
      114208:data<=16'd6736;
      114209:data<=16'd7019;
      114210:data<=16'd8376;
      114211:data<=16'd8648;
      114212:data<=16'd8040;
      114213:data<=16'd8140;
      114214:data<=16'd7680;
      114215:data<=16'd7545;
      114216:data<=16'd7530;
      114217:data<=16'd6678;
      114218:data<=16'd7641;
      114219:data<=16'd8913;
      114220:data<=16'd8329;
      114221:data<=16'd8032;
      114222:data<=16'd7609;
      114223:data<=16'd7075;
      114224:data<=16'd7239;
      114225:data<=16'd6798;
      114226:data<=16'd6443;
      114227:data<=16'd6332;
      114228:data<=16'd6015;
      114229:data<=16'd6031;
      114230:data<=16'd5485;
      114231:data<=16'd5683;
      114232:data<=16'd7125;
      114233:data<=16'd7087;
      114234:data<=16'd6545;
      114235:data<=16'd6586;
      114236:data<=16'd6026;
      114237:data<=16'd5609;
      114238:data<=16'd5512;
      114239:data<=16'd5445;
      114240:data<=16'd5438;
      114241:data<=16'd5040;
      114242:data<=16'd4590;
      114243:data<=16'd4111;
      114244:data<=16'd4469;
      114245:data<=16'd5823;
      114246:data<=16'd5721;
      114247:data<=16'd5045;
      114248:data<=16'd5388;
      114249:data<=16'd5096;
      114250:data<=16'd4437;
      114251:data<=16'd4212;
      114252:data<=16'd4030;
      114253:data<=16'd3891;
      114254:data<=16'd3526;
      114255:data<=16'd3274;
      114256:data<=16'd2767;
      114257:data<=16'd2626;
      114258:data<=16'd4472;
      114259:data<=16'd5275;
      114260:data<=16'd4202;
      114261:data<=16'd4394;
      114262:data<=16'd3838;
      114263:data<=16'd1844;
      114264:data<=16'd1333;
      114265:data<=16'd1287;
      114266:data<=16'd843;
      114267:data<=16'd745;
      114268:data<=16'd597;
      114269:data<=16'd281;
      114270:data<=16'd92;
      114271:data<=16'd1039;
      114272:data<=16'd2350;
      114273:data<=16'd2083;
      114274:data<=16'd1597;
      114275:data<=16'd1597;
      114276:data<=16'd1242;
      114277:data<=16'd1260;
      114278:data<=16'd1251;
      114279:data<=16'd741;
      114280:data<=16'd484;
      114281:data<=16'd557;
      114282:data<=16'd654;
      114283:data<=16'd180;
      114284:data<=16'd193;
      114285:data<=16'd1527;
      114286:data<=16'd1967;
      114287:data<=16'd1589;
      114288:data<=16'd1627;
      114289:data<=16'd1045;
      114290:data<=16'd675;
      114291:data<=16'd967;
      114292:data<=16'd544;
      114293:data<=-16'd15;
      114294:data<=-16'd79;
      114295:data<=-16'd62;
      114296:data<=-16'd218;
      114297:data<=-16'd76;
      114298:data<=16'd1077;
      114299:data<=16'd1733;
      114300:data<=16'd1272;
      114301:data<=16'd1257;
      114302:data<=16'd1045;
      114303:data<=16'd393;
      114304:data<=16'd411;
      114305:data<=16'd318;
      114306:data<=-16'd21;
      114307:data<=16'd9;
      114308:data<=-16'd123;
      114309:data<=-16'd459;
      114310:data<=-16'd241;
      114311:data<=16'd881;
      114312:data<=16'd1785;
      114313:data<=16'd1434;
      114314:data<=16'd863;
      114315:data<=16'd1139;
      114316:data<=16'd2017;
      114317:data<=16'd2438;
      114318:data<=16'd2030;
      114319:data<=16'd1823;
      114320:data<=16'd1704;
      114321:data<=16'd1368;
      114322:data<=16'd1154;
      114323:data<=16'd567;
      114324:data<=16'd963;
      114325:data<=16'd2708;
      114326:data<=16'd2801;
      114327:data<=16'd1839;
      114328:data<=16'd1773;
      114329:data<=16'd1453;
      114330:data<=16'd1057;
      114331:data<=16'd1001;
      114332:data<=16'd493;
      114333:data<=16'd112;
      114334:data<=16'd253;
      114335:data<=16'd179;
      114336:data<=-16'd314;
      114337:data<=16'd5;
      114338:data<=16'd1403;
      114339:data<=16'd1771;
      114340:data<=16'd1172;
      114341:data<=16'd999;
      114342:data<=16'd575;
      114343:data<=16'd211;
      114344:data<=16'd212;
      114345:data<=-16'd162;
      114346:data<=-16'd265;
      114347:data<=-16'd250;
      114348:data<=-16'd766;
      114349:data<=-16'd1137;
      114350:data<=-16'd708;
      114351:data<=16'd535;
      114352:data<=16'd995;
      114353:data<=16'd321;
      114354:data<=16'd340;
      114355:data<=16'd299;
      114356:data<=-16'd335;
      114357:data<=-16'd400;
      114358:data<=-16'd594;
      114359:data<=-16'd816;
      114360:data<=-16'd798;
      114361:data<=-16'd1375;
      114362:data<=-16'd1709;
      114363:data<=-16'd1727;
      114364:data<=-16'd1985;
      114365:data<=-16'd2061;
      114366:data<=-16'd2328;
      114367:data<=-16'd2334;
      114368:data<=-16'd2366;
      114369:data<=-16'd3776;
      114370:data<=-16'd5033;
      114371:data<=-16'd5221;
      114372:data<=-16'd5125;
      114373:data<=-16'd4704;
      114374:data<=-16'd4786;
      114375:data<=-16'd4996;
      114376:data<=-16'd4610;
      114377:data<=-16'd5327;
      114378:data<=-16'd6690;
      114379:data<=-16'd6884;
      114380:data<=-16'd6595;
      114381:data<=-16'd6516;
      114382:data<=-16'd6476;
      114383:data<=-16'd6364;
      114384:data<=-16'd6367;
      114385:data<=-16'd6511;
      114386:data<=-16'd6256;
      114387:data<=-16'd6184;
      114388:data<=-16'd6408;
      114389:data<=-16'd6061;
      114390:data<=-16'd6376;
      114391:data<=-16'd7576;
      114392:data<=-16'd7749;
      114393:data<=-16'd7356;
      114394:data<=-16'd7464;
      114395:data<=-16'd7439;
      114396:data<=-16'd7124;
      114397:data<=-16'd6998;
      114398:data<=-16'd6960;
      114399:data<=-16'd6667;
      114400:data<=-16'd6539;
      114401:data<=-16'd6558;
      114402:data<=-16'd6187;
      114403:data<=-16'd6478;
      114404:data<=-16'd7592;
      114405:data<=-16'd7814;
      114406:data<=-16'd7474;
      114407:data<=-16'd7497;
      114408:data<=-16'd7368;
      114409:data<=-16'd7028;
      114410:data<=-16'd6610;
      114411:data<=-16'd6281;
      114412:data<=-16'd6347;
      114413:data<=-16'd6425;
      114414:data<=-16'd6223;
      114415:data<=-16'd5811;
      114416:data<=-16'd5585;
      114417:data<=-16'd6209;
      114418:data<=-16'd7209;
      114419:data<=-16'd7441;
      114420:data<=-16'd6951;
      114421:data<=-16'd6525;
      114422:data<=-16'd5762;
      114423:data<=-16'd4305;
      114424:data<=-16'd3748;
      114425:data<=-16'd4118;
      114426:data<=-16'd3817;
      114427:data<=-16'd3802;
      114428:data<=-16'd4129;
      114429:data<=-16'd3527;
      114430:data<=-16'd3815;
      114431:data<=-16'd5256;
      114432:data<=-16'd5527;
      114433:data<=-16'd5151;
      114434:data<=-16'd4905;
      114435:data<=-16'd4429;
      114436:data<=-16'd4598;
      114437:data<=-16'd5045;
      114438:data<=-16'd4498;
      114439:data<=-16'd3882;
      114440:data<=-16'd4088;
      114441:data<=-16'd4047;
      114442:data<=-16'd3512;
      114443:data<=-16'd3882;
      114444:data<=-16'd5086;
      114445:data<=-16'd5517;
      114446:data<=-16'd5071;
      114447:data<=-16'd4808;
      114448:data<=-16'd4764;
      114449:data<=-16'd4334;
      114450:data<=-16'd3896;
      114451:data<=-16'd3974;
      114452:data<=-16'd3953;
      114453:data<=-16'd3755;
      114454:data<=-16'd3641;
      114455:data<=-16'd3156;
      114456:data<=-16'd3219;
      114457:data<=-16'd4416;
      114458:data<=-16'd5031;
      114459:data<=-16'd4796;
      114460:data<=-16'd4689;
      114461:data<=-16'd4519;
      114462:data<=-16'd4128;
      114463:data<=-16'd3607;
      114464:data<=-16'd3272;
      114465:data<=-16'd3262;
      114466:data<=-16'd3201;
      114467:data<=-16'd3247;
      114468:data<=-16'd2925;
      114469:data<=-16'd2376;
      114470:data<=-16'd3495;
      114471:data<=-16'd5165;
      114472:data<=-16'd5113;
      114473:data<=-16'd4393;
      114474:data<=-16'd3944;
      114475:data<=-16'd4290;
      114476:data<=-16'd5698;
      114477:data<=-16'd6011;
      114478:data<=-16'd4996;
      114479:data<=-16'd4711;
      114480:data<=-16'd4863;
      114481:data<=-16'd4520;
      114482:data<=-16'd3955;
      114483:data<=-16'd4176;
      114484:data<=-16'd5556;
      114485:data<=-16'd6128;
      114486:data<=-16'd5366;
      114487:data<=-16'd4975;
      114488:data<=-16'd4560;
      114489:data<=-16'd3952;
      114490:data<=-16'd4121;
      114491:data<=-16'd3974;
      114492:data<=-16'd3187;
      114493:data<=-16'd3027;
      114494:data<=-16'd2984;
      114495:data<=-16'd2629;
      114496:data<=-16'd2974;
      114497:data<=-16'd3802;
      114498:data<=-16'd4030;
      114499:data<=-16'd3815;
      114500:data<=-16'd3632;
      114501:data<=-16'd3157;
      114502:data<=-16'd2596;
      114503:data<=-16'd2499;
      114504:data<=-16'd2252;
      114505:data<=-16'd1632;
      114506:data<=-16'd1495;
      114507:data<=-16'd1579;
      114508:data<=-16'd1237;
      114509:data<=-16'd1275;
      114510:data<=-16'd2182;
      114511:data<=-16'd2799;
      114512:data<=-16'd2441;
      114513:data<=-16'd2011;
      114514:data<=-16'd1970;
      114515:data<=-16'd1721;
      114516:data<=-16'd1236;
      114517:data<=-16'd939;
      114518:data<=-16'd699;
      114519:data<=-16'd440;
      114520:data<=-16'd397;
      114521:data<=-16'd115;
      114522:data<=16'd623;
      114523:data<=16'd202;
      114524:data<=-16'd1500;
      114525:data<=-16'd1750;
      114526:data<=-16'd883;
      114527:data<=-16'd1005;
      114528:data<=-16'd315;
      114529:data<=16'd1616;
      114530:data<=16'd2215;
      114531:data<=16'd2273;
      114532:data<=16'd2828;
      114533:data<=16'd2579;
      114534:data<=16'd2472;
      114535:data<=16'd3116;
      114536:data<=16'd2519;
      114537:data<=16'd955;
      114538:data<=16'd511;
      114539:data<=16'd990;
      114540:data<=16'd1309;
      114541:data<=16'd1595;
      114542:data<=16'd1833;
      114543:data<=16'd1770;
      114544:data<=16'd2070;
      114545:data<=16'd2631;
      114546:data<=16'd2554;
      114547:data<=16'd2385;
      114548:data<=16'd2564;
      114549:data<=16'd2258;
      114550:data<=16'd1292;
      114551:data<=16'd505;
      114552:data<=16'd651;
      114553:data<=16'd1118;
      114554:data<=16'd1022;
      114555:data<=16'd1231;
      114556:data<=16'd1745;
      114557:data<=16'd1489;
      114558:data<=16'd1483;
      114559:data<=16'd2140;
      114560:data<=16'd2315;
      114561:data<=16'd2420;
      114562:data<=16'd2379;
      114563:data<=16'd1348;
      114564:data<=16'd628;
      114565:data<=16'd975;
      114566:data<=16'd1061;
      114567:data<=16'd826;
      114568:data<=16'd1145;
      114569:data<=16'd1569;
      114570:data<=16'd1709;
      114571:data<=16'd1944;
      114572:data<=16'd2114;
      114573:data<=16'd2134;
      114574:data<=16'd2256;
      114575:data<=16'd2188;
      114576:data<=16'd2161;
      114577:data<=16'd2558;
      114578:data<=16'd2648;
      114579:data<=16'd2587;
      114580:data<=16'd2984;
      114581:data<=16'd2499;
      114582:data<=16'd999;
      114583:data<=16'd787;
      114584:data<=16'd1510;
      114585:data<=16'd1283;
      114586:data<=16'd1162;
      114587:data<=16'd1629;
      114588:data<=16'd1639;
      114589:data<=16'd2438;
      114590:data<=16'd4002;
      114591:data<=16'd4108;
      114592:data<=16'd3647;
      114593:data<=16'd4026;
      114594:data<=16'd4249;
      114595:data<=16'd4064;
      114596:data<=16'd3988;
      114597:data<=16'd4178;
      114598:data<=16'd4376;
      114599:data<=16'd4140;
      114600:data<=16'd3983;
      114601:data<=16'd4049;
      114602:data<=16'd4272;
      114603:data<=16'd5465;
      114604:data<=16'd6581;
      114605:data<=16'd6391;
      114606:data<=16'd6197;
      114607:data<=16'd6451;
      114608:data<=16'd6344;
      114609:data<=16'd5962;
      114610:data<=16'd5817;
      114611:data<=16'd5967;
      114612:data<=16'd5873;
      114613:data<=16'd5717;
      114614:data<=16'd5727;
      114615:data<=16'd5526;
      114616:data<=16'd6143;
      114617:data<=16'd7498;
      114618:data<=16'd7686;
      114619:data<=16'd7282;
      114620:data<=16'd7201;
      114621:data<=16'd6927;
      114622:data<=16'd6717;
      114623:data<=16'd6438;
      114624:data<=16'd6073;
      114625:data<=16'd6276;
      114626:data<=16'd6516;
      114627:data<=16'd6187;
      114628:data<=16'd5691;
      114629:data<=16'd6037;
      114630:data<=16'd7348;
      114631:data<=16'd7923;
      114632:data<=16'd7394;
      114633:data<=16'd7054;
      114634:data<=16'd7447;
      114635:data<=16'd8511;
      114636:data<=16'd9062;
      114637:data<=16'd8616;
      114638:data<=16'd8407;
      114639:data<=16'd8240;
      114640:data<=16'd7761;
      114641:data<=16'd7527;
      114642:data<=16'd7641;
      114643:data<=16'd8495;
      114644:data<=16'd9104;
      114645:data<=16'd8490;
      114646:data<=16'd8219;
      114647:data<=16'd8193;
      114648:data<=16'd7506;
      114649:data<=16'd7279;
      114650:data<=16'd7233;
      114651:data<=16'd6766;
      114652:data<=16'd6673;
      114653:data<=16'd6525;
      114654:data<=16'd5815;
      114655:data<=16'd5721;
      114656:data<=16'd6878;
      114657:data<=16'd7688;
      114658:data<=16'd7013;
      114659:data<=16'd6358;
      114660:data<=16'd6479;
      114661:data<=16'd6414;
      114662:data<=16'd6058;
      114663:data<=16'd5609;
      114664:data<=16'd5190;
      114665:data<=16'd5043;
      114666:data<=16'd4921;
      114667:data<=16'd4485;
      114668:data<=16'd3897;
      114669:data<=16'd4356;
      114670:data<=16'd5779;
      114671:data<=16'd5858;
      114672:data<=16'd4913;
      114673:data<=16'd4801;
      114674:data<=16'd4836;
      114675:data<=16'd4523;
      114676:data<=16'd4234;
      114677:data<=16'd3817;
      114678:data<=16'd3527;
      114679:data<=16'd3582;
      114680:data<=16'd3595;
      114681:data<=16'd3021;
      114682:data<=16'd2939;
      114683:data<=16'd4437;
      114684:data<=16'd5095;
      114685:data<=16'd4320;
      114686:data<=16'd4326;
      114687:data<=16'd3745;
      114688:data<=16'd2024;
      114689:data<=16'd1260;
      114690:data<=16'd899;
      114691:data<=16'd479;
      114692:data<=16'd502;
      114693:data<=16'd376;
      114694:data<=16'd246;
      114695:data<=16'd535;
      114696:data<=16'd1339;
      114697:data<=16'd2011;
      114698:data<=16'd1739;
      114699:data<=16'd1538;
      114700:data<=16'd1454;
      114701:data<=16'd913;
      114702:data<=16'd920;
      114703:data<=16'd945;
      114704:data<=16'd576;
      114705:data<=16'd578;
      114706:data<=16'd297;
      114707:data<=16'd0;
      114708:data<=16'd265;
      114709:data<=16'd836;
      114710:data<=16'd1782;
      114711:data<=16'd1800;
      114712:data<=16'd1084;
      114713:data<=16'd1313;
      114714:data<=16'd1155;
      114715:data<=16'd462;
      114716:data<=16'd491;
      114717:data<=16'd276;
      114718:data<=16'd133;
      114719:data<=16'd440;
      114720:data<=-16'd168;
      114721:data<=-16'd869;
      114722:data<=-16'd5;
      114723:data<=16'd1556;
      114724:data<=16'd1809;
      114725:data<=16'd955;
      114726:data<=16'd785;
      114727:data<=16'd916;
      114728:data<=16'd558;
      114729:data<=16'd162;
      114730:data<=-16'd506;
      114731:data<=-16'd848;
      114732:data<=-16'd297;
      114733:data<=-16'd281;
      114734:data<=-16'd925;
      114735:data<=-16'd687;
      114736:data<=16'd604;
      114737:data<=16'd1474;
      114738:data<=16'd1119;
      114739:data<=16'd473;
      114740:data<=16'd352;
      114741:data<=16'd1146;
      114742:data<=16'd2320;
      114743:data<=16'd2068;
      114744:data<=16'd1136;
      114745:data<=16'd1271;
      114746:data<=16'd1333;
      114747:data<=16'd798;
      114748:data<=16'd790;
      114749:data<=16'd1557;
      114750:data<=16'd2353;
      114751:data<=16'd2334;
      114752:data<=16'd2067;
      114753:data<=16'd1889;
      114754:data<=16'd1190;
      114755:data<=16'd769;
      114756:data<=16'd660;
      114757:data<=16'd155;
      114758:data<=16'd18;
      114759:data<=16'd20;
      114760:data<=-16'd334;
      114761:data<=-16'd321;
      114762:data<=16'd249;
      114763:data<=16'd951;
      114764:data<=16'd981;
      114765:data<=16'd673;
      114766:data<=16'd776;
      114767:data<=16'd281;
      114768:data<=-16'd485;
      114769:data<=-16'd566;
      114770:data<=-16'd842;
      114771:data<=-16'd1051;
      114772:data<=-16'd948;
      114773:data<=-16'd1345;
      114774:data<=-16'd1747;
      114775:data<=-16'd1253;
      114776:data<=16'd82;
      114777:data<=16'd482;
      114778:data<=-16'd519;
      114779:data<=-16'd594;
      114780:data<=-16'd346;
      114781:data<=-16'd946;
      114782:data<=-16'd1005;
      114783:data<=-16'd1295;
      114784:data<=-16'd1895;
      114785:data<=-16'd1639;
      114786:data<=-16'd1848;
      114787:data<=-16'd2397;
      114788:data<=-16'd2491;
      114789:data<=-16'd2590;
      114790:data<=-16'd2411;
      114791:data<=-16'd2684;
      114792:data<=-16'd3209;
      114793:data<=-16'd3045;
      114794:data<=-16'd3785;
      114795:data<=-16'd5342;
      114796:data<=-16'd6034;
      114797:data<=-16'd5981;
      114798:data<=-16'd5812;
      114799:data<=-16'd5970;
      114800:data<=-16'd5723;
      114801:data<=-16'd5495;
      114802:data<=-16'd6942;
      114803:data<=-16'd8026;
      114804:data<=-16'd7591;
      114805:data<=-16'd7521;
      114806:data<=-16'd7586;
      114807:data<=-16'd7514;
      114808:data<=-16'd7491;
      114809:data<=-16'd7245;
      114810:data<=-16'd7413;
      114811:data<=-16'd7460;
      114812:data<=-16'd7319;
      114813:data<=-16'd7272;
      114814:data<=-16'd6654;
      114815:data<=-16'd7418;
      114816:data<=-16'd9306;
      114817:data<=-16'd9163;
      114818:data<=-16'd8505;
      114819:data<=-16'd8645;
      114820:data<=-16'd8351;
      114821:data<=-16'd8252;
      114822:data<=-16'd8254;
      114823:data<=-16'd7871;
      114824:data<=-16'd7524;
      114825:data<=-16'd7291;
      114826:data<=-16'd7363;
      114827:data<=-16'd7150;
      114828:data<=-16'd7224;
      114829:data<=-16'd8563;
      114830:data<=-16'd9110;
      114831:data<=-16'd8573;
      114832:data<=-16'd8508;
      114833:data<=-16'd8301;
      114834:data<=-16'd8041;
      114835:data<=-16'd8105;
      114836:data<=-16'd7959;
      114837:data<=-16'd7726;
      114838:data<=-16'd7373;
      114839:data<=-16'd7127;
      114840:data<=-16'd7060;
      114841:data<=-16'd7166;
      114842:data<=-16'd8093;
      114843:data<=-16'd8546;
      114844:data<=-16'd7802;
      114845:data<=-16'd7827;
      114846:data<=-16'd8191;
      114847:data<=-16'd6919;
      114848:data<=-16'd4978;
      114849:data<=-16'd4498;
      114850:data<=-16'd5090;
      114851:data<=-16'd4984;
      114852:data<=-16'd4531;
      114853:data<=-16'd4302;
      114854:data<=-16'd4272;
      114855:data<=-16'd5360;
      114856:data<=-16'd6208;
      114857:data<=-16'd5656;
      114858:data<=-16'd5641;
      114859:data<=-16'd5962;
      114860:data<=-16'd5618;
      114861:data<=-16'd5325;
      114862:data<=-16'd5174;
      114863:data<=-16'd5204;
      114864:data<=-16'd4940;
      114865:data<=-16'd4478;
      114866:data<=-16'd4510;
      114867:data<=-16'd3959;
      114868:data<=-16'd4026;
      114869:data<=-16'd5745;
      114870:data<=-16'd6076;
      114871:data<=-16'd5213;
      114872:data<=-16'd5110;
      114873:data<=-16'd4975;
      114874:data<=-16'd4951;
      114875:data<=-16'd4861;
      114876:data<=-16'd4320;
      114877:data<=-16'd4172;
      114878:data<=-16'd4147;
      114879:data<=-16'd4003;
      114880:data<=-16'd3627;
      114881:data<=-16'd3548;
      114882:data<=-16'd4890;
      114883:data<=-16'd5709;
      114884:data<=-16'd5125;
      114885:data<=-16'd4931;
      114886:data<=-16'd4575;
      114887:data<=-16'd3971;
      114888:data<=-16'd3956;
      114889:data<=-16'd3703;
      114890:data<=-16'd3189;
      114891:data<=-16'd2983;
      114892:data<=-16'd3018;
      114893:data<=-16'd2701;
      114894:data<=-16'd2587;
      114895:data<=-16'd4087;
      114896:data<=-16'd4992;
      114897:data<=-16'd4284;
      114898:data<=-16'd4375;
      114899:data<=-16'd4143;
      114900:data<=-16'd3844;
      114901:data<=-16'd5363;
      114902:data<=-16'd5833;
      114903:data<=-16'd5042;
      114904:data<=-16'd4948;
      114905:data<=-16'd4410;
      114906:data<=-16'd3953;
      114907:data<=-16'd4027;
      114908:data<=-16'd4217;
      114909:data<=-16'd5065;
      114910:data<=-16'd5181;
      114911:data<=-16'd4578;
      114912:data<=-16'd4534;
      114913:data<=-16'd4126;
      114914:data<=-16'd3554;
      114915:data<=-16'd3280;
      114916:data<=-16'd2954;
      114917:data<=-16'd2919;
      114918:data<=-16'd2784;
      114919:data<=-16'd2353;
      114920:data<=-16'd1750;
      114921:data<=-16'd1821;
      114922:data<=-16'd3469;
      114923:data<=-16'd4081;
      114924:data<=-16'd3021;
      114925:data<=-16'd2961;
      114926:data<=-16'd2889;
      114927:data<=-16'd2255;
      114928:data<=-16'd2188;
      114929:data<=-16'd1613;
      114930:data<=-16'd1158;
      114931:data<=-16'd1535;
      114932:data<=-16'd1216;
      114933:data<=-16'd502;
      114934:data<=-16'd746;
      114935:data<=-16'd1844;
      114936:data<=-16'd2314;
      114937:data<=-16'd1770;
      114938:data<=-16'd1524;
      114939:data<=-16'd1187;
      114940:data<=-16'd655;
      114941:data<=-16'd883;
      114942:data<=-16'd792;
      114943:data<=-16'd318;
      114944:data<=-16'd246;
      114945:data<=-16'd11;
      114946:data<=16'd100;
      114947:data<=16'd5;
      114948:data<=-16'd459;
      114949:data<=-16'd1444;
      114950:data<=-16'd1353;
      114951:data<=-16'd714;
      114952:data<=-16'd707;
      114953:data<=16'd211;
      114954:data<=16'd1707;
      114955:data<=16'd2279;
      114956:data<=16'd2488;
      114957:data<=16'd2693;
      114958:data<=16'd2675;
      114959:data<=16'd2877;
      114960:data<=16'd3324;
      114961:data<=16'd2596;
      114962:data<=16'd1049;
      114963:data<=16'd1171;
      114964:data<=16'd1879;
      114965:data<=16'd1503;
      114966:data<=16'd1674;
      114967:data<=16'd2205;
      114968:data<=16'd2203;
      114969:data<=16'd2332;
      114970:data<=16'd2224;
      114971:data<=16'd2126;
      114972:data<=16'd2657;
      114973:data<=16'd3107;
      114974:data<=16'd2500;
      114975:data<=16'd931;
      114976:data<=16'd587;
      114977:data<=16'd1438;
      114978:data<=16'd1243;
      114979:data<=16'd1192;
      114980:data<=16'd1800;
      114981:data<=16'd1842;
      114982:data<=16'd2261;
      114983:data<=16'd2635;
      114984:data<=16'd2249;
      114985:data<=16'd2265;
      114986:data<=16'd2646;
      114987:data<=16'd2575;
      114988:data<=16'd1445;
      114989:data<=16'd406;
      114990:data<=16'd875;
      114991:data<=16'd1122;
      114992:data<=16'd1016;
      114993:data<=16'd1612;
      114994:data<=16'd1750;
      114995:data<=16'd2012;
      114996:data<=16'd2499;
      114997:data<=16'd2234;
      114998:data<=16'd2355;
      114999:data<=16'd2522;
      115000:data<=16'd2496;
      115001:data<=16'd3046;
      115002:data<=16'd3021;
      115003:data<=16'd2795;
      115004:data<=16'd3024;
      115005:data<=16'd3098;
      115006:data<=16'd3145;
      115007:data<=16'd2209;
      115008:data<=16'd1074;
      115009:data<=16'd1401;
      115010:data<=16'd1674;
      115011:data<=16'd1911;
      115012:data<=16'd2353;
      115013:data<=16'd2021;
      115014:data<=16'd2736;
      115015:data<=16'd4319;
      115016:data<=16'd4645;
      115017:data<=16'd4382;
      115018:data<=16'd4250;
      115019:data<=16'd4449;
      115020:data<=16'd4720;
      115021:data<=16'd4511;
      115022:data<=16'd4484;
      115023:data<=16'd4573;
      115024:data<=16'd4781;
      115025:data<=16'd4918;
      115026:data<=16'd4181;
      115027:data<=16'd4620;
      115028:data<=16'd6517;
      115029:data<=16'd7043;
      115030:data<=16'd6733;
      115031:data<=16'd6768;
      115032:data<=16'd6654;
      115033:data<=16'd6399;
      115034:data<=16'd6187;
      115035:data<=16'd6363;
      115036:data<=16'd6243;
      115037:data<=16'd5817;
      115038:data<=16'd6059;
      115039:data<=16'd5767;
      115040:data<=16'd5726;
      115041:data<=16'd7292;
      115042:data<=16'd7978;
      115043:data<=16'd7720;
      115044:data<=16'd7785;
      115045:data<=16'd7371;
      115046:data<=16'd7089;
      115047:data<=16'd6915;
      115048:data<=16'd6583;
      115049:data<=16'd6714;
      115050:data<=16'd6522;
      115051:data<=16'd6222;
      115052:data<=16'd5967;
      115053:data<=16'd5689;
      115054:data<=16'd6951;
      115055:data<=16'd8132;
      115056:data<=16'd7680;
      115057:data<=16'd7611;
      115058:data<=16'd7592;
      115059:data<=16'd7219;
      115060:data<=16'd7882;
      115061:data<=16'd8810;
      115062:data<=16'd8883;
      115063:data<=16'd8357;
      115064:data<=16'd8072;
      115065:data<=16'd7867;
      115066:data<=16'd7195;
      115067:data<=16'd7738;
      115068:data<=16'd9191;
      115069:data<=16'd9142;
      115070:data<=16'd8569;
      115071:data<=16'd8392;
      115072:data<=16'd7917;
      115073:data<=16'd7579;
      115074:data<=16'd7388;
      115075:data<=16'd6990;
      115076:data<=16'd6589;
      115077:data<=16'd6645;
      115078:data<=16'd6728;
      115079:data<=16'd5949;
      115080:data<=16'd5918;
      115081:data<=16'd7060;
      115082:data<=16'd7295;
      115083:data<=16'd7160;
      115084:data<=16'd6954;
      115085:data<=16'd6252;
      115086:data<=16'd6252;
      115087:data<=16'd6128;
      115088:data<=16'd5517;
      115089:data<=16'd5442;
      115090:data<=16'd5171;
      115091:data<=16'd4915;
      115092:data<=16'd4687;
      115093:data<=16'd4396;
      115094:data<=16'd5288;
      115095:data<=16'd5812;
      115096:data<=16'd5336;
      115097:data<=16'd5500;
      115098:data<=16'd5125;
      115099:data<=16'd4258;
      115100:data<=16'd4320;
      115101:data<=16'd4413;
      115102:data<=16'd4181;
      115103:data<=16'd3888;
      115104:data<=16'd3679;
      115105:data<=16'd3385;
      115106:data<=16'd2872;
      115107:data<=16'd3707;
      115108:data<=16'd5168;
      115109:data<=16'd4998;
      115110:data<=16'd4293;
      115111:data<=16'd4131;
      115112:data<=16'd4088;
      115113:data<=16'd3372;
      115114:data<=16'd1814;
      115115:data<=16'd1265;
      115116:data<=16'd1418;
      115117:data<=16'd1057;
      115118:data<=16'd1033;
      115119:data<=16'd741;
      115120:data<=16'd1022;
      115121:data<=16'd2708;
      115122:data<=16'd2805;
      115123:data<=16'd1938;
      115124:data<=16'd2205;
      115125:data<=16'd2093;
      115126:data<=16'd1829;
      115127:data<=16'd1856;
      115128:data<=16'd1404;
      115129:data<=16'd1243;
      115130:data<=16'd1424;
      115131:data<=16'd1225;
      115132:data<=16'd667;
      115133:data<=16'd869;
      115134:data<=16'd2347;
      115135:data<=16'd2946;
      115136:data<=16'd2447;
      115137:data<=16'd2397;
      115138:data<=16'd2085;
      115139:data<=16'd1757;
      115140:data<=16'd1801;
      115141:data<=16'd1404;
      115142:data<=16'd1157;
      115143:data<=16'd1145;
      115144:data<=16'd1089;
      115145:data<=16'd999;
      115146:data<=16'd804;
      115147:data<=16'd1639;
      115148:data<=16'd2641;
      115149:data<=16'd2391;
      115150:data<=16'd2275;
      115151:data<=16'd2193;
      115152:data<=16'd1671;
      115153:data<=16'd1497;
      115154:data<=16'd1259;
      115155:data<=16'd1008;
      115156:data<=16'd713;
      115157:data<=16'd441;
      115158:data<=16'd640;
      115159:data<=16'd211;
      115160:data<=16'd379;
      115161:data<=16'd1932;
      115162:data<=16'd2036;
      115163:data<=16'd1585;
      115164:data<=16'd1754;
      115165:data<=16'd964;
      115166:data<=16'd1017;
      115167:data<=16'd2306;
      115168:data<=16'd2393;
      115169:data<=16'd1933;
      115170:data<=16'd1859;
      115171:data<=16'd1515;
      115172:data<=16'd974;
      115173:data<=16'd1381;
      115174:data<=16'd2643;
      115175:data<=16'd2834;
      115176:data<=16'd2472;
      115177:data<=16'd2579;
      115178:data<=16'd1996;
      115179:data<=16'd1328;
      115180:data<=16'd1108;
      115181:data<=16'd804;
      115182:data<=16'd843;
      115183:data<=16'd619;
      115184:data<=16'd223;
      115185:data<=-16'd3;
      115186:data<=-16'd365;
      115187:data<=16'd637;
      115188:data<=16'd1736;
      115189:data<=16'd1052;
      115190:data<=16'd808;
      115191:data<=16'd719;
      115192:data<=-16'd76;
      115193:data<=-16'd36;
      115194:data<=-16'd45;
      115195:data<=-16'd423;
      115196:data<=-16'd513;
      115197:data<=-16'd916;
      115198:data<=-16'd1110;
      115199:data<=-16'd1055;
      115200:data<=-16'd755;
      115201:data<=-16'd68;
      115202:data<=-16'd206;
      115203:data<=-16'd506;
      115204:data<=-16'd494;
      115205:data<=-16'd963;
      115206:data<=-16'd936;
      115207:data<=-16'd776;
      115208:data<=-16'd1201;
      115209:data<=-16'd1478;
      115210:data<=-16'd1973;
      115211:data<=-16'd2202;
      115212:data<=-16'd1962;
      115213:data<=-16'd2202;
      115214:data<=-16'd2375;
      115215:data<=-16'd2640;
      115216:data<=-16'd3018;
      115217:data<=-16'd2717;
      115218:data<=-16'd2796;
      115219:data<=-16'd3741;
      115220:data<=-16'd4916;
      115221:data<=-16'd5529;
      115222:data<=-16'd5203;
      115223:data<=-16'd5385;
      115224:data<=-16'd5727;
      115225:data<=-16'd5386;
      115226:data<=-16'd5984;
      115227:data<=-16'd7100;
      115228:data<=-16'd7750;
      115229:data<=-16'd8070;
      115230:data<=-16'd7603;
      115231:data<=-16'd7488;
      115232:data<=-16'd7746;
      115233:data<=-16'd7362;
      115234:data<=-16'd7326;
      115235:data<=-16'd7235;
      115236:data<=-16'd7071;
      115237:data<=-16'd7359;
      115238:data<=-16'd6910;
      115239:data<=-16'd7103;
      115240:data<=-16'd8375;
      115241:data<=-16'd8671;
      115242:data<=-16'd8739;
      115243:data<=-16'd8636;
      115244:data<=-16'd8155;
      115245:data<=-16'd8355;
      115246:data<=-16'd8019;
      115247:data<=-16'd7498;
      115248:data<=-16'd7746;
      115249:data<=-16'd7504;
      115250:data<=-16'd7377;
      115251:data<=-16'd7330;
      115252:data<=-16'd6943;
      115253:data<=-16'd7859;
      115254:data<=-16'd9077;
      115255:data<=-16'd9041;
      115256:data<=-16'd8702;
      115257:data<=-16'd8564;
      115258:data<=-16'd8498;
      115259:data<=-16'd8146;
      115260:data<=-16'd7770;
      115261:data<=-16'd7756;
      115262:data<=-16'd7555;
      115263:data<=-16'd7621;
      115264:data<=-16'd7615;
      115265:data<=-16'd6984;
      115266:data<=-16'd7573;
      115267:data<=-16'd9018;
      115268:data<=-16'd9277;
      115269:data<=-16'd8560;
      115270:data<=-16'd7858;
      115271:data<=-16'd7884;
      115272:data<=-16'd7498;
      115273:data<=-16'd5961;
      115274:data<=-16'd5125;
      115275:data<=-16'd4971;
      115276:data<=-16'd4975;
      115277:data<=-16'd5245;
      115278:data<=-16'd4628;
      115279:data<=-16'd4658;
      115280:data<=-16'd6181;
      115281:data<=-16'd6643;
      115282:data<=-16'd6261;
      115283:data<=-16'd5915;
      115284:data<=-16'd5366;
      115285:data<=-16'd5451;
      115286:data<=-16'd5586;
      115287:data<=-16'd5190;
      115288:data<=-16'd4767;
      115289:data<=-16'd4413;
      115290:data<=-16'd4508;
      115291:data<=-16'd4373;
      115292:data<=-16'd4215;
      115293:data<=-16'd5392;
      115294:data<=-16'd6252;
      115295:data<=-16'd5909;
      115296:data<=-16'd5752;
      115297:data<=-16'd5635;
      115298:data<=-16'd5485;
      115299:data<=-16'd5483;
      115300:data<=-16'd5301;
      115301:data<=-16'd4942;
      115302:data<=-16'd4416;
      115303:data<=-16'd4491;
      115304:data<=-16'd4742;
      115305:data<=-16'd4131;
      115306:data<=-16'd4476;
      115307:data<=-16'd5841;
      115308:data<=-16'd5941;
      115309:data<=-16'd5515;
      115310:data<=-16'd5611;
      115311:data<=-16'd5495;
      115312:data<=-16'd5016;
      115313:data<=-16'd4446;
      115314:data<=-16'd3961;
      115315:data<=-16'd3768;
      115316:data<=-16'd4109;
      115317:data<=-16'd4158;
      115318:data<=-16'd3247;
      115319:data<=-16'd3542;
      115320:data<=-16'd5350;
      115321:data<=-16'd5758;
      115322:data<=-16'd5204;
      115323:data<=-16'd5357;
      115324:data<=-16'd5222;
      115325:data<=-16'd4928;
      115326:data<=-16'd5520;
      115327:data<=-16'd5990;
      115328:data<=-16'd5644;
      115329:data<=-16'd5673;
      115330:data<=-16'd5771;
      115331:data<=-16'd4889;
      115332:data<=-16'd4864;
      115333:data<=-16'd6205;
      115334:data<=-16'd6590;
      115335:data<=-16'd6199;
      115336:data<=-16'd5841;
      115337:data<=-16'd5177;
      115338:data<=-16'd4911;
      115339:data<=-16'd4868;
      115340:data<=-16'd4457;
      115341:data<=-16'd4026;
      115342:data<=-16'd3677;
      115343:data<=-16'd3736;
      115344:data<=-16'd3644;
      115345:data<=-16'd3159;
      115346:data<=-16'd3761;
      115347:data<=-16'd4699;
      115348:data<=-16'd4534;
      115349:data<=-16'd4034;
      115350:data<=-16'd3509;
      115351:data<=-16'd3122;
      115352:data<=-16'd3084;
      115353:data<=-16'd2852;
      115354:data<=-16'd2464;
      115355:data<=-16'd2008;
      115356:data<=-16'd1753;
      115357:data<=-16'd1650;
      115358:data<=-16'd993;
      115359:data<=-16'd1133;
      115360:data<=-16'd2469;
      115361:data<=-16'd2693;
      115362:data<=-16'd2100;
      115363:data<=-16'd2093;
      115364:data<=-16'd1867;
      115365:data<=-16'd1178;
      115366:data<=-16'd758;
      115367:data<=-16'd672;
      115368:data<=-16'd534;
      115369:data<=-16'd399;
      115370:data<=-16'd262;
      115371:data<=16'd191;
      115372:data<=-16'd106;
      115373:data<=-16'd1350;
      115374:data<=-16'd1548;
      115375:data<=-16'd916;
      115376:data<=-16'd631;
      115377:data<=-16'd397;
      115378:data<=-16'd291;
      115379:data<=16'd555;
      115380:data<=16'd2390;
      115381:data<=16'd3093;
      115382:data<=16'd2670;
      115383:data<=16'd2666;
      115384:data<=16'd3022;
      115385:data<=16'd3015;
      115386:data<=16'd2012;
      115387:data<=16'd1092;
      115388:data<=16'd1515;
      115389:data<=16'd1929;
      115390:data<=16'd1889;
      115391:data<=16'd2334;
      115392:data<=16'd2508;
      115393:data<=16'd2315;
      115394:data<=16'd2663;
      115395:data<=16'd2880;
      115396:data<=16'd2605;
      115397:data<=16'd2949;
      115398:data<=16'd3551;
      115399:data<=16'd2742;
      115400:data<=16'd1227;
      115401:data<=16'd967;
      115402:data<=16'd1533;
      115403:data<=16'd1703;
      115404:data<=16'd1741;
      115405:data<=16'd2033;
      115406:data<=16'd2259;
      115407:data<=16'd2223;
      115408:data<=16'd2312;
      115409:data<=16'd2570;
      115410:data<=16'd2634;
      115411:data<=16'd2696;
      115412:data<=16'd2382;
      115413:data<=16'd1187;
      115414:data<=16'd570;
      115415:data<=16'd1219;
      115416:data<=16'd1648;
      115417:data<=16'd1682;
      115418:data<=16'd1859;
      115419:data<=16'd1545;
      115420:data<=16'd1195;
      115421:data<=16'd1760;
      115422:data<=16'd2325;
      115423:data<=16'd2413;
      115424:data<=16'd2760;
      115425:data<=16'd2990;
      115426:data<=16'd2914;
      115427:data<=16'd3266;
      115428:data<=16'd3591;
      115429:data<=16'd3448;
      115430:data<=16'd3338;
      115431:data<=16'd3087;
      115432:data<=16'd2790;
      115433:data<=16'd3071;
      115434:data<=16'd3530;
      115435:data<=16'd3683;
      115436:data<=16'd3732;
      115437:data<=16'd3900;
      115438:data<=16'd4487;
      115439:data<=16'd5401;
      115440:data<=16'd5893;
      115441:data<=16'd5897;
      115442:data<=16'd5958;
      115443:data<=16'd5829;
      115444:data<=16'd5398;
      115445:data<=16'd5272;
      115446:data<=16'd5382;
      115447:data<=16'd5535;
      115448:data<=16'd5682;
      115449:data<=16'd5448;
      115450:data<=16'd5421;
      115451:data<=16'd5862;
      115452:data<=16'd6260;
      115453:data<=16'd7145;
      115454:data<=16'd7652;
      115455:data<=16'd6872;
      115456:data<=16'd6936;
      115457:data<=16'd7595;
      115458:data<=16'd6887;
      115459:data<=16'd6338;
      115460:data<=16'd6570;
      115461:data<=16'd6361;
      115462:data<=16'd6153;
      115463:data<=16'd6044;
      115464:data<=16'd5953;
      115465:data<=16'd6721;
      115466:data<=16'd7914;
      115467:data<=16'd8184;
      115468:data<=16'd7389;
      115469:data<=16'd6899;
      115470:data<=16'd7259;
      115471:data<=16'd7365;
      115472:data<=16'd7122;
      115473:data<=16'd6907;
      115474:data<=16'd6475;
      115475:data<=16'd6388;
      115476:data<=16'd6625;
      115477:data<=16'd6413;
      115478:data<=16'd6311;
      115479:data<=16'd6978;
      115480:data<=16'd7749;
      115481:data<=16'd7662;
      115482:data<=16'd7181;
      115483:data<=16'd7230;
      115484:data<=16'd7077;
      115485:data<=16'd6620;
      115486:data<=16'd6631;
      115487:data<=16'd6240;
      115488:data<=16'd5604;
      115489:data<=16'd5786;
      115490:data<=16'd5968;
      115491:data<=16'd6082;
      115492:data<=16'd6769;
      115493:data<=16'd7262;
      115494:data<=16'd7059;
      115495:data<=16'd6531;
      115496:data<=16'd6404;
      115497:data<=16'd6669;
      115498:data<=16'd6355;
      115499:data<=16'd5921;
      115500:data<=16'd5853;
      115501:data<=16'd5524;
      115502:data<=16'd5697;
      115503:data<=16'd6088;
      115504:data<=16'd5333;
      115505:data<=16'd5183;
      115506:data<=16'd6432;
      115507:data<=16'd6675;
      115508:data<=16'd5967;
      115509:data<=16'd5782;
      115510:data<=16'd5491;
      115511:data<=16'd4908;
      115512:data<=16'd4915;
      115513:data<=16'd5309;
      115514:data<=16'd5198;
      115515:data<=16'd4549;
      115516:data<=16'd4058;
      115517:data<=16'd3836;
      115518:data<=16'd4132;
      115519:data<=16'd5328;
      115520:data<=16'd5868;
      115521:data<=16'd5043;
      115522:data<=16'd4790;
      115523:data<=16'd5127;
      115524:data<=16'd4833;
      115525:data<=16'd4322;
      115526:data<=16'd3782;
      115527:data<=16'd3571;
      115528:data<=16'd3786;
      115529:data<=16'd3365;
      115530:data<=16'd3137;
      115531:data<=16'd3899;
      115532:data<=16'd4513;
      115533:data<=16'd5021;
      115534:data<=16'd5112;
      115535:data<=16'd4346;
      115536:data<=16'd4159;
      115537:data<=16'd4262;
      115538:data<=16'd3803;
      115539:data<=16'd3510;
      115540:data<=16'd2955;
      115541:data<=16'd2475;
      115542:data<=16'd2995;
      115543:data<=16'd3065;
      115544:data<=16'd2648;
      115545:data<=16'd3316;
      115546:data<=16'd4299;
      115547:data<=16'd4347;
      115548:data<=16'd3798;
      115549:data<=16'd3495;
      115550:data<=16'd3422;
      115551:data<=16'd2995;
      115552:data<=16'd2751;
      115553:data<=16'd2863;
      115554:data<=16'd2294;
      115555:data<=16'd1522;
      115556:data<=16'd1450;
      115557:data<=16'd1553;
      115558:data<=16'd2024;
      115559:data<=16'd3037;
      115560:data<=16'd3112;
      115561:data<=16'd2229;
      115562:data<=16'd2006;
      115563:data<=16'd2030;
      115564:data<=16'd1639;
      115565:data<=16'd1712;
      115566:data<=16'd1629;
      115567:data<=16'd1081;
      115568:data<=16'd1472;
      115569:data<=16'd1524;
      115570:data<=16'd449;
      115571:data<=16'd1052;
      115572:data<=16'd2602;
      115573:data<=16'd2226;
      115574:data<=16'd1480;
      115575:data<=16'd1613;
      115576:data<=16'd1547;
      115577:data<=16'd1532;
      115578:data<=16'd1343;
      115579:data<=16'd587;
      115580:data<=16'd403;
      115581:data<=16'd528;
      115582:data<=16'd102;
      115583:data<=-16'd294;
      115584:data<=-16'd212;
      115585:data<=16'd696;
      115586:data<=16'd1770;
      115587:data<=16'd1598;
      115588:data<=16'd1190;
      115589:data<=16'd1277;
      115590:data<=16'd843;
      115591:data<=16'd696;
      115592:data<=16'd817;
      115593:data<=-16'd42;
      115594:data<=-16'd476;
      115595:data<=-16'd246;
      115596:data<=-16'd622;
      115597:data<=-16'd356;
      115598:data<=16'd434;
      115599:data<=16'd296;
      115600:data<=16'd346;
      115601:data<=16'd658;
      115602:data<=16'd218;
      115603:data<=16'd74;
      115604:data<=16'd343;
      115605:data<=16'd182;
      115606:data<=-16'd146;
      115607:data<=-16'd895;
      115608:data<=-16'd1548;
      115609:data<=-16'd1154;
      115610:data<=-16'd1230;
      115611:data<=-16'd1603;
      115612:data<=-16'd190;
      115613:data<=16'd1025;
      115614:data<=16'd523;
      115615:data<=16'd475;
      115616:data<=16'd497;
      115617:data<=-16'd262;
      115618:data<=-16'd243;
      115619:data<=-16'd152;
      115620:data<=-16'd887;
      115621:data<=-16'd1207;
      115622:data<=-16'd1316;
      115623:data<=-16'd1513;
      115624:data<=-16'd1066;
      115625:data<=-16'd491;
      115626:data<=-16'd334;
      115627:data<=-16'd372;
      115628:data<=-16'd459;
      115629:data<=-16'd406;
      115630:data<=-16'd564;
      115631:data<=-16'd1107;
      115632:data<=-16'd1246;
      115633:data<=-16'd1165;
      115634:data<=-16'd1641;
      115635:data<=-16'd2087;
      115636:data<=-16'd2206;
      115637:data<=-16'd2526;
      115638:data<=-16'd2591;
      115639:data<=-16'd2493;
      115640:data<=-16'd2881;
      115641:data<=-16'd2925;
      115642:data<=-16'd2652;
      115643:data<=-16'd2725;
      115644:data<=-16'd2435;
      115645:data<=-16'd2554;
      115646:data<=-16'd3748;
      115647:data<=-16'd4115;
      115648:data<=-16'd3491;
      115649:data<=-16'd3099;
      115650:data<=-16'd2969;
      115651:data<=-16'd3530;
      115652:data<=-16'd4581;
      115653:data<=-16'd5109;
      115654:data<=-16'd5394;
      115655:data<=-16'd5747;
      115656:data<=-16'd5674;
      115657:data<=-16'd5473;
      115658:data<=-16'd5821;
      115659:data<=-16'd5723;
      115660:data<=-16'd5048;
      115661:data<=-16'd5817;
      115662:data<=-16'd6425;
      115663:data<=-16'd5059;
      115664:data<=-16'd5379;
      115665:data<=-16'd7515;
      115666:data<=-16'd7999;
      115667:data<=-16'd7691;
      115668:data<=-16'd7159;
      115669:data<=-16'd6448;
      115670:data<=-16'd6881;
      115671:data<=-16'd6953;
      115672:data<=-16'd6454;
      115673:data<=-16'd6815;
      115674:data<=-16'd6931;
      115675:data<=-16'd6645;
      115676:data<=-16'd6284;
      115677:data<=-16'd6358;
      115678:data<=-16'd8170;
      115679:data<=-16'd9397;
      115680:data<=-16'd8575;
      115681:data<=-16'd7749;
      115682:data<=-16'd7007;
      115683:data<=-16'd7015;
      115684:data<=-16'd8166;
      115685:data<=-16'd7987;
      115686:data<=-16'd7185;
      115687:data<=-16'd7356;
      115688:data<=-16'd6975;
      115689:data<=-16'd6238;
      115690:data<=-16'd6545;
      115691:data<=-16'd7583;
      115692:data<=-16'd8495;
      115693:data<=-16'd8755;
      115694:data<=-16'd8755;
      115695:data<=-16'd8537;
      115696:data<=-16'd7635;
      115697:data<=-16'd6942;
      115698:data<=-16'd6824;
      115699:data<=-16'd6399;
      115700:data<=-16'd6090;
      115701:data<=-16'd6182;
      115702:data<=-16'd5577;
      115703:data<=-16'd4952;
      115704:data<=-16'd5897;
      115705:data<=-16'd7495;
      115706:data<=-16'd8513;
      115707:data<=-16'd8628;
      115708:data<=-16'd7514;
      115709:data<=-16'd6669;
      115710:data<=-16'd6984;
      115711:data<=-16'd6811;
      115712:data<=-16'd6319;
      115713:data<=-16'd6404;
      115714:data<=-16'd6043;
      115715:data<=-16'd5106;
      115716:data<=-16'd4683;
      115717:data<=-16'd5574;
      115718:data<=-16'd7169;
      115719:data<=-16'd7755;
      115720:data<=-16'd7171;
      115721:data<=-16'd6354;
      115722:data<=-16'd6029;
      115723:data<=-16'd6170;
      115724:data<=-16'd5600;
      115725:data<=-16'd5063;
      115726:data<=-16'd5733;
      115727:data<=-16'd6128;
      115728:data<=-16'd5749;
      115729:data<=-16'd5092;
      115730:data<=-16'd4810;
      115731:data<=-16'd6258;
      115732:data<=-16'd7659;
      115733:data<=-16'd7131;
      115734:data<=-16'd6125;
      115735:data<=-16'd5247;
      115736:data<=-16'd5125;
      115737:data<=-16'd5921;
      115738:data<=-16'd5727;
      115739:data<=-16'd5007;
      115740:data<=-16'd4931;
      115741:data<=-16'd4849;
      115742:data<=-16'd4543;
      115743:data<=-16'd3829;
      115744:data<=-16'd3849;
      115745:data<=-16'd5644;
      115746:data<=-16'd6871;
      115747:data<=-16'd6146;
      115748:data<=-16'd4884;
      115749:data<=-16'd4504;
      115750:data<=-16'd5130;
      115751:data<=-16'd5100;
      115752:data<=-16'd4293;
      115753:data<=-16'd4297;
      115754:data<=-16'd4275;
      115755:data<=-16'd3121;
      115756:data<=-16'd2112;
      115757:data<=-16'd2874;
      115758:data<=-16'd4516;
      115759:data<=-16'd4613;
      115760:data<=-16'd4214;
      115761:data<=-16'd4948;
      115762:data<=-16'd4743;
      115763:data<=-16'd3633;
      115764:data<=-16'd3383;
      115765:data<=-16'd2948;
      115766:data<=-16'd2422;
      115767:data<=-16'd2646;
      115768:data<=-16'd2312;
      115769:data<=-16'd1639;
      115770:data<=-16'd2099;
      115771:data<=-16'd3269;
      115772:data<=-16'd4126;
      115773:data<=-16'd3711;
      115774:data<=-16'd2373;
      115775:data<=-16'd2390;
      115776:data<=-16'd2808;
      115777:data<=-16'd1240;
      115778:data<=-16'd472;
      115779:data<=-16'd1607;
      115780:data<=-16'd1501;
      115781:data<=-16'd917;
      115782:data<=-16'd599;
      115783:data<=16'd311;
      115784:data<=-16'd611;
      115785:data<=-16'd2438;
      115786:data<=-16'd2349;
      115787:data<=-16'd2191;
      115788:data<=-16'd2325;
      115789:data<=-16'd1933;
      115790:data<=-16'd1783;
      115791:data<=-16'd1098;
      115792:data<=-16'd400;
      115793:data<=-16'd875;
      115794:data<=-16'd1289;
      115795:data<=-16'd672;
      115796:data<=16'd312;
      115797:data<=-16'd376;
      115798:data<=-16'd2159;
      115799:data<=-16'd2147;
      115800:data<=-16'd1759;
      115801:data<=-16'd1970;
      115802:data<=-16'd873;
      115803:data<=16'd190;
      115804:data<=-16'd155;
      115805:data<=-16'd831;
      115806:data<=-16'd397;
      115807:data<=16'd1007;
      115808:data<=16'd832;
      115809:data<=16'd270;
      115810:data<=16'd752;
      115811:data<=-16'd705;
      115812:data<=-16'd1864;
      115813:data<=-16'd522;
      115814:data<=-16'd281;
      115815:data<=-16'd167;
      115816:data<=16'd887;
      115817:data<=16'd746;
      115818:data<=16'd375;
      115819:data<=-16'd199;
      115820:data<=-16'd321;
      115821:data<=16'd1503;
      115822:data<=16'd1921;
      115823:data<=16'd255;
      115824:data<=-16'd274;
      115825:data<=-16'd267;
      115826:data<=-16'd793;
      115827:data<=-16'd547;
      115828:data<=16'd479;
      115829:data<=16'd591;
      115830:data<=16'd168;
      115831:data<=16'd482;
      115832:data<=16'd230;
      115833:data<=-16'd117;
      115834:data<=16'd572;
      115835:data<=16'd732;
      115836:data<=16'd1237;
      115837:data<=16'd1811;
      115838:data<=16'd431;
      115839:data<=-16'd466;
      115840:data<=-16'd373;
      115841:data<=-16'd265;
      115842:data<=16'd970;
      115843:data<=16'd1119;
      115844:data<=16'd252;
      115845:data<=16'd1187;
      115846:data<=16'd1894;
      115847:data<=16'd881;
      115848:data<=16'd167;
      115849:data<=16'd1292;
      115850:data<=16'd2362;
      115851:data<=16'd1327;
      115852:data<=16'd1465;
      115853:data<=16'd2958;
      115854:data<=16'd3046;
      115855:data<=16'd3676;
      115856:data<=16'd3797;
      115857:data<=16'd3115;
      115858:data<=16'd3785;
      115859:data<=16'd2773;
      115860:data<=16'd2594;
      115861:data<=16'd4658;
      115862:data<=16'd3127;
      115863:data<=16'd3095;
      115864:data<=16'd6828;
      115865:data<=16'd6868;
      115866:data<=16'd6178;
      115867:data<=16'd7075;
      115868:data<=16'd6423;
      115869:data<=16'd5815;
      115870:data<=16'd5503;
      115871:data<=16'd5900;
      115872:data<=16'd6000;
      115873:data<=16'd4367;
      115874:data<=16'd5850;
      115875:data<=16'd7605;
      115876:data<=16'd5595;
      115877:data<=16'd6648;
      115878:data<=16'd8966;
      115879:data<=16'd7843;
      115880:data<=16'd8088;
      115881:data<=16'd9300;
      115882:data<=16'd8419;
      115883:data<=16'd7285;
      115884:data<=16'd7342;
      115885:data<=16'd8225;
      115886:data<=16'd8078;
      115887:data<=16'd7504;
      115888:data<=16'd7996;
      115889:data<=16'd8044;
      115890:data<=16'd8254;
      115891:data<=16'd9101;
      115892:data<=16'd9544;
      115893:data<=16'd10210;
      115894:data<=16'd9806;
      115895:data<=16'd8235;
      115896:data<=16'd7834;
      115897:data<=16'd8255;
      115898:data<=16'd8721;
      115899:data<=16'd8507;
      115900:data<=16'd7612;
      115901:data<=16'd7198;
      115902:data<=16'd6780;
      115903:data<=16'd7665;
      115904:data<=16'd9577;
      115905:data<=16'd8813;
      115906:data<=16'd7603;
      115907:data<=16'd8345;
      115908:data<=16'd8008;
      115909:data<=16'd6642;
      115910:data<=16'd6181;
      115911:data<=16'd6558;
      115912:data<=16'd6925;
      115913:data<=16'd6429;
      115914:data<=16'd6003;
      115915:data<=16'd6517;
      115916:data<=16'd7450;
      115917:data<=16'd7979;
      115918:data<=16'd7733;
      115919:data<=16'd8216;
      115920:data<=16'd8633;
      115921:data<=16'd6610;
      115922:data<=16'd5121;
      115923:data<=16'd6361;
      115924:data<=16'd7083;
      115925:data<=16'd6250;
      115926:data<=16'd5855;
      115927:data<=16'd5611;
      115928:data<=16'd4525;
      115929:data<=16'd4469;
      115930:data<=16'd6088;
      115931:data<=16'd6980;
      115932:data<=16'd6798;
      115933:data<=16'd6131;
      115934:data<=16'd5198;
      115935:data<=16'd4948;
      115936:data<=16'd4889;
      115937:data<=16'd4996;
      115938:data<=16'd4963;
      115939:data<=16'd4134;
      115940:data<=16'd4143;
      115941:data<=16'd3327;
      115942:data<=16'd1715;
      115943:data<=16'd3207;
      115944:data<=16'd4131;
      115945:data<=16'd3621;
      115946:data<=16'd5695;
      115947:data<=16'd6343;
      115948:data<=16'd5165;
      115949:data<=16'd4887;
      115950:data<=16'd3538;
      115951:data<=16'd3230;
      115952:data<=16'd3597;
      115953:data<=16'd2585;
      115954:data<=16'd3189;
      115955:data<=16'd3479;
      115956:data<=16'd3018;
      115957:data<=16'd4919;
      115958:data<=16'd5560;
      115959:data<=16'd4085;
      115960:data<=16'd4481;
      115961:data<=16'd6159;
      115962:data<=16'd5412;
      115963:data<=16'd2855;
      115964:data<=16'd3580;
      115965:data<=16'd5172;
      115966:data<=16'd3764;
      115967:data<=16'd3025;
      115968:data<=16'd2215;
      115969:data<=16'd2326;
      115970:data<=16'd5703;
      115971:data<=16'd5418;
      115972:data<=16'd3109;
      115973:data<=16'd3474;
      115974:data<=16'd1958;
      115975:data<=16'd933;
      115976:data<=16'd1889;
      115977:data<=16'd1524;
      115978:data<=16'd2015;
      115979:data<=16'd2199;
      115980:data<=16'd1365;
      115981:data<=16'd1281;
      115982:data<=16'd455;
      115983:data<=16'd1049;
      115984:data<=16'd3227;
      115985:data<=16'd3219;
      115986:data<=-16'd18;
      115987:data<=-16'd5028;
      115988:data<=-16'd6675;
      115989:data<=-16'd6231;
      115990:data<=-16'd7518;
      115991:data<=-16'd6282;
      115992:data<=-16'd4855;
      115993:data<=-16'd5896;
      115994:data<=-16'd5530;
      115995:data<=-16'd5891;
      115996:data<=-16'd6125;
      115997:data<=-16'd4622;
      115998:data<=-16'd3808;
      115999:data<=-16'd2634;
      116000:data<=-16'd3668;
      116001:data<=-16'd4875;
      116002:data<=-16'd2710;
      116003:data<=-16'd3427;
      116004:data<=-16'd3694;
      116005:data<=-16'd1477;
      116006:data<=-16'd3128;
      116007:data<=-16'd4000;
      116008:data<=-16'd3935;
      116009:data<=-16'd3356;
      116010:data<=16'd2564;
      116011:data<=16'd4710;
      116012:data<=16'd326;
      116013:data<=-16'd3744;
      116014:data<=-16'd6860;
      116015:data<=-16'd6219;
      116016:data<=-16'd5069;
      116017:data<=-16'd5767;
      116018:data<=-16'd3224;
      116019:data<=16'd578;
      116020:data<=16'd4322;
      116021:data<=16'd3767;
      116022:data<=16'd1670;
      116023:data<=16'd11338;
      116024:data<=16'd16610;
      116025:data<=16'd6992;
      116026:data<=16'd4024;
      116027:data<=16'd4764;
      116028:data<=16'd259;
      116029:data<=-16'd138;
      116030:data<=16'd2117;
      116031:data<=16'd5075;
      116032:data<=16'd6279;
      116033:data<=16'd1982;
      116034:data<=-16'd135;
      116035:data<=16'd161;
      116036:data<=-16'd1221;
      116037:data<=-16'd1753;
      116038:data<=16'd1184;
      116039:data<=16'd5970;
      116040:data<=16'd2696;
      116041:data<=-16'd3190;
      116042:data<=-16'd647;
      116043:data<=-16'd3413;
      116044:data<=-16'd12957;
      116045:data<=-16'd16977;
      116046:data<=-16'd19064;
      116047:data<=-16'd21696;
      116048:data<=-16'd25388;
      116049:data<=-16'd25299;
      116050:data<=-16'd16769;
      116051:data<=-16'd13110;
      116052:data<=-16'd16183;
      116053:data<=-16'd18806;
      116054:data<=-16'd20019;
      116055:data<=-16'd15723;
      116056:data<=-16'd15153;
      116057:data<=-16'd17750;
      116058:data<=-16'd12455;
      116059:data<=-16'd10863;
      116060:data<=-16'd10437;
      116061:data<=-16'd8784;
      116062:data<=-16'd16337;
      116063:data<=-16'd13289;
      116064:data<=-16'd3815;
      116065:data<=-16'd11435;
      116066:data<=-16'd18829;
      116067:data<=-16'd21100;
      116068:data<=-16'd22946;
      116069:data<=-16'd17256;
      116070:data<=-16'd15053;
      116071:data<=-16'd14055;
      116072:data<=-16'd11242;
      116073:data<=-16'd16084;
      116074:data<=-16'd16736;
      116075:data<=-16'd15474;
      116076:data<=-16'd19378;
      116077:data<=-16'd18618;
      116078:data<=-16'd21675;
      116079:data<=-16'd26538;
      116080:data<=-16'd24090;
      116081:data<=-16'd22151;
      116082:data<=-16'd16583;
      116083:data<=-16'd13509;
      116084:data<=-16'd15406;
      116085:data<=-16'd5036;
      116086:data<=16'd1177;
      116087:data<=-16'd4426;
      116088:data<=-16'd1397;
      116089:data<=16'd1162;
      116090:data<=16'd140;
      116091:data<=16'd5101;
      116092:data<=16'd5711;
      116093:data<=16'd2775;
      116094:data<=16'd3588;
      116095:data<=16'd4946;
      116096:data<=16'd5096;
      116097:data<=16'd3579;
      116098:data<=16'd1524;
      116099:data<=-16'd2701;
      116100:data<=-16'd3791;
      116101:data<=16'd3052;
      116102:data<=16'd2165;
      116103:data<=-16'd2699;
      116104:data<=16'd901;
      116105:data<=-16'd3093;
      116106:data<=-16'd10466;
      116107:data<=-16'd8052;
      116108:data<=-16'd5300;
      116109:data<=16'd822;
      116110:data<=16'd3758;
      116111:data<=-16'd6711;
      116112:data<=-16'd8678;
      116113:data<=-16'd3083;
      116114:data<=-16'd8990;
      116115:data<=-16'd13308;
      116116:data<=-16'd7885;
      116117:data<=-16'd3051;
      116118:data<=-16'd2299;
      116119:data<=-16'd3795;
      116120:data<=-16'd3627;
      116121:data<=-16'd2138;
      116122:data<=-16'd632;
      116123:data<=16'd1530;
      116124:data<=16'd778;
      116125:data<=16'd3983;
      116126:data<=16'd12398;
      116127:data<=16'd4910;
      116128:data<=-16'd10079;
      116129:data<=-16'd4667;
      116130:data<=16'd2494;
      116131:data<=-16'd6789;
      116132:data<=-16'd9080;
      116133:data<=-16'd4417;
      116134:data<=-16'd8455;
      116135:data<=-16'd8234;
      116136:data<=-16'd5333;
      116137:data<=-16'd7594;
      116138:data<=16'd39;
      116139:data<=16'd6654;
      116140:data<=16'd253;
      116141:data<=16'd570;
      116142:data<=16'd2036;
      116143:data<=-16'd1472;
      116144:data<=16'd5165;
      116145:data<=16'd6667;
      116146:data<=-16'd591;
      116147:data<=16'd2440;
      116148:data<=16'd4099;
      116149:data<=16'd3219;
      116150:data<=16'd8046;
      116151:data<=16'd4449;
      116152:data<=16'd1512;
      116153:data<=16'd6184;
      116154:data<=16'd2742;
      116155:data<=16'd3544;
      116156:data<=16'd11092;
      116157:data<=16'd6070;
      116158:data<=16'd4043;
      116159:data<=16'd14242;
      116160:data<=16'd15358;
      116161:data<=16'd9764;
      116162:data<=16'd10014;
      116163:data<=16'd8413;
      116164:data<=16'd5007;
      116165:data<=16'd10288;
      116166:data<=16'd16686;
      116167:data<=16'd12643;
      116168:data<=16'd7861;
      116169:data<=16'd13735;
      116170:data<=16'd24344;
      116171:data<=16'd27972;
      116172:data<=16'd24234;
      116173:data<=16'd23358;
      116174:data<=16'd21998;
      116175:data<=16'd13201;
      116176:data<=16'd10795;
      116177:data<=16'd15713;
      116178:data<=16'd14001;
      116179:data<=16'd12737;
      116180:data<=16'd15042;
      116181:data<=16'd13226;
      116182:data<=16'd13279;
      116183:data<=16'd15826;
      116184:data<=16'd14762;
      116185:data<=16'd13171;
      116186:data<=16'd11200;
      116187:data<=16'd7172;
      116188:data<=16'd6331;
      116189:data<=16'd9570;
      116190:data<=16'd10364;
      116191:data<=16'd11920;
      116192:data<=16'd18553;
      116193:data<=16'd17337;
      116194:data<=16'd11724;
      116195:data<=16'd17370;
      116196:data<=16'd16868;
      116197:data<=16'd4781;
      116198:data<=16'd4819;
      116199:data<=16'd10954;
      116200:data<=16'd9000;
      116201:data<=16'd5717;
      116202:data<=16'd5826;
      116203:data<=16'd9655;
      116204:data<=16'd11536;
      116205:data<=16'd10793;
      116206:data<=16'd12325;
      116207:data<=16'd8075;
      116208:data<=16'd3172;
      116209:data<=16'd6801;
      116210:data<=16'd5162;
      116211:data<=-16'd1656;
      116212:data<=-16'd5685;
      116213:data<=-16'd11309;
      116214:data<=-16'd11697;
      116215:data<=-16'd5006;
      116216:data<=-16'd3163;
      116217:data<=-16'd7001;
      116218:data<=-16'd8082;
      116219:data<=-16'd4737;
      116220:data<=-16'd5406;
      116221:data<=-16'd7602;
      116222:data<=-16'd4952;
      116223:data<=-16'd6304;
      116224:data<=-16'd4831;
      116225:data<=16'd4356;
      116226:data<=16'd4085;
      116227:data<=16'd3704;
      116228:data<=16'd10892;
      116229:data<=16'd8038;
      116230:data<=16'd1403;
      116231:data<=-16'd851;
      116232:data<=-16'd3319;
      116233:data<=-16'd2607;
      116234:data<=-16'd2488;
      116235:data<=-16'd196;
      116236:data<=16'd7235;
      116237:data<=16'd5001;
      116238:data<=-16'd3453;
      116239:data<=-16'd5450;
      116240:data<=-16'd4211;
      116241:data<=-16'd3204;
      116242:data<=-16'd3008;
      116243:data<=-16'd623;
      116244:data<=-16'd440;
      116245:data<=-16'd8023;
      116246:data<=-16'd8486;
      116247:data<=-16'd3627;
      116248:data<=-16'd8690;
      116249:data<=-16'd10082;
      116250:data<=-16'd3560;
      116251:data<=-16'd5148;
      116252:data<=-16'd7288;
      116253:data<=16'd4173;
      116254:data<=16'd15065;
      116255:data<=16'd11133;
      116256:data<=16'd10575;
      116257:data<=16'd16954;
      116258:data<=16'd9078;
      116259:data<=16'd4053;
      116260:data<=16'd12787;
      116261:data<=16'd8445;
      116262:data<=16'd2877;
      116263:data<=16'd11103;
      116264:data<=16'd9970;
      116265:data<=16'd2934;
      116266:data<=16'd2974;
      116267:data<=16'd1016;
      116268:data<=-16'd796;
      116269:data<=16'd3400;
      116270:data<=16'd6246;
      116271:data<=16'd1773;
      116272:data<=-16'd1125;
      116273:data<=16'd2555;
      116274:data<=-16'd390;
      116275:data<=-16'd5251;
      116276:data<=-16'd2707;
      116277:data<=-16'd8475;
      116278:data<=-16'd17738;
      116279:data<=-16'd15321;
      116280:data<=-16'd10795;
      116281:data<=-16'd9213;
      116282:data<=-16'd10558;
      116283:data<=-16'd12160;
      116284:data<=-16'd9320;
      116285:data<=-16'd11888;
      116286:data<=-16'd15235;
      116287:data<=-16'd11424;
      116288:data<=-16'd12081;
      116289:data<=-16'd9782;
      116290:data<=-16'd2864;
      116291:data<=-16'd9448;
      116292:data<=-16'd17785;
      116293:data<=-16'd14578;
      116294:data<=-16'd10675;
      116295:data<=-16'd14334;
      116296:data<=-16'd26554;
      116297:data<=-16'd33386;
      116298:data<=-16'd27223;
      116299:data<=-16'd24539;
      116300:data<=-16'd26177;
      116301:data<=-16'd22380;
      116302:data<=-16'd20287;
      116303:data<=-16'd23247;
      116304:data<=-16'd22375;
      116305:data<=-16'd16847;
      116306:data<=-16'd19658;
      116307:data<=-16'd27616;
      116308:data<=-16'd24118;
      116309:data<=-16'd21238;
      116310:data<=-16'd26100;
      116311:data<=-16'd21281;
      116312:data<=-16'd16651;
      116313:data<=-16'd22213;
      116314:data<=-16'd21312;
      116315:data<=-16'd14078;
      116316:data<=-16'd10936;
      116317:data<=-16'd13717;
      116318:data<=-16'd17145;
      116319:data<=-16'd15214;
      116320:data<=-16'd18236;
      116321:data<=-16'd21435;
      116322:data<=-16'd11430;
      116323:data<=-16'd10715;
      116324:data<=-16'd19159;
      116325:data<=-16'd10577;
      116326:data<=-16'd1742;
      116327:data<=-16'd2749;
      116328:data<=16'd1666;
      116329:data<=16'd2090;
      116330:data<=-16'd3442;
      116331:data<=-16'd1710;
      116332:data<=16'd2484;
      116333:data<=16'd3852;
      116334:data<=16'd3519;
      116335:data<=16'd1146;
      116336:data<=16'd631;
      116337:data<=16'd5447;
      116338:data<=16'd12369;
      116339:data<=16'd15873;
      116340:data<=16'd18468;
      116341:data<=16'd21631;
      116342:data<=16'd18691;
      116343:data<=16'd15646;
      116344:data<=16'd19331;
      116345:data<=16'd21930;
      116346:data<=16'd22312;
      116347:data<=16'd19050;
      116348:data<=16'd11038;
      116349:data<=16'd10997;
      116350:data<=16'd15465;
      116351:data<=16'd11966;
      116352:data<=16'd8818;
      116353:data<=16'd10753;
      116354:data<=16'd12862;
      116355:data<=16'd16010;
      116356:data<=16'd18524;
      116357:data<=16'd17705;
      116358:data<=16'd16019;
      116359:data<=16'd17014;
      116360:data<=16'd19036;
      116361:data<=16'd15462;
      116362:data<=16'd9762;
      116363:data<=16'd11145;
      116364:data<=16'd15274;
      116365:data<=16'd15987;
      116366:data<=16'd16959;
      116367:data<=16'd17937;
      116368:data<=16'd14581;
      116369:data<=16'd9806;
      116370:data<=16'd7815;
      116371:data<=16'd8528;
      116372:data<=16'd10887;
      116373:data<=16'd12598;
      116374:data<=16'd12966;
      116375:data<=16'd8452;
      116376:data<=-16'd1248;
      116377:data<=16'd1949;
      116378:data<=16'd13361;
      116379:data<=16'd3143;
      116380:data<=-16'd13878;
      116381:data<=-16'd16098;
      116382:data<=-16'd17199;
      116383:data<=-16'd12508;
      116384:data<=-16'd4034;
      116385:data<=-16'd7344;
      116386:data<=-16'd5792;
      116387:data<=-16'd1519;
      116388:data<=-16'd6840;
      116389:data<=-16'd4752;
      116390:data<=-16'd3817;
      116391:data<=-16'd11015;
      116392:data<=-16'd7000;
      116393:data<=-16'd688;
      116394:data<=-16'd1306;
      116395:data<=-16'd3577;
      116396:data<=-16'd7417;
      116397:data<=-16'd2187;
      116398:data<=16'd5139;
      116399:data<=16'd419;
      116400:data<=-16'd1735;
      116401:data<=16'd1850;
      116402:data<=16'd2093;
      116403:data<=16'd1677;
      116404:data<=16'd262;
      116405:data<=-16'd1155;
      116406:data<=16'd996;
      116407:data<=16'd5833;
      116408:data<=16'd5350;
      116409:data<=-16'd3313;
      116410:data<=-16'd1806;
      116411:data<=16'd7347;
      116412:data<=16'd4074;
      116413:data<=16'd1610;
      116414:data<=16'd6202;
      116415:data<=16'd7078;
      116416:data<=16'd8267;
      116417:data<=16'd7195;
      116418:data<=16'd6640;
      116419:data<=16'd8636;
      116420:data<=16'd4382;
      116421:data<=16'd10184;
      116422:data<=16'd21960;
      116423:data<=16'd17390;
      116424:data<=16'd18393;
      116425:data<=16'd27830;
      116426:data<=16'd25631;
      116427:data<=16'd24388;
      116428:data<=16'd25364;
      116429:data<=16'd24432;
      116430:data<=16'd28107;
      116431:data<=16'd28758;
      116432:data<=16'd29207;
      116433:data<=16'd27943;
      116434:data<=16'd18613;
      116435:data<=16'd19230;
      116436:data<=16'd22971;
      116437:data<=16'd14684;
      116438:data<=16'd13899;
      116439:data<=16'd19801;
      116440:data<=16'd17095;
      116441:data<=16'd13191;
      116442:data<=16'd12922;
      116443:data<=16'd13030;
      116444:data<=16'd11471;
      116445:data<=16'd10822;
      116446:data<=16'd10560;
      116447:data<=16'd6819;
      116448:data<=16'd10683;
      116449:data<=16'd14774;
      116450:data<=16'd1296;
      116451:data<=-16'd4147;
      116452:data<=16'd6299;
      116453:data<=16'd4623;
      116454:data<=-16'd2602;
      116455:data<=-16'd2413;
      116456:data<=16'd147;
      116457:data<=16'd1770;
      116458:data<=-16'd1985;
      116459:data<=-16'd1876;
      116460:data<=16'd415;
      116461:data<=-16'd6024;
      116462:data<=-16'd1666;
      116463:data<=16'd4046;
      116464:data<=-16'd13303;
      116465:data<=-16'd24780;
      116466:data<=-16'd23783;
      116467:data<=-16'd27223;
      116468:data<=-16'd19238;
      116469:data<=-16'd10746;
      116470:data<=-16'd19450;
      116471:data<=-16'd23910;
      116472:data<=-16'd18936;
      116473:data<=-16'd15603;
      116474:data<=-16'd16659;
      116475:data<=-16'd23643;
      116476:data<=-16'd27995;
      116477:data<=-16'd24938;
      116478:data<=-16'd21667;
      116479:data<=-16'd24415;
      116480:data<=-16'd30426;
      116481:data<=-16'd27492;
      116482:data<=-16'd23135;
      116483:data<=-16'd27513;
      116484:data<=-16'd23388;
      116485:data<=-16'd18139;
      116486:data<=-16'd28172;
      116487:data<=-16'd30236;
      116488:data<=-16'd20274;
      116489:data<=-16'd18084;
      116490:data<=-16'd20964;
      116491:data<=-16'd25314;
      116492:data<=-16'd27395;
      116493:data<=-16'd21094;
      116494:data<=-16'd16681;
      116495:data<=-16'd16319;
      116496:data<=-16'd14155;
      116497:data<=-16'd18130;
      116498:data<=-16'd25002;
      116499:data<=-16'd20436;
      116500:data<=-16'd13391;
      116501:data<=-16'd15264;
      116502:data<=-16'd13297;
      116503:data<=-16'd9398;
      116504:data<=-16'd16365;
      116505:data<=-16'd13045;
      116506:data<=16'd4438;
      116507:data<=16'd5479;
      116508:data<=16'd954;
      116509:data<=16'd7908;
      116510:data<=16'd6639;
      116511:data<=16'd2905;
      116512:data<=16'd6610;
      116513:data<=16'd1920;
      116514:data<=-16'd1263;
      116515:data<=16'd4176;
      116516:data<=16'd884;
      116517:data<=-16'd2992;
      116518:data<=-16'd638;
      116519:data<=-16'd3442;
      116520:data<=-16'd3815;
      116521:data<=-16'd1068;
      116522:data<=-16'd2285;
      116523:data<=16'd1994;
      116524:data<=16'd3548;
      116525:data<=-16'd1568;
      116526:data<=16'd6064;
      116527:data<=16'd12387;
      116528:data<=16'd3921;
      116529:data<=16'd1733;
      116530:data<=16'd1914;
      116531:data<=-16'd2977;
      116532:data<=16'd769;
      116533:data<=16'd6575;
      116534:data<=16'd7809;
      116535:data<=16'd6223;
      116536:data<=-16'd1501;
      116537:data<=-16'd3359;
      116538:data<=16'd1486;
      116539:data<=16'd635;
      116540:data<=16'd1895;
      116541:data<=16'd4041;
      116542:data<=-16'd1780;
      116543:data<=-16'd5641;
      116544:data<=-16'd3436;
      116545:data<=-16'd2397;
      116546:data<=-16'd5198;
      116547:data<=-16'd7122;
      116548:data<=-16'd9277;
      116549:data<=-16'd19227;
      116550:data<=-16'd20729;
      116551:data<=-16'd7467;
      116552:data<=-16'd7230;
      116553:data<=-16'd12904;
      116554:data<=-16'd6760;
      116555:data<=-16'd8381;
      116556:data<=-16'd12346;
      116557:data<=-16'd5118;
      116558:data<=-16'd6264;
      116559:data<=-16'd12387;
      116560:data<=-16'd8049;
      116561:data<=-16'd6851;
      116562:data<=-16'd12051;
      116563:data<=-16'd8449;
      116564:data<=16'd543;
      116565:data<=16'd2029;
      116566:data<=-16'd1108;
      116567:data<=-16'd2896;
      116568:data<=-16'd3410;
      116569:data<=-16'd761;
      116570:data<=16'd2238;
      116571:data<=16'd4087;
      116572:data<=16'd6190;
      116573:data<=16'd2153;
      116574:data<=-16'd469;
      116575:data<=16'd4211;
      116576:data<=-16'd1507;
      116577:data<=-16'd8627;
      116578:data<=-16'd746;
      116579:data<=16'd1116;
      116580:data<=-16'd4288;
      116581:data<=-16'd713;
      116582:data<=16'd359;
      116583:data<=-16'd2532;
      116584:data<=-16'd297;
      116585:data<=16'd579;
      116586:data<=16'd2664;
      116587:data<=16'd6555;
      116588:data<=16'd2422;
      116589:data<=16'd4008;
      116590:data<=16'd17494;
      116591:data<=16'd18776;
      116592:data<=16'd16199;
      116593:data<=16'd27883;
      116594:data<=16'd26321;
      116595:data<=16'd12919;
      116596:data<=16'd17475;
      116597:data<=16'd20237;
      116598:data<=16'd14082;
      116599:data<=16'd17887;
      116600:data<=16'd17047;
      116601:data<=16'd15435;
      116602:data<=16'd22870;
      116603:data<=16'd18648;
      116604:data<=16'd15427;
      116605:data<=16'd21463;
      116606:data<=16'd16477;
      116607:data<=16'd15767;
      116608:data<=16'd19355;
      116609:data<=16'd11144;
      116610:data<=16'd12945;
      116611:data<=16'd18621;
      116612:data<=16'd12507;
      116613:data<=16'd15209;
      116614:data<=16'd18516;
      116615:data<=16'd13136;
      116616:data<=16'd17942;
      116617:data<=16'd22924;
      116618:data<=16'd17453;
      116619:data<=16'd13797;
      116620:data<=16'd14706;
      116621:data<=16'd17132;
      116622:data<=16'd15352;
      116623:data<=16'd11721;
      116624:data<=16'd12722;
      116625:data<=16'd10116;
      116626:data<=16'd11681;
      116627:data<=16'd22013;
      116628:data<=16'd18554;
      116629:data<=16'd12217;
      116630:data<=16'd20804;
      116631:data<=16'd20428;
      116632:data<=16'd6907;
      116633:data<=16'd1110;
      116634:data<=16'd3921;
      116635:data<=16'd3906;
      116636:data<=-16'd2943;
      116637:data<=-16'd1753;
      116638:data<=16'd8995;
      116639:data<=16'd5903;
      116640:data<=-16'd2823;
      116641:data<=16'd811;
      116642:data<=16'd1154;
      116643:data<=-16'd4519;
      116644:data<=-16'd1909;
      116645:data<=16'd3604;
      116646:data<=16'd2343;
      116647:data<=-16'd1054;
      116648:data<=16'd1334;
      116649:data<=16'd3565;
      116650:data<=16'd20;
      116651:data<=16'd555;
      116652:data<=16'd2328;
      116653:data<=-16'd4481;
      116654:data<=-16'd7674;
      116655:data<=-16'd83;
      116656:data<=16'd4538;
      116657:data<=-16'd908;
      116658:data<=-16'd6123;
      116659:data<=-16'd3084;
      116660:data<=-16'd164;
      116661:data<=-16'd1242;
      116662:data<=16'd112;
      116663:data<=-16'd857;
      116664:data<=-16'd5247;
      116665:data<=-16'd3500;
      116666:data<=-16'd2208;
      116667:data<=-16'd7709;
      116668:data<=-16'd5338;
      116669:data<=16'd3770;
      116670:data<=-16'd640;
      116671:data<=-16'd10796;
      116672:data<=-16'd10604;
      116673:data<=-16'd8009;
      116674:data<=-16'd185;
      116675:data<=16'd12627;
      116676:data<=16'd9104;
      116677:data<=16'd159;
      116678:data<=16'd2024;
      116679:data<=-16'd1589;
      116680:data<=-16'd7030;
      116681:data<=-16'd4640;
      116682:data<=-16'd6229;
      116683:data<=-16'd8822;
      116684:data<=-16'd5510;
      116685:data<=-16'd1765;
      116686:data<=-16'd2858;
      116687:data<=-16'd8208;
      116688:data<=-16'd5489;
      116689:data<=16'd2165;
      116690:data<=-16'd2265;
      116691:data<=-16'd8804;
      116692:data<=-16'd6990;
      116693:data<=-16'd5510;
      116694:data<=-16'd4105;
      116695:data<=-16'd1145;
      116696:data<=-16'd1671;
      116697:data<=-16'd4059;
      116698:data<=-16'd4020;
      116699:data<=-16'd4185;
      116700:data<=-16'd6326;
      116701:data<=-16'd6851;
      116702:data<=-16'd9404;
      116703:data<=-16'd12023;
      116704:data<=-16'd7447;
      116705:data<=-16'd7336;
      116706:data<=-16'd9594;
      116707:data<=-16'd3286;
      116708:data<=-16'd2896;
      116709:data<=-16'd3747;
      116710:data<=16'd778;
      116711:data<=-16'd5034;
      116712:data<=-16'd7178;
      116713:data<=-16'd2711;
      116714:data<=-16'd9307;
      116715:data<=-16'd12202;
      116716:data<=-16'd13333;
      116717:data<=-16'd22348;
      116718:data<=-16'd23378;
      116719:data<=-16'd23777;
      116720:data<=-16'd28019;
      116721:data<=-16'd24838;
      116722:data<=-16'd21626;
      116723:data<=-16'd21652;
      116724:data<=-16'd25350;
      116725:data<=-16'd26467;
      116726:data<=-16'd14410;
      116727:data<=-16'd8276;
      116728:data<=-16'd12810;
      116729:data<=-16'd11571;
      116730:data<=-16'd9505;
      116731:data<=-16'd6205;
      116732:data<=-16'd3284;
      116733:data<=-16'd8392;
      116734:data<=-16'd9486;
      116735:data<=-16'd7045;
      116736:data<=-16'd8736;
      116737:data<=-16'd9262;
      116738:data<=-16'd8758;
      116739:data<=-16'd6141;
      116740:data<=-16'd4886;
      116741:data<=-16'd7806;
      116742:data<=-16'd6839;
      116743:data<=-16'd6695;
      116744:data<=-16'd7874;
      116745:data<=-16'd4087;
      116746:data<=-16'd3677;
      116747:data<=-16'd7453;
      116748:data<=-16'd9034;
      116749:data<=-16'd4331;
      116750:data<=16'd364;
      116751:data<=-16'd7768;
      116752:data<=-16'd9878;
      116753:data<=16'd623;
      116754:data<=-16'd429;
      116755:data<=-16'd3401;
      116756:data<=-16'd3153;
      116757:data<=-16'd6551;
      116758:data<=16'd3312;
      116759:data<=16'd14487;
      116760:data<=16'd14063;
      116761:data<=16'd13535;
      116762:data<=16'd9532;
      116763:data<=16'd13265;
      116764:data<=16'd20554;
      116765:data<=16'd10607;
      116766:data<=16'd8652;
      116767:data<=16'd16134;
      116768:data<=16'd10937;
      116769:data<=16'd8144;
      116770:data<=16'd8978;
      116771:data<=16'd12819;
      116772:data<=16'd20654;
      116773:data<=16'd13593;
      116774:data<=16'd9165;
      116775:data<=16'd17728;
      116776:data<=16'd16269;
      116777:data<=16'd10812;
      116778:data<=16'd4889;
      116779:data<=16'd83;
      116780:data<=16'd6438;
      116781:data<=16'd6608;
      116782:data<=16'd4705;
      116783:data<=16'd12731;
      116784:data<=16'd11304;
      116785:data<=16'd5488;
      116786:data<=16'd4252;
      116787:data<=16'd974;
      116788:data<=16'd3052;
      116789:data<=16'd7115;
      116790:data<=16'd10593;
      116791:data<=16'd13526;
      116792:data<=16'd7124;
      116793:data<=16'd7010;
      116794:data<=16'd12267;
      116795:data<=16'd3830;
      116796:data<=16'd848;
      116797:data<=16'd7794;
      116798:data<=16'd8479;
      116799:data<=16'd7200;
      116800:data<=16'd89;
      116801:data<=-16'd8345;
      116802:data<=-16'd6863;
      116803:data<=-16'd5943;
      116804:data<=-16'd4543;
      116805:data<=-16'd3586;
      116806:data<=-16'd9900;
      116807:data<=-16'd7717;
      116808:data<=-16'd1577;
      116809:data<=-16'd3667;
      116810:data<=16'd39;
      116811:data<=16'd4270;
      116812:data<=16'd585;
      116813:data<=16'd408;
      116814:data<=-16'd241;
      116815:data<=-16'd4203;
      116816:data<=-16'd3686;
      116817:data<=-16'd1368;
      116818:data<=16'd704;
      116819:data<=16'd2361;
      116820:data<=16'd1434;
      116821:data<=16'd268;
      116822:data<=16'd2355;
      116823:data<=16'd5177;
      116824:data<=16'd100;
      116825:data<=-16'd3133;
      116826:data<=16'd9576;
      116827:data<=16'd16301;
      116828:data<=16'd8608;
      116829:data<=16'd10228;
      116830:data<=16'd15864;
      116831:data<=16'd12787;
      116832:data<=16'd8008;
      116833:data<=16'd5165;
      116834:data<=16'd8608;
      116835:data<=16'd11300;
      116836:data<=16'd9197;
      116837:data<=16'd16509;
      116838:data<=16'd19136;
      116839:data<=16'd9480;
      116840:data<=16'd10445;
      116841:data<=16'd12205;
      116842:data<=16'd11781;
      116843:data<=16'd24839;
      116844:data<=16'd28128;
      116845:data<=16'd21567;
      116846:data<=16'd28459;
      116847:data<=16'd29959;
      116848:data<=16'd23027;
      116849:data<=16'd24771;
      116850:data<=16'd24539;
      116851:data<=16'd20948;
      116852:data<=16'd21029;
      116853:data<=16'd18882;
      116854:data<=16'd17896;
      116855:data<=16'd21535;
      116856:data<=16'd21936;
      116857:data<=16'd18095;
      116858:data<=16'd18591;
      116859:data<=16'd22063;
      116860:data<=16'd18174;
      116861:data<=16'd13420;
      116862:data<=16'd15324;
      116863:data<=16'd14798;
      116864:data<=16'd13236;
      116865:data<=16'd14786;
      116866:data<=16'd14650;
      116867:data<=16'd14149;
      116868:data<=16'd10530;
      116869:data<=16'd5785;
      116870:data<=16'd7926;
      116871:data<=16'd7633;
      116872:data<=16'd5190;
      116873:data<=16'd8943;
      116874:data<=16'd8243;
      116875:data<=16'd5406;
      116876:data<=16'd6476;
      116877:data<=-16'd1580;
      116878:data<=-16'd11753;
      116879:data<=-16'd9338;
      116880:data<=-16'd5216;
      116881:data<=-16'd6757;
      116882:data<=-16'd7952;
      116883:data<=-16'd10599;
      116884:data<=-16'd19519;
      116885:data<=-16'd27761;
      116886:data<=-16'd27234;
      116887:data<=-16'd24404;
      116888:data<=-16'd25167;
      116889:data<=-16'd25261;
      116890:data<=-16'd23819;
      116891:data<=-16'd23497;
      116892:data<=-16'd25062;
      116893:data<=-16'd24416;
      116894:data<=-16'd19241;
      116895:data<=-16'd19265;
      116896:data<=-16'd23555;
      116897:data<=-16'd19070;
      116898:data<=-16'd13849;
      116899:data<=-16'd18768;
      116900:data<=-16'd23276;
      116901:data<=-16'd20130;
      116902:data<=-16'd17004;
      116903:data<=-16'd19804;
      116904:data<=-16'd22645;
      116905:data<=-16'd21634;
      116906:data<=-16'd21819;
      116907:data<=-16'd21185;
      116908:data<=-16'd18042;
      116909:data<=-16'd16989;
      116910:data<=-16'd16208;
      116911:data<=-16'd15913;
      116912:data<=-16'd15070;
      116913:data<=-16'd12232;
      116914:data<=-16'd15479;
      116915:data<=-16'd17617;
      116916:data<=-16'd13998;
      116917:data<=-16'd18506;
      116918:data<=-16'd19281;
      116919:data<=-16'd9592;
      116920:data<=-16'd9623;
      116921:data<=-16'd13668;
      116922:data<=-16'd14515;
      116923:data<=-16'd17286;
      116924:data<=-16'd14754;
      116925:data<=-16'd14314;
      116926:data<=-16'd13370;
      116927:data<=16'd4889;
      116928:data<=16'd18956;
      116929:data<=16'd15320;
      116930:data<=16'd12451;
      116931:data<=16'd13459;
      116932:data<=16'd14020;
      116933:data<=16'd10064;
      116934:data<=16'd3228;
      116935:data<=16'd5024;
      116936:data<=16'd9647;
      116937:data<=16'd10921;
      116938:data<=16'd9658;
      116939:data<=16'd1384;
      116940:data<=-16'd1077;
      116941:data<=16'd5768;
      116942:data<=16'd6805;
      116943:data<=16'd5806;
      116944:data<=16'd4375;
      116945:data<=16'd890;
      116946:data<=16'd582;
      116947:data<=-16'd2629;
      116948:data<=-16'd3802;
      116949:data<=16'd376;
      116950:data<=16'd282;
      116951:data<=16'd3063;
      116952:data<=16'd3755;
      116953:data<=-16'd958;
      116954:data<=16'd4739;
      116955:data<=16'd2819;
      116956:data<=-16'd9098;
      116957:data<=-16'd4003;
      116958:data<=16'd24;
      116959:data<=-16'd3562;
      116960:data<=16'd2135;
      116961:data<=16'd922;
      116962:data<=-16'd3436;
      116963:data<=16'd1680;
      116964:data<=16'd616;
      116965:data<=-16'd2564;
      116966:data<=-16'd930;
      116967:data<=-16'd2217;
      116968:data<=-16'd7291;
      116969:data<=-16'd18494;
      116970:data<=-16'd23047;
      116971:data<=-16'd14246;
      116972:data<=-16'd14254;
      116973:data<=-16'd18166;
      116974:data<=-16'd12813;
      116975:data<=-16'd14005;
      116976:data<=-16'd19526;
      116977:data<=-16'd18266;
      116978:data<=-16'd17603;
      116979:data<=-16'd19114;
      116980:data<=-16'd19667;
      116981:data<=-16'd17452;
      116982:data<=-16'd13344;
      116983:data<=-16'd14929;
      116984:data<=-16'd17447;
      116985:data<=-16'd13012;
      116986:data<=-16'd10413;
      116987:data<=-16'd11529;
      116988:data<=-16'd8247;
      116989:data<=-16'd5682;
      116990:data<=-16'd7750;
      116991:data<=-16'd5847;
      116992:data<=-16'd3336;
      116993:data<=-16'd7031;
      116994:data<=-16'd5835;
      116995:data<=-16'd861;
      116996:data<=-16'd4094;
      116997:data<=-16'd6176;
      116998:data<=-16'd4592;
      116999:data<=-16'd5877;
      117000:data<=-16'd892;
      117001:data<=16'd2992;
      117002:data<=-16'd3674;
      117003:data<=-16'd3864;
      117004:data<=-16'd136;
      117005:data<=-16'd2692;
      117006:data<=16'd873;
      117007:data<=16'd4470;
      117008:data<=-16'd1064;
      117009:data<=16'd544;
      117010:data<=16'd10934;
      117011:data<=16'd17744;
      117012:data<=16'd20527;
      117013:data<=16'd22271;
      117014:data<=16'd24516;
      117015:data<=16'd24156;
      117016:data<=16'd20319;
      117017:data<=16'd19872;
      117018:data<=16'd19834;
      117019:data<=16'd18340;
      117020:data<=16'd21911;
      117021:data<=16'd22777;
      117022:data<=16'd18818;
      117023:data<=16'd21053;
      117024:data<=16'd21798;
      117025:data<=16'd16163;
      117026:data<=16'd16345;
      117027:data<=16'd20879;
      117028:data<=16'd24577;
      117029:data<=16'd28990;
      117030:data<=16'd30039;
      117031:data<=16'd29821;
      117032:data<=16'd31345;
      117033:data<=16'd29431;
      117034:data<=16'd27299;
      117035:data<=16'd28192;
      117036:data<=16'd28289;
      117037:data<=16'd28104;
      117038:data<=16'd26133;
      117039:data<=16'd23168;
      117040:data<=16'd23960;
      117041:data<=16'd23987;
      117042:data<=16'd23111;
      117043:data<=16'd25332;
      117044:data<=16'd24762;
      117045:data<=16'd21872;
      117046:data<=16'd20585;
      117047:data<=16'd18736;
      117048:data<=16'd19023;
      117049:data<=16'd19456;
      117050:data<=16'd17450;
      117051:data<=16'd18022;
      117052:data<=16'd13579;
      117053:data<=16'd1539;
      117054:data<=-16'd3435;
      117055:data<=-16'd2184;
      117056:data<=-16'd2065;
      117057:data<=-16'd1510;
      117058:data<=-16'd2196;
      117059:data<=-16'd2029;
      117060:data<=-16'd1300;
      117061:data<=-16'd3480;
      117062:data<=-16'd1078;
      117063:data<=16'd2426;
      117064:data<=-16'd1292;
      117065:data<=-16'd2560;
      117066:data<=-16'd1011;
      117067:data<=-16'd2444;
      117068:data<=-16'd858;
      117069:data<=16'd751;
      117070:data<=-16'd1309;
      117071:data<=-16'd1343;
      117072:data<=-16'd3;
      117073:data<=16'd637;
      117074:data<=-16'd309;
      117075:data<=-16'd1868;
      117076:data<=-16'd643;
      117077:data<=-16'd2673;
      117078:data<=-16'd8543;
      117079:data<=-16'd9536;
      117080:data<=-16'd9406;
      117081:data<=-16'd11001;
      117082:data<=-16'd10903;
      117083:data<=-16'd12094;
      117084:data<=-16'd12695;
      117085:data<=-16'd10302;
      117086:data<=-16'd9774;
      117087:data<=-16'd10724;
      117088:data<=-16'd11177;
      117089:data<=-16'd13036;
      117090:data<=-16'd14692;
      117091:data<=-16'd12481;
      117092:data<=-16'd10408;
      117093:data<=-16'd12787;
      117094:data<=-16'd8851;
      117095:data<=16'd3142;
      117096:data<=16'd6293;
      117097:data<=16'd3638;
      117098:data<=16'd5372;
      117099:data<=16'd4898;
      117100:data<=16'd4143;
      117101:data<=16'd4834;
      117102:data<=16'd1773;
      117103:data<=16'd1202;
      117104:data<=16'd2137;
      117105:data<=-16'd159;
      117106:data<=16'd761;
      117107:data<=16'd1853;
      117108:data<=-16'd989;
      117109:data<=-16'd2352;
      117110:data<=-16'd2917;
      117111:data<=-16'd3450;
      117112:data<=-16'd2378;
      117113:data<=-16'd2323;
      117114:data<=-16'd3548;
      117115:data<=-16'd3997;
      117116:data<=-16'd3873;
      117117:data<=-16'd4632;
      117118:data<=-16'd5065;
      117119:data<=-16'd4590;
      117120:data<=-16'd5789;
      117121:data<=-16'd5742;
      117122:data<=-16'd4514;
      117123:data<=-16'd6487;
      117124:data<=-16'd6003;
      117125:data<=-16'd4601;
      117126:data<=-16'd7523;
      117127:data<=-16'd5415;
      117128:data<=-16'd155;
      117129:data<=16'd146;
      117130:data<=16'd303;
      117131:data<=16'd161;
      117132:data<=-16'd513;
      117133:data<=-16'd438;
      117134:data<=-16'd1782;
      117135:data<=-16'd614;
      117136:data<=-16'd4690;
      117137:data<=-16'd18067;
      117138:data<=-16'd21855;
      117139:data<=-16'd18301;
      117140:data<=-16'd19358;
      117141:data<=-16'd17656;
      117142:data<=-16'd17349;
      117143:data<=-16'd21238;
      117144:data<=-16'd19784;
      117145:data<=-16'd17896;
      117146:data<=-16'd18117;
      117147:data<=-16'd16137;
      117148:data<=-16'd16043;
      117149:data<=-16'd17180;
      117150:data<=-16'd16763;
      117151:data<=-16'd16051;
      117152:data<=-16'd14598;
      117153:data<=-16'd13847;
      117154:data<=-16'd14481;
      117155:data<=-16'd15242;
      117156:data<=-16'd15515;
      117157:data<=-16'd14898;
      117158:data<=-16'd14713;
      117159:data<=-16'd13585;
      117160:data<=-16'd11982;
      117161:data<=-16'd13600;
      117162:data<=-16'd14266;
      117163:data<=-16'd12540;
      117164:data<=-16'd12584;
      117165:data<=-16'd12392;
      117166:data<=-16'd11694;
      117167:data<=-16'd11359;
      117168:data<=-16'd10989;
      117169:data<=-16'd12276;
      117170:data<=-16'd12041;
      117171:data<=-16'd11036;
      117172:data<=-16'd11869;
      117173:data<=-16'd9624;
      117174:data<=-16'd8050;
      117175:data<=-16'd9159;
      117176:data<=-16'd8768;
      117177:data<=-16'd12957;
      117178:data<=-16'd13990;
      117179:data<=-16'd2963;
      117180:data<=16'd3065;
      117181:data<=16'd2174;
      117182:data<=16'd3797;
      117183:data<=16'd2036;
      117184:data<=16'd1090;
      117185:data<=16'd3724;
      117186:data<=16'd2705;
      117187:data<=16'd3045;
      117188:data<=16'd4654;
      117189:data<=16'd3286;
      117190:data<=16'd4090;
      117191:data<=16'd4607;
      117192:data<=16'd3378;
      117193:data<=16'd4390;
      117194:data<=16'd4629;
      117195:data<=16'd5412;
      117196:data<=16'd7744;
      117197:data<=16'd6513;
      117198:data<=16'd4911;
      117199:data<=16'd5765;
      117200:data<=16'd5961;
      117201:data<=16'd6945;
      117202:data<=16'd9053;
      117203:data<=16'd9512;
      117204:data<=16'd8906;
      117205:data<=16'd8278;
      117206:data<=16'd7511;
      117207:data<=16'd7840;
      117208:data<=16'd9257;
      117209:data<=16'd9265;
      117210:data<=16'd8540;
      117211:data<=16'd8851;
      117212:data<=16'd8537;
      117213:data<=16'd8337;
      117214:data<=16'd8916;
      117215:data<=16'd8849;
      117216:data<=16'd9737;
      117217:data<=16'd9765;
      117218:data<=16'd8786;
      117219:data<=16'd10527;
      117220:data<=16'd6684;
      117221:data<=-16'd4499;
      117222:data<=-16'd8699;
      117223:data<=-16'd6909;
      117224:data<=-16'd7104;
      117225:data<=-16'd6849;
      117226:data<=-16'd6711;
      117227:data<=-16'd4643;
      117228:data<=16'd1709;
      117229:data<=16'd4683;
      117230:data<=16'd4259;
      117231:data<=16'd5971;
      117232:data<=16'd6634;
      117233:data<=16'd5192;
      117234:data<=16'd5081;
      117235:data<=16'd6881;
      117236:data<=16'd8843;
      117237:data<=16'd8473;
      117238:data<=16'd6622;
      117239:data<=16'd6141;
      117240:data<=16'd6764;
      117241:data<=16'd7576;
      117242:data<=16'd8226;
      117243:data<=16'd8008;
      117244:data<=16'd7714;
      117245:data<=16'd8358;
      117246:data<=16'd8513;
      117247:data<=16'd7342;
      117248:data<=16'd7306;
      117249:data<=16'd8766;
      117250:data<=16'd9130;
      117251:data<=16'd8539;
      117252:data<=16'd7971;
      117253:data<=16'd7946;
      117254:data<=16'd8963;
      117255:data<=16'd9330;
      117256:data<=16'd9198;
      117257:data<=16'd8859;
      117258:data<=16'd7242;
      117259:data<=16'd7993;
      117260:data<=16'd8771;
      117261:data<=16'd5130;
      117262:data<=16'd9051;
      117263:data<=16'd22375;
      117264:data<=16'd27269;
      117265:data<=16'd24497;
      117266:data<=16'd24224;
      117267:data<=16'd22683;
      117268:data<=16'd20788;
      117269:data<=16'd22031;
      117270:data<=16'd22109;
      117271:data<=16'd21146;
      117272:data<=16'd20521;
      117273:data<=16'd18704;
      117274:data<=16'd17707;
      117275:data<=16'd18255;
      117276:data<=16'd18234;
      117277:data<=16'd15931;
      117278:data<=16'd10924;
      117279:data<=16'd6775;
      117280:data<=16'd5832;
      117281:data<=16'd6384;
      117282:data<=16'd7420;
      117283:data<=16'd7360;
      117284:data<=16'd6240;
      117285:data<=16'd6354;
      117286:data<=16'd6091;
      117287:data<=16'd4593;
      117288:data<=16'd4332;
      117289:data<=16'd4937;
      117290:data<=16'd4690;
      117291:data<=16'd3469;
      117292:data<=16'd3116;
      117293:data<=16'd4444;
      117294:data<=16'd3673;
      117295:data<=16'd367;
      117296:data<=-16'd811;
      117297:data<=-16'd36;
      117298:data<=-16'd136;
      117299:data<=-16'd449;
      117300:data<=16'd117;
      117301:data<=-16'd441;
      117302:data<=-16'd2617;
      117303:data<=-16'd2437;
      117304:data<=-16'd3764;
      117305:data<=-16'd13317;
      117306:data<=-16'd21138;
      117307:data<=-16'd20262;
      117308:data<=-16'd19931;
      117309:data<=-16'd20870;
      117310:data<=-16'd19338;
      117311:data<=-16'd19024;
      117312:data<=-16'd18712;
      117313:data<=-16'd17790;
      117314:data<=-16'd19214;
      117315:data<=-16'd19523;
      117316:data<=-16'd17772;
      117317:data<=-16'd17420;
      117318:data<=-16'd17509;
      117319:data<=-16'd17277;
      117320:data<=-16'd17170;
      117321:data<=-16'd16286;
      117322:data<=-16'd15838;
      117323:data<=-16'd16527;
      117324:data<=-16'd16120;
      117325:data<=-16'd14965;
      117326:data<=-16'd14966;
      117327:data<=-16'd13749;
      117328:data<=-16'd10125;
      117329:data<=-16'd7567;
      117330:data<=-16'd6484;
      117331:data<=-16'd5974;
      117332:data<=-16'd6740;
      117333:data<=-16'd6451;
      117334:data<=-16'd5589;
      117335:data<=-16'd7518;
      117336:data<=-16'd9309;
      117337:data<=-16'd8405;
      117338:data<=-16'd7087;
      117339:data<=-16'd5999;
      117340:data<=-16'd5090;
      117341:data<=-16'd5655;
      117342:data<=-16'd7947;
      117343:data<=-16'd8963;
      117344:data<=-16'd7459;
      117345:data<=-16'd7653;
      117346:data<=-16'd6173;
      117347:data<=16'd3146;
      117348:data<=16'd10190;
      117349:data<=16'd8607;
      117350:data<=16'd7849;
      117351:data<=16'd8188;
      117352:data<=16'd5633;
      117353:data<=16'd5283;
      117354:data<=16'd6370;
      117355:data<=16'd4874;
      117356:data<=16'd3868;
      117357:data<=16'd4272;
      117358:data<=16'd3849;
      117359:data<=16'd3533;
      117360:data<=16'd4070;
      117361:data<=16'd3254;
      117362:data<=16'd751;
      117363:data<=-16'd44;
      117364:data<=16'd581;
      117365:data<=-16'd255;
      117366:data<=-16'd411;
      117367:data<=16'd337;
      117368:data<=-16'd1075;
      117369:data<=-16'd2403;
      117370:data<=-16'd1757;
      117371:data<=-16'd911;
      117372:data<=-16'd224;
      117373:data<=-16'd44;
      117374:data<=-16'd657;
      117375:data<=-16'd2002;
      117376:data<=-16'd3046;
      117377:data<=-16'd2434;
      117378:data<=-16'd4705;
      117379:data<=-16'd10292;
      117380:data<=-16'd11317;
      117381:data<=-16'd10480;
      117382:data<=-16'd12787;
      117383:data<=-16'd12781;
      117384:data<=-16'd10709;
      117385:data<=-16'd10000;
      117386:data<=-16'd8771;
      117387:data<=-16'd8120;
      117388:data<=-16'd10871;
      117389:data<=-16'd18835;
      117390:data<=-16'd28041;
      117391:data<=-16'd29804;
      117392:data<=-16'd27002;
      117393:data<=-16'd25228;
      117394:data<=-16'd22369;
      117395:data<=-16'd21017;
      117396:data<=-16'd21325;
      117397:data<=-16'd19411;
      117398:data<=-16'd18813;
      117399:data<=-16'd19549;
      117400:data<=-16'd18125;
      117401:data<=-16'd16064;
      117402:data<=-16'd13829;
      117403:data<=-16'd12499;
      117404:data<=-16'd12390;
      117405:data<=-16'd11294;
      117406:data<=-16'd11100;
      117407:data<=-16'd10895;
      117408:data<=-16'd7864;
      117409:data<=-16'd6492;
      117410:data<=-16'd7676;
      117411:data<=-16'd6390;
      117412:data<=-16'd4343;
      117413:data<=-16'd5400;
      117414:data<=-16'd6055;
      117415:data<=-16'd3680;
      117416:data<=-16'd2461;
      117417:data<=-16'd2977;
      117418:data<=-16'd2328;
      117419:data<=-16'd1718;
      117420:data<=-16'd1128;
      117421:data<=16'd176;
      117422:data<=16'd1395;
      117423:data<=16'd2831;
      117424:data<=16'd2974;
      117425:data<=16'd2585;
      117426:data<=16'd2115;
      117427:data<=16'd299;
      117428:data<=16'd4581;
      117429:data<=16'd11903;
      117430:data<=16'd11819;
      117431:data<=16'd17117;
      117432:data<=16'd29037;
      117433:data<=16'd29323;
      117434:data<=16'd26436;
      117435:data<=16'd28976;
      117436:data<=16'd27348;
      117437:data<=16'd25397;
      117438:data<=16'd25711;
      117439:data<=16'd23620;
      117440:data<=16'd23214;
      117441:data<=16'd24362;
      117442:data<=16'd24153;
      117443:data<=16'd23490;
      117444:data<=16'd22010;
      117445:data<=16'd21479;
      117446:data<=16'd21238;
      117447:data<=16'd19896;
      117448:data<=16'd20729;
      117449:data<=16'd21836;
      117450:data<=16'd20128;
      117451:data<=16'd18392;
      117452:data<=16'd17710;
      117453:data<=16'd16537;
      117454:data<=16'd15365;
      117455:data<=16'd16492;
      117456:data<=16'd18218;
      117457:data<=16'd17367;
      117458:data<=16'd16398;
      117459:data<=16'd15960;
      117460:data<=16'd15277;
      117461:data<=16'd15850;
      117462:data<=16'd15085;
      117463:data<=16'd13770;
      117464:data<=16'd14040;
      117465:data<=16'd12417;
      117466:data<=16'd11183;
      117467:data<=16'd11822;
      117468:data<=16'd12057;
      117469:data<=16'd13274;
      117470:data<=16'd12110;
      117471:data<=16'd11186;
      117472:data<=16'd13500;
      117473:data<=16'd6308;
      117474:data<=-16'd5433;
      117475:data<=-16'd6928;
      117476:data<=-16'd6091;
      117477:data<=-16'd5824;
      117478:data<=-16'd5395;
      117479:data<=-16'd10833;
      117480:data<=-16'd12842;
      117481:data<=-16'd9174;
      117482:data<=-16'd9799;
      117483:data<=-16'd10226;
      117484:data<=-16'd8113;
      117485:data<=-16'd7817;
      117486:data<=-16'd8516;
      117487:data<=-16'd9454;
      117488:data<=-16'd7897;
      117489:data<=-16'd5485;
      117490:data<=-16'd6131;
      117491:data<=-16'd5386;
      117492:data<=-16'd3776;
      117493:data<=-16'd4012;
      117494:data<=-16'd2883;
      117495:data<=-16'd1812;
      117496:data<=-16'd1912;
      117497:data<=-16'd1906;
      117498:data<=-16'd2290;
      117499:data<=-16'd2215;
      117500:data<=-16'd2995;
      117501:data<=-16'd3704;
      117502:data<=-16'd2610;
      117503:data<=-16'd3169;
      117504:data<=-16'd3457;
      117505:data<=-16'd2120;
      117506:data<=-16'd2613;
      117507:data<=-16'd3275;
      117508:data<=-16'd4440;
      117509:data<=-16'd5156;
      117510:data<=-16'd3585;
      117511:data<=-16'd4749;
      117512:data<=-16'd5013;
      117513:data<=-16'd3553;
      117514:data<=-16'd6514;
      117515:data<=-16'd1906;
      117516:data<=16'd10328;
      117517:data<=16'd12236;
      117518:data<=16'd10243;
      117519:data<=16'd11761;
      117520:data<=16'd9485;
      117521:data<=16'd7141;
      117522:data<=16'd7065;
      117523:data<=16'd5667;
      117524:data<=16'd4872;
      117525:data<=16'd5027;
      117526:data<=16'd5078;
      117527:data<=16'd4053;
      117528:data<=16'd3732;
      117529:data<=16'd7309;
      117530:data<=16'd9091;
      117531:data<=16'd7109;
      117532:data<=16'd6928;
      117533:data<=16'd6504;
      117534:data<=16'd4237;
      117535:data<=16'd2901;
      117536:data<=16'd2396;
      117537:data<=16'd2300;
      117538:data<=16'd1953;
      117539:data<=16'd2023;
      117540:data<=16'd2030;
      117541:data<=-16'd130;
      117542:data<=-16'd763;
      117543:data<=16'd68;
      117544:data<=-16'd1345;
      117545:data<=-16'd1162;
      117546:data<=16'd296;
      117547:data<=-16'd1008;
      117548:data<=-16'd3021;
      117549:data<=-16'd3588;
      117550:data<=-16'd2328;
      117551:data<=-16'd2419;
      117552:data<=-16'd4077;
      117553:data<=-16'd2717;
      117554:data<=-16'd3786;
      117555:data<=-16'd6684;
      117556:data<=-16'd4011;
      117557:data<=-16'd8434;
      117558:data<=-16'd21391;
      117559:data<=-16'd24013;
      117560:data<=-16'd21161;
      117561:data<=-16'd22682;
      117562:data<=-16'd21687;
      117563:data<=-16'd19728;
      117564:data<=-16'd20491;
      117565:data<=-16'd20149;
      117566:data<=-16'd19129;
      117567:data<=-16'd19052;
      117568:data<=-16'd19678;
      117569:data<=-16'd20371;
      117570:data<=-16'd19543;
      117571:data<=-16'd17590;
      117572:data<=-16'd16187;
      117573:data<=-16'd15938;
      117574:data<=-16'd15878;
      117575:data<=-16'd15543;
      117576:data<=-16'd15274;
      117577:data<=-16'd13973;
      117578:data<=-16'd14104;
      117579:data<=-16'd17547;
      117580:data<=-16'd19402;
      117581:data<=-16'd19773;
      117582:data<=-16'd20707;
      117583:data<=-16'd19240;
      117584:data<=-16'd17801;
      117585:data<=-16'd17465;
      117586:data<=-16'd15403;
      117587:data<=-16'd15133;
      117588:data<=-16'd16595;
      117589:data<=-16'd15967;
      117590:data<=-16'd14775;
      117591:data<=-16'd14114;
      117592:data<=-16'd13808;
      117593:data<=-16'd12659;
      117594:data<=-16'd11409;
      117595:data<=-16'd12809;
      117596:data<=-16'd12117;
      117597:data<=-16'd10646;
      117598:data<=-16'd12871;
      117599:data<=-16'd6270;
      117600:data<=16'd7042;
      117601:data<=16'd8592;
      117602:data<=16'd5577;
      117603:data<=16'd7410;
      117604:data<=16'd7215;
      117605:data<=16'd6766;
      117606:data<=16'd7717;
      117607:data<=16'd7157;
      117608:data<=16'd7213;
      117609:data<=16'd7075;
      117610:data<=16'd6889;
      117611:data<=16'd7738;
      117612:data<=16'd6945;
      117613:data<=16'd6376;
      117614:data<=16'd7303;
      117615:data<=16'd7877;
      117616:data<=16'd8730;
      117617:data<=16'd8288;
      117618:data<=16'd6655;
      117619:data<=16'd6687;
      117620:data<=16'd7345;
      117621:data<=16'd7739;
      117622:data<=16'd8220;
      117623:data<=16'd8909;
      117624:data<=16'd9394;
      117625:data<=16'd8323;
      117626:data<=16'd7559;
      117627:data<=16'd8319;
      117628:data<=16'd10311;
      117629:data<=16'd14270;
      117630:data<=16'd16166;
      117631:data<=16'd15424;
      117632:data<=16'd15696;
      117633:data<=16'd14906;
      117634:data<=16'd14963;
      117635:data<=16'd16271;
      117636:data<=16'd14650;
      117637:data<=16'd14842;
      117638:data<=16'd15107;
      117639:data<=16'd12915;
      117640:data<=16'd15791;
      117641:data<=16'd12898;
      117642:data<=-16'd698;
      117643:data<=-16'd4496;
      117644:data<=-16'd855;
      117645:data<=-16'd2616;
      117646:data<=-16'd2582;
      117647:data<=-16'd212;
      117648:data<=16'd49;
      117649:data<=-16'd50;
      117650:data<=-16'd693;
      117651:data<=-16'd171;
      117652:data<=16'd353;
      117653:data<=-16'd411;
      117654:data<=16'd1494;
      117655:data<=16'd2854;
      117656:data<=16'd1905;
      117657:data<=16'd2857;
      117658:data<=16'd2989;
      117659:data<=16'd2159;
      117660:data<=16'd4044;
      117661:data<=16'd5680;
      117662:data<=16'd5303;
      117663:data<=16'd5066;
      117664:data<=16'd5457;
      117665:data<=16'd5275;
      117666:data<=16'd4604;
      117667:data<=16'd5667;
      117668:data<=16'd7285;
      117669:data<=16'd6883;
      117670:data<=16'd5785;
      117671:data<=16'd5178;
      117672:data<=16'd4895;
      117673:data<=16'd4640;
      117674:data<=16'd5491;
      117675:data<=16'd7250;
      117676:data<=16'd6164;
      117677:data<=16'd5682;
      117678:data<=16'd7297;
      117679:data<=16'd2892;
      117680:data<=-16'd1017;
      117681:data<=16'd1333;
      117682:data<=16'd176;
      117683:data<=16'd3495;
      117684:data<=16'd15829;
      117685:data<=16'd19331;
      117686:data<=16'd17047;
      117687:data<=16'd19155;
      117688:data<=16'd18412;
      117689:data<=16'd16449;
      117690:data<=16'd16672;
      117691:data<=16'd15356;
      117692:data<=16'd14374;
      117693:data<=16'd13835;
      117694:data<=16'd14081;
      117695:data<=16'd15923;
      117696:data<=16'd14748;
      117697:data<=16'd12792;
      117698:data<=16'd13349;
      117699:data<=16'd12885;
      117700:data<=16'd12207;
      117701:data<=16'd12401;
      117702:data<=16'd12038;
      117703:data<=16'd11691;
      117704:data<=16'd10715;
      117705:data<=16'd9740;
      117706:data<=16'd9771;
      117707:data<=16'd9824;
      117708:data<=16'd10430;
      117709:data<=16'd10715;
      117710:data<=16'd9395;
      117711:data<=16'd8126;
      117712:data<=16'd8085;
      117713:data<=16'd8320;
      117714:data<=16'd7260;
      117715:data<=16'd6567;
      117716:data<=16'd7045;
      117717:data<=16'd6047;
      117718:data<=16'd5940;
      117719:data<=16'd6552;
      117720:data<=16'd4226;
      117721:data<=16'd3394;
      117722:data<=16'd3620;
      117723:data<=16'd2598;
      117724:data<=16'd3952;
      117725:data<=-16'd1037;
      117726:data<=-16'd14022;
      117727:data<=-16'd19484;
      117728:data<=-16'd18386;
      117729:data<=-16'd16272;
      117730:data<=-16'd10568;
      117731:data<=-16'd8160;
      117732:data<=-16'd10202;
      117733:data<=-16'd10621;
      117734:data<=-16'd11348;
      117735:data<=-16'd11788;
      117736:data<=-16'd11095;
      117737:data<=-16'd11408;
      117738:data<=-16'd10762;
      117739:data<=-16'd10025;
      117740:data<=-16'd10942;
      117741:data<=-16'd12037;
      117742:data<=-16'd12631;
      117743:data<=-16'd11421;
      117744:data<=-16'd9906;
      117745:data<=-16'd10211;
      117746:data<=-16'd10451;
      117747:data<=-16'd10830;
      117748:data<=-16'd11213;
      117749:data<=-16'd10615;
      117750:data<=-16'd10890;
      117751:data<=-16'd11097;
      117752:data<=-16'd10276;
      117753:data<=-16'd10378;
      117754:data<=-16'd11318;
      117755:data<=-16'd11972;
      117756:data<=-16'd11502;
      117757:data<=-16'd10801;
      117758:data<=-16'd10695;
      117759:data<=-16'd10437;
      117760:data<=-16'd11641;
      117761:data<=-16'd12443;
      117762:data<=-16'd11189;
      117763:data<=-16'd12022;
      117764:data<=-16'd11336;
      117765:data<=-16'd9175;
      117766:data<=-16'd12361;
      117767:data<=-16'd9603;
      117768:data<=16'd2723;
      117769:data<=16'd6998;
      117770:data<=16'd4478;
      117771:data<=16'd5256;
      117772:data<=16'd5128;
      117773:data<=16'd3378;
      117774:data<=16'd2916;
      117775:data<=16'd2960;
      117776:data<=16'd2770;
      117777:data<=16'd2452;
      117778:data<=16'd3130;
      117779:data<=16'd1218;
      117780:data<=-16'd4457;
      117781:data<=-16'd6575;
      117782:data<=-16'd5662;
      117783:data<=-16'd5961;
      117784:data<=-16'd5683;
      117785:data<=-16'd5736;
      117786:data<=-16'd6426;
      117787:data<=-16'd6998;
      117788:data<=-16'd8076;
      117789:data<=-16'd7415;
      117790:data<=-16'd6680;
      117791:data<=-16'd6972;
      117792:data<=-16'd5280;
      117793:data<=-16'd5435;
      117794:data<=-16'd8141;
      117795:data<=-16'd8263;
      117796:data<=-16'd7412;
      117797:data<=-16'd7160;
      117798:data<=-16'd6602;
      117799:data<=-16'd6258;
      117800:data<=-16'd6507;
      117801:data<=-16'd7794;
      117802:data<=-16'd7530;
      117803:data<=-16'd6487;
      117804:data<=-16'd7436;
      117805:data<=-16'd6216;
      117806:data<=-16'd5943;
      117807:data<=-16'd8758;
      117808:data<=-16'd6843;
      117809:data<=-16'd9174;
      117810:data<=-16'd21114;
      117811:data<=-16'd25628;
      117812:data<=-16'd23020;
      117813:data<=-16'd23877;
      117814:data<=-16'd24119;
      117815:data<=-16'd22798;
      117816:data<=-16'd22046;
      117817:data<=-16'd20929;
      117818:data<=-16'd20195;
      117819:data<=-16'd19194;
      117820:data<=-16'd18472;
      117821:data<=-16'd18036;
      117822:data<=-16'd16695;
      117823:data<=-16'd15879;
      117824:data<=-16'd14907;
      117825:data<=-16'd14240;
      117826:data<=-16'd13861;
      117827:data<=-16'd11583;
      117828:data<=-16'd10947;
      117829:data<=-16'd9335;
      117830:data<=-16'd3260;
      117831:data<=-16'd1750;
      117832:data<=-16'd2971;
      117833:data<=-16'd211;
      117834:data<=16'd779;
      117835:data<=16'd864;
      117836:data<=16'd2262;
      117837:data<=16'd1674;
      117838:data<=16'd1726;
      117839:data<=16'd2549;
      117840:data<=16'd2981;
      117841:data<=16'd3665;
      117842:data<=16'd2955;
      117843:data<=16'd3617;
      117844:data<=16'd4686;
      117845:data<=16'd3497;
      117846:data<=16'd4399;
      117847:data<=16'd5236;
      117848:data<=16'd5356;
      117849:data<=16'd7115;
      117850:data<=16'd5489;
      117851:data<=16'd8196;
      117852:data<=16'd20286;
      117853:data<=16'd26078;
      117854:data<=16'd24786;
      117855:data<=16'd25335;
      117856:data<=16'd24359;
      117857:data<=16'd22689;
      117858:data<=16'd22518;
      117859:data<=16'd22028;
      117860:data<=16'd22377;
      117861:data<=16'd22660;
      117862:data<=16'd22316;
      117863:data<=16'd22093;
      117864:data<=16'd21039;
      117865:data<=16'd19887;
      117866:data<=16'd19153;
      117867:data<=16'd19520;
      117868:data<=16'd20350;
      117869:data<=16'd19220;
      117870:data<=16'd18116;
      117871:data<=16'd17556;
      117872:data<=16'd16836;
      117873:data<=16'd17922;
      117874:data<=16'd18086;
      117875:data<=16'd16929;
      117876:data<=16'd16877;
      117877:data<=16'd15869;
      117878:data<=16'd15238;
      117879:data<=16'd14054;
      117880:data<=16'd10219;
      117881:data<=16'd9295;
      117882:data<=16'd9908;
      117883:data<=16'd8962;
      117884:data<=16'd9119;
      117885:data<=16'd7738;
      117886:data<=16'd7215;
      117887:data<=16'd9580;
      117888:data<=16'd8727;
      117889:data<=16'd8040;
      117890:data<=16'd8137;
      117891:data<=16'd5786;
      117892:data<=16'd7353;
      117893:data<=16'd5818;
      117894:data<=-16'd5142;
      117895:data<=-16'd10698;
      117896:data<=-16'd9182;
      117897:data<=-16'd9574;
      117898:data<=-16'd9612;
      117899:data<=-16'd8731;
      117900:data<=-16'd7791;
      117901:data<=-16'd6631;
      117902:data<=-16'd7054;
      117903:data<=-16'd7050;
      117904:data<=-16'd6786;
      117905:data<=-16'd7456;
      117906:data<=-16'd6172;
      117907:data<=-16'd4366;
      117908:data<=-16'd4308;
      117909:data<=-16'd4405;
      117910:data<=-16'd4200;
      117911:data<=-16'd3908;
      117912:data<=-16'd3483;
      117913:data<=-16'd2199;
      117914:data<=-16'd960;
      117915:data<=-16'd1642;
      117916:data<=-16'd1348;
      117917:data<=-16'd9;
      117918:data<=-16'd992;
      117919:data<=-16'd1162;
      117920:data<=16'd711;
      117921:data<=16'd1160;
      117922:data<=16'd535;
      117923:data<=16'd331;
      117924:data<=16'd651;
      117925:data<=16'd560;
      117926:data<=16'd156;
      117927:data<=16'd52;
      117928:data<=-16'd1462;
      117929:data<=-16'd214;
      117930:data<=16'd5644;
      117931:data<=16'd6878;
      117932:data<=16'd5089;
      117933:data<=16'd5125;
      117934:data<=16'd1848;
      117935:data<=16'd3479;
      117936:data<=16'd14747;
      117937:data<=16'd20378;
      117938:data<=16'd19308;
      117939:data<=16'd19068;
      117940:data<=16'd16654;
      117941:data<=16'd14463;
      117942:data<=16'd14803;
      117943:data<=16'd13905;
      117944:data<=16'd13104;
      117945:data<=16'd12930;
      117946:data<=16'd11388;
      117947:data<=16'd9535;
      117948:data<=16'd8417;
      117949:data<=16'd7888;
      117950:data<=16'd7380;
      117951:data<=16'd7491;
      117952:data<=16'd7597;
      117953:data<=16'd5319;
      117954:data<=16'd3424;
      117955:data<=16'd3477;
      117956:data<=16'd2505;
      117957:data<=16'd2428;
      117958:data<=16'd3392;
      117959:data<=16'd1738;
      117960:data<=-16'd347;
      117961:data<=-16'd975;
      117962:data<=-16'd1671;
      117963:data<=-16'd1996;
      117964:data<=-16'd1422;
      117965:data<=-16'd1162;
      117966:data<=-16'd2693;
      117967:data<=-16'd4203;
      117968:data<=-16'd3676;
      117969:data<=-16'd3715;
      117970:data<=-16'd4131;
      117971:data<=-16'd3595;
      117972:data<=-16'd4573;
      117973:data<=-16'd5976;
      117974:data<=-16'd6828;
      117975:data<=-16'd7277;
      117976:data<=-16'd5260;
      117977:data<=-16'd6661;
      117978:data<=-16'd15529;
      117979:data<=-16'd23928;
      117980:data<=-16'd29040;
      117981:data<=-16'd31907;
      117982:data<=-16'd30702;
      117983:data<=-16'd28744;
      117984:data<=-16'd27924;
      117985:data<=-16'd26861;
      117986:data<=-16'd27132;
      117987:data<=-16'd27604;
      117988:data<=-16'd26617;
      117989:data<=-16'd25539;
      117990:data<=-16'd24186;
      117991:data<=-16'd22651;
      117992:data<=-16'd22260;
      117993:data<=-16'd23302;
      117994:data<=-16'd24071;
      117995:data<=-16'd22563;
      117996:data<=-16'd20773;
      117997:data<=-16'd19916;
      117998:data<=-16'd18418;
      117999:data<=-16'd18271;
      118000:data<=-16'd19749;
      118001:data<=-16'd19657;
      118002:data<=-16'd18434;
      118003:data<=-16'd17014;
      118004:data<=-16'd15449;
      118005:data<=-16'd14918;
      118006:data<=-16'd15494;
      118007:data<=-16'd16427;
      118008:data<=-16'd15993;
      118009:data<=-16'd14424;
      118010:data<=-16'd14028;
      118011:data<=-16'd13227;
      118012:data<=-16'd12234;
      118013:data<=-16'd13365;
      118014:data<=-16'd13588;
      118015:data<=-16'd12659;
      118016:data<=-16'd12120;
      118017:data<=-16'd10328;
      118018:data<=-16'd10404;
      118019:data<=-16'd10097;
      118020:data<=-16'd1697;
      118021:data<=16'd7072;
      118022:data<=16'd7862;
      118023:data<=16'd7145;
      118024:data<=16'd7812;
      118025:data<=16'd7292;
      118026:data<=16'd6376;
      118027:data<=16'd5394;
      118028:data<=16'd4772;
      118029:data<=16'd5944;
      118030:data<=16'd8947;
      118031:data<=16'd11850;
      118032:data<=16'd12146;
      118033:data<=16'd10866;
      118034:data<=16'd9999;
      118035:data<=16'd9412;
      118036:data<=16'd9890;
      118037:data<=16'd10624;
      118038:data<=16'd10225;
      118039:data<=16'd10313;
      118040:data<=16'd10596;
      118041:data<=16'd10417;
      118042:data<=16'd10965;
      118043:data<=16'd10901;
      118044:data<=16'd9975;
      118045:data<=16'd10116;
      118046:data<=16'd10836;
      118047:data<=16'd11166;
      118048:data<=16'd11098;
      118049:data<=16'd10986;
      118050:data<=16'd10916;
      118051:data<=16'd10554;
      118052:data<=16'd11033;
      118053:data<=16'd12038;
      118054:data<=16'd11884;
      118055:data<=16'd11635;
      118056:data<=16'd11605;
      118057:data<=16'd11247;
      118058:data<=16'd10850;
      118059:data<=16'd10425;
      118060:data<=16'd12107;
      118061:data<=16'd12225;
      118062:data<=16'd3230;
      118063:data<=-16'd6966;
      118064:data<=-16'd8081;
      118065:data<=-16'd5591;
      118066:data<=-16'd4149;
      118067:data<=-16'd2996;
      118068:data<=-16'd3040;
      118069:data<=-16'd2822;
      118070:data<=-16'd2549;
      118071:data<=-16'd3435;
      118072:data<=-16'd2441;
      118073:data<=-16'd224;
      118074:data<=-16'd79;
      118075:data<=-16'd293;
      118076:data<=16'd406;
      118077:data<=16'd350;
      118078:data<=16'd563;
      118079:data<=16'd2184;
      118080:data<=16'd1368;
      118081:data<=-16'd2338;
      118082:data<=-16'd3036;
      118083:data<=-16'd1726;
      118084:data<=-16'd2544;
      118085:data<=-16'd2085;
      118086:data<=16'd365;
      118087:data<=16'd1204;
      118088:data<=16'd1071;
      118089:data<=16'd1186;
      118090:data<=16'd1398;
      118091:data<=16'd1434;
      118092:data<=16'd1935;
      118093:data<=16'd4032;
      118094:data<=16'd4687;
      118095:data<=16'd3309;
      118096:data<=16'd3530;
      118097:data<=16'd3662;
      118098:data<=16'd3635;
      118099:data<=16'd5113;
      118100:data<=16'd4945;
      118101:data<=16'd4725;
      118102:data<=16'd5096;
      118103:data<=16'd4592;
      118104:data<=16'd11035;
      118105:data<=16'd21971;
      118106:data<=16'd24811;
      118107:data<=16'd23193;
      118108:data<=16'd23056;
      118109:data<=16'd21893;
      118110:data<=16'd20744;
      118111:data<=16'd20028;
      118112:data<=16'd20111;
      118113:data<=16'd21849;
      118114:data<=16'd21291;
      118115:data<=16'd19243;
      118116:data<=16'd19139;
      118117:data<=16'd18430;
      118118:data<=16'd17011;
      118119:data<=16'd17111;
      118120:data<=16'd17227;
      118121:data<=16'd16571;
      118122:data<=16'd16318;
      118123:data<=16'd15932;
      118124:data<=16'd14580;
      118125:data<=16'd14222;
      118126:data<=16'd15239;
      118127:data<=16'd15111;
      118128:data<=16'd13925;
      118129:data<=16'd12665;
      118130:data<=16'd13449;
      118131:data<=16'd17546;
      118132:data<=16'd19136;
      118133:data<=16'd17644;
      118134:data<=16'd17939;
      118135:data<=16'd17015;
      118136:data<=16'd15650;
      118137:data<=16'd16524;
      118138:data<=16'd15123;
      118139:data<=16'd13600;
      118140:data<=16'd13864;
      118141:data<=16'd12815;
      118142:data<=16'd12627;
      118143:data<=16'd11423;
      118144:data<=16'd10008;
      118145:data<=16'd11409;
      118146:data<=16'd4238;
      118147:data<=-16'd9033;
      118148:data<=-16'd11809;
      118149:data<=-16'd10191;
      118150:data<=-16'd11247;
      118151:data<=-16'd9903;
      118152:data<=-16'd9931;
      118153:data<=-16'd12184;
      118154:data<=-16'd12389;
      118155:data<=-16'd12320;
      118156:data<=-16'd11732;
      118157:data<=-16'd10786;
      118158:data<=-16'd11931;
      118159:data<=-16'd13100;
      118160:data<=-16'd12622;
      118161:data<=-16'd11879;
      118162:data<=-16'd11994;
      118163:data<=-16'd12082;
      118164:data<=-16'd11006;
      118165:data<=-16'd10813;
      118166:data<=-16'd11978;
      118167:data<=-16'd12323;
      118168:data<=-16'd12314;
      118169:data<=-16'd12246;
      118170:data<=-16'd11321;
      118171:data<=-16'd10598;
      118172:data<=-16'd11307;
      118173:data<=-16'd12613;
      118174:data<=-16'd12725;
      118175:data<=-16'd12220;
      118176:data<=-16'd11626;
      118177:data<=-16'd10648;
      118178:data<=-16'd11215;
      118179:data<=-16'd12208;
      118180:data<=-16'd13432;
      118181:data<=-16'd17810;
      118182:data<=-16'd19406;
      118183:data<=-16'd16750;
      118184:data<=-16'd17387;
      118185:data<=-16'd17481;
      118186:data<=-16'd16986;
      118187:data<=-16'd20086;
      118188:data<=-16'd13958;
      118189:data<=-16'd94;
      118190:data<=16'd3298;
      118191:data<=16'd911;
      118192:data<=16'd1198;
      118193:data<=-16'd247;
      118194:data<=-16'd1287;
      118195:data<=-16'd544;
      118196:data<=-16'd660;
      118197:data<=-16'd256;
      118198:data<=-16'd564;
      118199:data<=-16'd2091;
      118200:data<=-16'd2469;
      118201:data<=-16'd2872;
      118202:data<=-16'd3755;
      118203:data<=-16'd3539;
      118204:data<=-16'd2702;
      118205:data<=-16'd3065;
      118206:data<=-16'd4764;
      118207:data<=-16'd5466;
      118208:data<=-16'd5204;
      118209:data<=-16'd5140;
      118210:data<=-16'd4276;
      118211:data<=-16'd4311;
      118212:data<=-16'd5850;
      118213:data<=-16'd5918;
      118214:data<=-16'd5394;
      118215:data<=-16'd5512;
      118216:data<=-16'd5289;
      118217:data<=-16'd5280;
      118218:data<=-16'd5468;
      118219:data<=-16'd6184;
      118220:data<=-16'd7227;
      118221:data<=-16'd6799;
      118222:data<=-16'd6072;
      118223:data<=-16'd5550;
      118224:data<=-16'd4663;
      118225:data<=-16'd5260;
      118226:data<=-16'd6543;
      118227:data<=-16'd7104;
      118228:data<=-16'd6516;
      118229:data<=-16'd5027;
      118230:data<=-16'd8472;
      118231:data<=-16'd16067;
      118232:data<=-16'd18697;
      118233:data<=-16'd17993;
      118234:data<=-16'd18195;
      118235:data<=-16'd17337;
      118236:data<=-16'd16736;
      118237:data<=-16'd16413;
      118238:data<=-16'd15659;
      118239:data<=-16'd16402;
      118240:data<=-16'd16389;
      118241:data<=-16'd15091;
      118242:data<=-16'd14645;
      118243:data<=-16'd13816;
      118244:data<=-16'd12895;
      118245:data<=-16'd12034;
      118246:data<=-16'd11003;
      118247:data<=-16'd11358;
      118248:data<=-16'd11071;
      118249:data<=-16'd9922;
      118250:data<=-16'd9781;
      118251:data<=-16'd7947;
      118252:data<=-16'd5492;
      118253:data<=-16'd5474;
      118254:data<=-16'd5465;
      118255:data<=-16'd4579;
      118256:data<=-16'd4056;
      118257:data<=-16'd3570;
      118258:data<=-16'd2549;
      118259:data<=-16'd1475;
      118260:data<=-16'd1651;
      118261:data<=-16'd1524;
      118262:data<=-16'd628;
      118263:data<=-16'd1356;
      118264:data<=-16'd1703;
      118265:data<=-16'd526;
      118266:data<=16'd743;
      118267:data<=16'd2015;
      118268:data<=16'd1295;
      118269:data<=16'd1002;
      118270:data<=16'd1983;
      118271:data<=16'd334;
      118272:data<=16'd5958;
      118273:data<=16'd19732;
      118274:data<=16'd22759;
      118275:data<=16'd19139;
      118276:data<=16'd20721;
      118277:data<=16'd19660;
      118278:data<=16'd18131;
      118279:data<=16'd21259;
      118280:data<=16'd20177;
      118281:data<=16'd15223;
      118282:data<=16'd13029;
      118283:data<=16'd12524;
      118284:data<=16'd12208;
      118285:data<=16'd12448;
      118286:data<=16'd12991;
      118287:data<=16'd12398;
      118288:data<=16'd11230;
      118289:data<=16'd11411;
      118290:data<=16'd11112;
      118291:data<=16'd10583;
      118292:data<=16'd11508;
      118293:data<=16'd11634;
      118294:data<=16'd11220;
      118295:data<=16'd11144;
      118296:data<=16'd10255;
      118297:data<=16'd9691;
      118298:data<=16'd10040;
      118299:data<=16'd11148;
      118300:data<=16'd11808;
      118301:data<=16'd10460;
      118302:data<=16'd9580;
      118303:data<=16'd9623;
      118304:data<=16'd9737;
      118305:data<=16'd11192;
      118306:data<=16'd11614;
      118307:data<=16'd10662;
      118308:data<=16'd9885;
      118309:data<=16'd8790;
      118310:data<=16'd9532;
      118311:data<=16'd9690;
      118312:data<=16'd9210;
      118313:data<=16'd12245;
      118314:data<=16'd7501;
      118315:data<=-16'd5984;
      118316:data<=-16'd10108;
      118317:data<=-16'd8267;
      118318:data<=-16'd8677;
      118319:data<=-16'd6344;
      118320:data<=-16'd5718;
      118321:data<=-16'd7200;
      118322:data<=-16'd5730;
      118323:data<=-16'd5874;
      118324:data<=-16'd5926;
      118325:data<=-16'd3506;
      118326:data<=-16'd3210;
      118327:data<=-16'd3046;
      118328:data<=-16'd2197;
      118329:data<=-16'd2507;
      118330:data<=-16'd943;
      118331:data<=16'd2664;
      118332:data<=16'd5943;
      118333:data<=16'd7341;
      118334:data<=16'd6717;
      118335:data<=16'd6357;
      118336:data<=16'd5915;
      118337:data<=16'd5134;
      118338:data<=16'd6028;
      118339:data<=16'd7415;
      118340:data<=16'd7363;
      118341:data<=16'd6281;
      118342:data<=16'd6093;
      118343:data<=16'd6516;
      118344:data<=16'd5482;
      118345:data<=16'd5694;
      118346:data<=16'd7039;
      118347:data<=16'd5820;
      118348:data<=16'd5034;
      118349:data<=16'd5274;
      118350:data<=16'd4949;
      118351:data<=16'd5750;
      118352:data<=16'd5269;
      118353:data<=16'd5163;
      118354:data<=16'd5888;
      118355:data<=16'd2646;
      118356:data<=16'd6660;
      118357:data<=16'd20272;
      118358:data<=16'd23394;
      118359:data<=16'd18393;
      118360:data<=16'd18048;
      118361:data<=16'd16856;
      118362:data<=16'd14938;
      118363:data<=16'd15377;
      118364:data<=16'd13521;
      118365:data<=16'd11069;
      118366:data<=16'd10560;
      118367:data<=16'd9837;
      118368:data<=16'd8599;
      118369:data<=16'd7746;
      118370:data<=16'd7244;
      118371:data<=16'd5344;
      118372:data<=16'd3136;
      118373:data<=16'd3030;
      118374:data<=16'd2331;
      118375:data<=16'd1196;
      118376:data<=16'd2105;
      118377:data<=16'd2281;
      118378:data<=16'd905;
      118379:data<=-16'd209;
      118380:data<=-16'd1833;
      118381:data<=-16'd4937;
      118382:data<=-16'd7943;
      118383:data<=-16'd8084;
      118384:data<=-16'd7679;
      118385:data<=-16'd9374;
      118386:data<=-16'd9671;
      118387:data<=-16'd8783;
      118388:data<=-16'd8913;
      118389:data<=-16'd8560;
      118390:data<=-16'd8539;
      118391:data<=-16'd9078;
      118392:data<=-16'd10273;
      118393:data<=-16'd11919;
      118394:data<=-16'd10707;
      118395:data<=-16'd10267;
      118396:data<=-16'd11079;
      118397:data<=-16'd8345;
      118398:data<=-16'd13077;
      118399:data<=-16'd26435;
      118400:data<=-16'd30198;
      118401:data<=-16'd27200;
      118402:data<=-16'd27577;
      118403:data<=-16'd26715;
      118404:data<=-16'd25713;
      118405:data<=-16'd26409;
      118406:data<=-16'd25542;
      118407:data<=-16'd24923;
      118408:data<=-16'd24674;
      118409:data<=-16'd23491;
      118410:data<=-16'd22430;
      118411:data<=-16'd21594;
      118412:data<=-16'd21584;
      118413:data<=-16'd20996;
      118414:data<=-16'd19183;
      118415:data<=-16'd18719;
      118416:data<=-16'd18283;
      118417:data<=-16'd17224;
      118418:data<=-16'd17811;
      118419:data<=-16'd18340;
      118420:data<=-16'd17302;
      118421:data<=-16'd16195;
      118422:data<=-16'd15696;
      118423:data<=-16'd14959;
      118424:data<=-16'd14142;
      118425:data<=-16'd14804;
      118426:data<=-16'd15229;
      118427:data<=-16'd14295;
      118428:data<=-16'd14448;
      118429:data<=-16'd14173;
      118430:data<=-16'd12380;
      118431:data<=-16'd10469;
      118432:data<=-16'd7683;
      118433:data<=-16'd6220;
      118434:data<=-16'd6015;
      118435:data<=-16'd4993;
      118436:data<=-16'd5850;
      118437:data<=-16'd5580;
      118438:data<=-16'd4540;
      118439:data<=-16'd7783;
      118440:data<=-16'd3674;
      118441:data<=16'd9571;
      118442:data<=16'd14316;
      118443:data<=16'd12601;
      118444:data<=16'd12777;
      118445:data<=16'd10936;
      118446:data<=16'd9670;
      118447:data<=16'd10266;
      118448:data<=16'd9338;
      118449:data<=16'd9094;
      118450:data<=16'd8901;
      118451:data<=16'd7629;
      118452:data<=16'd7235;
      118453:data<=16'd6930;
      118454:data<=16'd6534;
      118455:data<=16'd5876;
      118456:data<=16'd4884;
      118457:data<=16'd5271;
      118458:data<=16'd5632;
      118459:data<=16'd5112;
      118460:data<=16'd5109;
      118461:data<=16'd5248;
      118462:data<=16'd5422;
      118463:data<=16'd5257;
      118464:data<=16'd5310;
      118465:data<=16'd6936;
      118466:data<=16'd7815;
      118467:data<=16'd7429;
      118468:data<=16'd7808;
      118469:data<=16'd7837;
      118470:data<=16'd7024;
      118471:data<=16'd7043;
      118472:data<=16'd8390;
      118473:data<=16'd9098;
      118474:data<=16'd8272;
      118475:data<=16'd8084;
      118476:data<=16'd7709;
      118477:data<=16'd7665;
      118478:data<=16'd10396;
      118479:data<=16'd10587;
      118480:data<=16'd8898;
      118481:data<=16'd9166;
      118482:data<=16'd961;
      118483:data<=-16'd13089;
      118484:data<=-16'd16424;
      118485:data<=-16'd13224;
      118486:data<=-16'd11979;
      118487:data<=-16'd10756;
      118488:data<=-16'd10786;
      118489:data<=-16'd11019;
      118490:data<=-16'd9673;
      118491:data<=-16'd8461;
      118492:data<=-16'd6648;
      118493:data<=-16'd5947;
      118494:data<=-16'd6878;
      118495:data<=-16'd6125;
      118496:data<=-16'd5025;
      118497:data<=-16'd4162;
      118498:data<=-16'd2181;
      118499:data<=-16'd1017;
      118500:data<=-16'd855;
      118501:data<=-16'd485;
      118502:data<=-16'd247;
      118503:data<=-16'd664;
      118504:data<=-16'd937;
      118505:data<=16'd622;
      118506:data<=16'd1968;
      118507:data<=16'd1644;
      118508:data<=16'd1941;
      118509:data<=16'd1929;
      118510:data<=16'd1811;
      118511:data<=16'd3404;
      118512:data<=16'd4376;
      118513:data<=16'd4868;
      118514:data<=16'd5360;
      118515:data<=16'd4408;
      118516:data<=16'd4314;
      118517:data<=16'd5294;
      118518:data<=16'd6351;
      118519:data<=16'd7409;
      118520:data<=16'd6396;
      118521:data<=16'd6610;
      118522:data<=16'd7849;
      118523:data<=16'd5248;
      118524:data<=16'd8843;
      118525:data<=16'd21843;
      118526:data<=16'd27472;
      118527:data<=16'd24413;
      118528:data<=16'd23513;
      118529:data<=16'd23109;
      118530:data<=16'd21937;
      118531:data<=16'd24515;
      118532:data<=16'd28749;
      118533:data<=16'd29244;
      118534:data<=16'd27284;
      118535:data<=16'd26730;
      118536:data<=16'd26231;
      118537:data<=16'd25176;
      118538:data<=16'd25373;
      118539:data<=16'd25100;
      118540:data<=16'd23887;
      118541:data<=16'd22821;
      118542:data<=16'd21212;
      118543:data<=16'd20503;
      118544:data<=16'd21082;
      118545:data<=16'd21455;
      118546:data<=16'd21557;
      118547:data<=16'd20416;
      118548:data<=16'd18918;
      118549:data<=16'd18462;
      118550:data<=16'd17682;
      118551:data<=16'd17447;
      118552:data<=16'd17757;
      118553:data<=16'd17130;
      118554:data<=16'd16688;
      118555:data<=16'd15509;
      118556:data<=16'd14022;
      118557:data<=16'd14390;
      118558:data<=16'd14419;
      118559:data<=16'd14069;
      118560:data<=16'd13761;
      118561:data<=16'd12116;
      118562:data<=16'd11800;
      118563:data<=16'd11215;
      118564:data<=16'd9194;
      118565:data<=16'd10219;
      118566:data<=16'd7056;
      118567:data<=-16'd4469;
      118568:data<=-16'd10754;
      118569:data<=-16'd9365;
      118570:data<=-16'd9388;
      118571:data<=-16'd10784;
      118572:data<=-16'd11788;
      118573:data<=-16'd12020;
      118574:data<=-16'd11265;
      118575:data<=-16'd11876;
      118576:data<=-16'd12013;
      118577:data<=-16'd10959;
      118578:data<=-16'd12857;
      118579:data<=-16'd14205;
      118580:data<=-16'd11732;
      118581:data<=-16'd12692;
      118582:data<=-16'd17261;
      118583:data<=-16'd17681;
      118584:data<=-16'd16782;
      118585:data<=-16'd18651;
      118586:data<=-16'd18759;
      118587:data<=-16'd17576;
      118588:data<=-16'd17769;
      118589:data<=-16'd16891;
      118590:data<=-16'd16747;
      118591:data<=-16'd18342;
      118592:data<=-16'd17911;
      118593:data<=-16'd17179;
      118594:data<=-16'd17505;
      118595:data<=-16'd16671;
      118596:data<=-16'd15952;
      118597:data<=-16'd15571;
      118598:data<=-16'd15432;
      118599:data<=-16'd16569;
      118600:data<=-16'd16581;
      118601:data<=-16'd15506;
      118602:data<=-16'd14694;
      118603:data<=-16'd13502;
      118604:data<=-16'd14151;
      118605:data<=-16'd14886;
      118606:data<=-16'd13671;
      118607:data<=-16'd14680;
      118608:data<=-16'd12057;
      118609:data<=-16'd781;
      118610:data<=16'd5950;
      118611:data<=16'd3755;
      118612:data<=16'd2620;
      118613:data<=16'd3247;
      118614:data<=16'd2927;
      118615:data<=16'd3036;
      118616:data<=16'd2936;
      118617:data<=16'd2215;
      118618:data<=16'd843;
      118619:data<=-16'd511;
      118620:data<=16'd111;
      118621:data<=16'd790;
      118622:data<=16'd17;
      118623:data<=-16'd214;
      118624:data<=-16'd717;
      118625:data<=-16'd2141;
      118626:data<=-16'd2678;
      118627:data<=-16'd2713;
      118628:data<=-16'd2356;
      118629:data<=-16'd1624;
      118630:data<=-16'd2484;
      118631:data<=-16'd2652;
      118632:data<=16'd719;
      118633:data<=16'd3048;
      118634:data<=16'd2217;
      118635:data<=16'd2554;
      118636:data<=16'd3521;
      118637:data<=16'd2303;
      118638:data<=16'd647;
      118639:data<=-16'd397;
      118640:data<=-16'd719;
      118641:data<=-16'd11;
      118642:data<=16'd77;
      118643:data<=-16'd429;
      118644:data<=-16'd1522;
      118645:data<=-16'd3615;
      118646:data<=-16'd3413;
      118647:data<=-16'd2516;
      118648:data<=-16'd3859;
      118649:data<=-16'd2457;
      118650:data<=-16'd3196;
      118651:data<=-16'd14413;
      118652:data<=-16'd23450;
      118653:data<=-16'd22146;
      118654:data<=-16'd20947;
      118655:data<=-16'd20961;
      118656:data<=-16'd18671;
      118657:data<=-16'd18677;
      118658:data<=-16'd19923;
      118659:data<=-16'd19227;
      118660:data<=-16'd18691;
      118661:data<=-16'd18102;
      118662:data<=-16'd17139;
      118663:data<=-16'd17127;
      118664:data<=-16'd17006;
      118665:data<=-16'd16584;
      118666:data<=-16'd16550;
      118667:data<=-16'd15790;
      118668:data<=-16'd14481;
      118669:data<=-16'd13967;
      118670:data<=-16'd13512;
      118671:data<=-16'd12384;
      118672:data<=-16'd11861;
      118673:data<=-16'd11637;
      118674:data<=-16'd10439;
      118675:data<=-16'd9994;
      118676:data<=-16'd10355;
      118677:data<=-16'd8801;
      118678:data<=-16'd6799;
      118679:data<=-16'd6141;
      118680:data<=-16'd5016;
      118681:data<=-16'd5087;
      118682:data<=-16'd8677;
      118683:data<=-16'd11138;
      118684:data<=-16'd9004;
      118685:data<=-16'd6807;
      118686:data<=-16'd6837;
      118687:data<=-16'd5974;
      118688:data<=-16'd5339;
      118689:data<=-16'd5567;
      118690:data<=-16'd3388;
      118691:data<=-16'd2023;
      118692:data<=-16'd848;
      118693:data<=16'd8244;
      118694:data<=16'd17661;
      118695:data<=16'd17203;
      118696:data<=16'd15403;
      118697:data<=16'd16815;
      118698:data<=16'd16819;
      118699:data<=16'd16732;
      118700:data<=16'd16903;
      118701:data<=16'd16219;
      118702:data<=16'd16051;
      118703:data<=16'd16234;
      118704:data<=16'd17399;
      118705:data<=16'd18161;
      118706:data<=16'd16352;
      118707:data<=16'd15456;
      118708:data<=16'd15713;
      118709:data<=16'd14358;
      118710:data<=16'd13916;
      118711:data<=16'd15029;
      118712:data<=16'd15417;
      118713:data<=16'd15289;
      118714:data<=16'd14856;
      118715:data<=16'd13826;
      118716:data<=16'd12938;
      118717:data<=16'd13493;
      118718:data<=16'd14586;
      118719:data<=16'd14082;
      118720:data<=16'd13638;
      118721:data<=16'd13850;
      118722:data<=16'd12938;
      118723:data<=16'd12825;
      118724:data<=16'd13949;
      118725:data<=16'd14374;
      118726:data<=16'd14277;
      118727:data<=16'd13382;
      118728:data<=16'd12487;
      118729:data<=16'd12022;
      118730:data<=16'd11382;
      118731:data<=16'd12856;
      118732:data<=16'd15559;
      118733:data<=16'd17559;
      118734:data<=16'd17468;
      118735:data<=16'd8940;
      118736:data<=-16'd2003;
      118737:data<=-16'd2311;
      118738:data<=16'd661;
      118739:data<=-16'd214;
      118740:data<=16'd928;
      118741:data<=16'd1677;
      118742:data<=-16'd76;
      118743:data<=16'd347;
      118744:data<=16'd1651;
      118745:data<=16'd1579;
      118746:data<=16'd1052;
      118747:data<=16'd893;
      118748:data<=16'd1304;
      118749:data<=16'd1451;
      118750:data<=16'd2466;
      118751:data<=16'd4067;
      118752:data<=16'd3686;
      118753:data<=16'd3087;
      118754:data<=16'd3228;
      118755:data<=16'd2713;
      118756:data<=16'd2983;
      118757:data<=16'd4149;
      118758:data<=16'd4749;
      118759:data<=16'd4488;
      118760:data<=16'd3965;
      118761:data<=16'd3993;
      118762:data<=16'd3181;
      118763:data<=16'd2575;
      118764:data<=16'd4407;
      118765:data<=16'd5068;
      118766:data<=16'd3698;
      118767:data<=16'd3234;
      118768:data<=16'd3019;
      118769:data<=16'd3183;
      118770:data<=16'd3745;
      118771:data<=16'd3958;
      118772:data<=16'd4134;
      118773:data<=16'd3445;
      118774:data<=16'd4084;
      118775:data<=16'd4645;
      118776:data<=16'd2475;
      118777:data<=16'd8220;
      118778:data<=16'd20266;
      118779:data<=16'd21484;
      118780:data<=16'd17700;
      118781:data<=16'd18101;
      118782:data<=16'd14478;
      118783:data<=16'd9072;
      118784:data<=16'd7662;
      118785:data<=16'd6572;
      118786:data<=16'd6149;
      118787:data<=16'd6384;
      118788:data<=16'd5674;
      118789:data<=16'd5335;
      118790:data<=16'd3580;
      118791:data<=16'd734;
      118792:data<=16'd124;
      118793:data<=16'd346;
      118794:data<=-16'd27;
      118795:data<=-16'd9;
      118796:data<=-16'd564;
      118797:data<=-16'd2335;
      118798:data<=-16'd3168;
      118799:data<=-16'd3042;
      118800:data<=-16'd3892;
      118801:data<=-16'd3548;
      118802:data<=-16'd2220;
      118803:data<=-16'd3542;
      118804:data<=-16'd4813;
      118805:data<=-16'd4845;
      118806:data<=-16'd5873;
      118807:data<=-16'd5598;
      118808:data<=-16'd4872;
      118809:data<=-16'd5163;
      118810:data<=-16'd5269;
      118811:data<=-16'd7050;
      118812:data<=-16'd7861;
      118813:data<=-16'd7009;
      118814:data<=-16'd8522;
      118815:data<=-16'd8257;
      118816:data<=-16'd7650;
      118817:data<=-16'd9574;
      118818:data<=-16'd8200;
      118819:data<=-16'd12756;
      118820:data<=-16'd25680;
      118821:data<=-16'd27931;
      118822:data<=-16'd23293;
      118823:data<=-16'd24004;
      118824:data<=-16'd23845;
      118825:data<=-16'd23052;
      118826:data<=-16'd23278;
      118827:data<=-16'd21957;
      118828:data<=-16'd22368;
      118829:data<=-16'd22087;
      118830:data<=-16'd21058;
      118831:data<=-16'd22789;
      118832:data<=-16'd20102;
      118833:data<=-16'd13873;
      118834:data<=-16'd12408;
      118835:data<=-16'd12466;
      118836:data<=-16'd11922;
      118837:data<=-16'd12486;
      118838:data<=-16'd11699;
      118839:data<=-16'd9953;
      118840:data<=-16'd9415;
      118841:data<=-16'd9288;
      118842:data<=-16'd9077;
      118843:data<=-16'd9784;
      118844:data<=-16'd10768;
      118845:data<=-16'd10381;
      118846:data<=-16'd9997;
      118847:data<=-16'd9746;
      118848:data<=-16'd8287;
      118849:data<=-16'd8123;
      118850:data<=-16'd9291;
      118851:data<=-16'd9717;
      118852:data<=-16'd9834;
      118853:data<=-16'd9159;
      118854:data<=-16'd8968;
      118855:data<=-16'd9001;
      118856:data<=-16'd7949;
      118857:data<=-16'd9444;
      118858:data<=-16'd9976;
      118859:data<=-16'd7929;
      118860:data<=-16'd9996;
      118861:data<=-16'd5924;
      118862:data<=16'd7357;
      118863:data<=16'd9955;
      118864:data<=16'd5096;
      118865:data<=16'd5906;
      118866:data<=16'd5538;
      118867:data<=16'd4302;
      118868:data<=16'd5990;
      118869:data<=16'd5776;
      118870:data<=16'd4843;
      118871:data<=16'd4220;
      118872:data<=16'd3351;
      118873:data<=16'd3650;
      118874:data<=16'd2840;
      118875:data<=16'd2088;
      118876:data<=16'd2420;
      118877:data<=16'd1337;
      118878:data<=16'd1391;
      118879:data<=16'd1930;
      118880:data<=16'd983;
      118881:data<=16'd1595;
      118882:data<=16'd422;
      118883:data<=-16'd4111;
      118884:data<=-16'd5433;
      118885:data<=-16'd4020;
      118886:data<=-16'd3612;
      118887:data<=-16'd3219;
      118888:data<=-16'd2905;
      118889:data<=-16'd2893;
      118890:data<=-16'd1826;
      118891:data<=-16'd625;
      118892:data<=-16'd652;
      118893:data<=-16'd123;
      118894:data<=16'd825;
      118895:data<=16'd508;
      118896:data<=16'd1682;
      118897:data<=16'd3169;
      118898:data<=16'd2027;
      118899:data<=16'd2403;
      118900:data<=16'd2646;
      118901:data<=16'd1603;
      118902:data<=16'd4243;
      118903:data<=16'd1307;
      118904:data<=-16'd9392;
      118905:data<=-16'd11882;
      118906:data<=-16'd8771;
      118907:data<=-16'd8896;
      118908:data<=-16'd7855;
      118909:data<=-16'd6793;
      118910:data<=-16'd6178;
      118911:data<=-16'd4290;
      118912:data<=-16'd4463;
      118913:data<=-16'd4105;
      118914:data<=-16'd3160;
      118915:data<=-16'd4464;
      118916:data<=-16'd3268;
      118917:data<=-16'd607;
      118918:data<=-16'd320;
      118919:data<=-16'd332;
      118920:data<=-16'd458;
      118921:data<=-16'd155;
      118922:data<=16'd813;
      118923:data<=16'd1848;
      118924:data<=16'd3717;
      118925:data<=16'd3733;
      118926:data<=16'd3160;
      118927:data<=16'd4305;
      118928:data<=16'd3131;
      118929:data<=16'd2805;
      118930:data<=16'd5421;
      118931:data<=16'd5275;
      118932:data<=16'd6329;
      118933:data<=16'd11329;
      118934:data<=16'd13303;
      118935:data<=16'd12008;
      118936:data<=16'd12176;
      118937:data<=16'd13905;
      118938:data<=16'd13999;
      118939:data<=16'd13300;
      118940:data<=16'd14099;
      118941:data<=16'd13033;
      118942:data<=16'd12619;
      118943:data<=16'd14836;
      118944:data<=16'd13239;
      118945:data<=16'd16134;
      118946:data<=16'd27486;
      118947:data<=16'd30455;
      118948:data<=16'd27055;
      118949:data<=16'd27581;
      118950:data<=16'd26521;
      118951:data<=16'd25376;
      118952:data<=16'd25854;
      118953:data<=16'd24037;
      118954:data<=16'd23209;
      118955:data<=16'd22618;
      118956:data<=16'd21884;
      118957:data<=16'd23629;
      118958:data<=16'd22865;
      118959:data<=16'd20733;
      118960:data<=16'd20944;
      118961:data<=16'd19647;
      118962:data<=16'd18560;
      118963:data<=16'd19556;
      118964:data<=16'd19502;
      118965:data<=16'd18689;
      118966:data<=16'd17687;
      118967:data<=16'd16848;
      118968:data<=16'd16274;
      118969:data<=16'd15740;
      118970:data<=16'd17029;
      118971:data<=16'd17738;
      118972:data<=16'd15769;
      118973:data<=16'd14261;
      118974:data<=16'd13443;
      118975:data<=16'd12598;
      118976:data<=16'd12304;
      118977:data<=16'd12734;
      118978:data<=16'd13453;
      118979:data<=16'd11925;
      118980:data<=16'd10595;
      118981:data<=16'd11082;
      118982:data<=16'd8302;
      118983:data<=16'd5268;
      118984:data<=16'd4582;
      118985:data<=16'd3530;
      118986:data<=16'd4846;
      118987:data<=16'd1215;
      118988:data<=-16'd10731;
      118989:data<=-16'd14980;
      118990:data<=-16'd12575;
      118991:data<=-16'd13220;
      118992:data<=-16'd12007;
      118993:data<=-16'd11590;
      118994:data<=-16'd13819;
      118995:data<=-16'd12878;
      118996:data<=-16'd12445;
      118997:data<=-16'd13380;
      118998:data<=-16'd13132;
      118999:data<=-16'd13860;
      119000:data<=-16'd13641;
      119001:data<=-16'd12977;
      119002:data<=-16'd14041;
      119003:data<=-16'd14261;
      119004:data<=-16'd14010;
      119005:data<=-16'd13634;
      119006:data<=-16'd12756;
      119007:data<=-16'd12610;
      119008:data<=-16'd12129;
      119009:data<=-16'd12489;
      119010:data<=-16'd13966;
      119011:data<=-16'd13717;
      119012:data<=-16'd13265;
      119013:data<=-16'd13285;
      119014:data<=-16'd12433;
      119015:data<=-16'd11684;
      119016:data<=-16'd11873;
      119017:data<=-16'd13173;
      119018:data<=-16'd13109;
      119019:data<=-16'd11908;
      119020:data<=-16'd12631;
      119021:data<=-16'd12334;
      119022:data<=-16'd11709;
      119023:data<=-16'd12693;
      119024:data<=-16'd11937;
      119025:data<=-16'd12554;
      119026:data<=-16'd12859;
      119027:data<=-16'd10401;
      119028:data<=-16'd12326;
      119029:data<=-16'd8960;
      119030:data<=16'd2916;
      119031:data<=16'd4525;
      119032:data<=16'd3168;
      119033:data<=16'd8906;
      119034:data<=16'd9106;
      119035:data<=16'd7747;
      119036:data<=16'd9201;
      119037:data<=16'd6655;
      119038:data<=16'd5632;
      119039:data<=16'd6320;
      119040:data<=16'd5289;
      119041:data<=16'd5900;
      119042:data<=16'd4611;
      119043:data<=16'd2297;
      119044:data<=16'd2736;
      119045:data<=16'd2162;
      119046:data<=16'd1421;
      119047:data<=16'd1363;
      119048:data<=16'd770;
      119049:data<=16'd550;
      119050:data<=-16'd1384;
      119051:data<=-16'd2569;
      119052:data<=-16'd1146;
      119053:data<=-16'd1480;
      119054:data<=-16'd1770;
      119055:data<=-16'd1604;
      119056:data<=-16'd3539;
      119057:data<=-16'd4105;
      119058:data<=-16'd3386;
      119059:data<=-16'd3648;
      119060:data<=-16'd3871;
      119061:data<=-16'd4085;
      119062:data<=-16'd4423;
      119063:data<=-16'd5433;
      119064:data<=-16'd6053;
      119065:data<=-16'd5885;
      119066:data<=-16'd6516;
      119067:data<=-16'd5119;
      119068:data<=-16'd4331;
      119069:data<=-16'd6849;
      119070:data<=-16'd6193;
      119071:data<=-16'd9367;
      119072:data<=-16'd20460;
      119073:data<=-16'd23904;
      119074:data<=-16'd21208;
      119075:data<=-16'd21793;
      119076:data<=-16'd21411;
      119077:data<=-16'd21262;
      119078:data<=-16'd21293;
      119079:data<=-16'd19415;
      119080:data<=-16'd19396;
      119081:data<=-16'd17983;
      119082:data<=-16'd17691;
      119083:data<=-16'd23592;
      119084:data<=-16'd25693;
      119085:data<=-16'd23446;
      119086:data<=-16'd23864;
      119087:data<=-16'd22553;
      119088:data<=-16'd20254;
      119089:data<=-16'd20641;
      119090:data<=-16'd20742;
      119091:data<=-16'd20043;
      119092:data<=-16'd18882;
      119093:data<=-16'd17634;
      119094:data<=-16'd17191;
      119095:data<=-16'd16208;
      119096:data<=-16'd15292;
      119097:data<=-16'd15020;
      119098:data<=-16'd14079;
      119099:data<=-16'd12672;
      119100:data<=-16'd11318;
      119101:data<=-16'd10354;
      119102:data<=-16'd9174;
      119103:data<=-16'd7711;
      119104:data<=-16'd7080;
      119105:data<=-16'd6191;
      119106:data<=-16'd5201;
      119107:data<=-16'd4535;
      119108:data<=-16'd3576;
      119109:data<=-16'd3832;
      119110:data<=-16'd2444;
      119111:data<=-16'd80;
      119112:data<=-16'd2124;
      119113:data<=16'd1222;
      119114:data<=16'd12991;
      119115:data<=16'd17541;
      119116:data<=16'd16193;
      119117:data<=16'd17109;
      119118:data<=16'd16252;
      119119:data<=16'd15556;
      119120:data<=16'd16119;
      119121:data<=16'd14784;
      119122:data<=16'd14969;
      119123:data<=16'd16342;
      119124:data<=16'd16639;
      119125:data<=16'd16735;
      119126:data<=16'd15905;
      119127:data<=16'd15811;
      119128:data<=16'd15926;
      119129:data<=16'd15200;
      119130:data<=16'd16503;
      119131:data<=16'd16261;
      119132:data<=16'd14694;
      119133:data<=16'd18148;
      119134:data<=16'd21088;
      119135:data<=16'd20249;
      119136:data<=16'd21076;
      119137:data<=16'd21540;
      119138:data<=16'd20286;
      119139:data<=16'd20027;
      119140:data<=16'd19388;
      119141:data<=16'd18081;
      119142:data<=16'd17682;
      119143:data<=16'd18395;
      119144:data<=16'd18798;
      119145:data<=16'd17503;
      119146:data<=16'd16336;
      119147:data<=16'd16045;
      119148:data<=16'd15722;
      119149:data<=16'd15952;
      119150:data<=16'd16295;
      119151:data<=16'd16409;
      119152:data<=16'd15255;
      119153:data<=16'd13849;
      119154:data<=16'd15361;
      119155:data<=16'd12366;
      119156:data<=16'd2218;
      119157:data<=-16'd1689;
      119158:data<=16'd206;
      119159:data<=-16'd529;
      119160:data<=-16'd97;
      119161:data<=16'd337;
      119162:data<=-16'd550;
      119163:data<=16'd1624;
      119164:data<=16'd2291;
      119165:data<=16'd607;
      119166:data<=16'd1284;
      119167:data<=16'd1339;
      119168:data<=16'd596;
      119169:data<=16'd1315;
      119170:data<=16'd1753;
      119171:data<=16'd2106;
      119172:data<=16'd2443;
      119173:data<=16'd2522;
      119174:data<=16'd2613;
      119175:data<=16'd2426;
      119176:data<=16'd3635;
      119177:data<=16'd4561;
      119178:data<=16'd3454;
      119179:data<=16'd3315;
      119180:data<=16'd2666;
      119181:data<=16'd1683;
      119182:data<=16'd3551;
      119183:data<=16'd2554;
      119184:data<=-16'd2221;
      119185:data<=-16'd3371;
      119186:data<=-16'd2581;
      119187:data<=-16'd3160;
      119188:data<=-16'd2353;
      119189:data<=-16'd643;
      119190:data<=-16'd288;
      119191:data<=-16'd182;
      119192:data<=16'd111;
      119193:data<=-16'd892;
      119194:data<=-16'd1221;
      119195:data<=16'd240;
      119196:data<=16'd376;
      119197:data<=16'd3727;
      119198:data<=16'd13203;
      119199:data<=16'd17337;
      119200:data<=16'd14471;
      119201:data<=16'd14149;
      119202:data<=16'd14258;
      119203:data<=16'd12530;
      119204:data<=16'd12413;
      119205:data<=16'd11838;
      119206:data<=16'd10252;
      119207:data<=16'd9644;
      119208:data<=16'd8578;
      119209:data<=16'd6752;
      119210:data<=16'd5906;
      119211:data<=16'd6507;
      119212:data<=16'd6411;
      119213:data<=16'd4795;
      119214:data<=16'd4062;
      119215:data<=16'd3177;
      119216:data<=16'd1016;
      119217:data<=16'd596;
      119218:data<=16'd1254;
      119219:data<=16'd761;
      119220:data<=16'd241;
      119221:data<=16'd252;
      119222:data<=-16'd196;
      119223:data<=-16'd1986;
      119224:data<=-16'd3374;
      119225:data<=-16'd2972;
      119226:data<=-16'd2987;
      119227:data<=-16'd2969;
      119228:data<=-16'd2855;
      119229:data<=-16'd4748;
      119230:data<=-16'd5465;
      119231:data<=-16'd4965;
      119232:data<=-16'd6223;
      119233:data<=-16'd4710;
      119234:data<=-16'd109;
      119235:data<=16'd1061;
      119236:data<=-16'd1569;
      119237:data<=-16'd3112;
      119238:data<=-16'd1560;
      119239:data<=-16'd3962;
      119240:data<=-16'd13512;
      119241:data<=-16'd18971;
      119242:data<=-16'd18211;
      119243:data<=-16'd18983;
      119244:data<=-16'd18601;
      119245:data<=-16'd16854;
      119246:data<=-16'd17437;
      119247:data<=-16'd16647;
      119248:data<=-16'd15778;
      119249:data<=-16'd17576;
      119250:data<=-16'd17738;
      119251:data<=-16'd16531;
      119252:data<=-16'd16568;
      119253:data<=-16'd16522;
      119254:data<=-16'd16190;
      119255:data<=-16'd16381;
      119256:data<=-16'd17015;
      119257:data<=-16'd16775;
      119258:data<=-16'd15464;
      119259:data<=-16'd15153;
      119260:data<=-16'd15130;
      119261:data<=-16'd14643;
      119262:data<=-16'd15244;
      119263:data<=-16'd15708;
      119264:data<=-16'd15382;
      119265:data<=-16'd15039;
      119266:data<=-16'd13599;
      119267:data<=-16'd12248;
      119268:data<=-16'd12812;
      119269:data<=-16'd13806;
      119270:data<=-16'd13543;
      119271:data<=-16'd12637;
      119272:data<=-16'd12657;
      119273:data<=-16'd12328;
      119274:data<=-16'd10988;
      119275:data<=-16'd11521;
      119276:data<=-16'd12862;
      119277:data<=-16'd12649;
      119278:data<=-16'd11588;
      119279:data<=-16'd10293;
      119280:data<=-16'd11107;
      119281:data<=-16'd9523;
      119282:data<=16'd36;
      119283:data<=16'd4431;
      119284:data<=-16'd1717;
      119285:data<=-16'd3918;
      119286:data<=-16'd2419;
      119287:data<=-16'd3216;
      119288:data<=-16'd2413;
      119289:data<=-16'd2936;
      119290:data<=-16'd4807;
      119291:data<=-16'd3213;
      119292:data<=-16'd2485;
      119293:data<=-16'd3206;
      119294:data<=-16'd2605;
      119295:data<=-16'd3401;
      119296:data<=-16'd4470;
      119297:data<=-16'd3977;
      119298:data<=-16'd3562;
      119299:data<=-16'd3325;
      119300:data<=-16'd3425;
      119301:data<=-16'd3836;
      119302:data<=-16'd4410;
      119303:data<=-16'd5039;
      119304:data<=-16'd4422;
      119305:data<=-16'd3453;
      119306:data<=-16'd3071;
      119307:data<=-16'd2790;
      119308:data<=-16'd3219;
      119309:data<=-16'd3268;
      119310:data<=-16'd2484;
      119311:data<=-16'd2181;
      119312:data<=-16'd1820;
      119313:data<=-16'd1612;
      119314:data<=-16'd1439;
      119315:data<=-16'd281;
      119316:data<=16'd740;
      119317:data<=16'd1272;
      119318:data<=16'd1676;
      119319:data<=16'd2005;
      119320:data<=16'd2141;
      119321:data<=16'd2417;
      119322:data<=16'd5051;
      119323:data<=16'd4585;
      119324:data<=-16'd4557;
      119325:data<=-16'd11103;
      119326:data<=-16'd9824;
      119327:data<=-16'd9047;
      119328:data<=-16'd7840;
      119329:data<=-16'd5457;
      119330:data<=-16'd5259;
      119331:data<=-16'd4739;
      119332:data<=-16'd4404;
      119333:data<=-16'd3153;
      119334:data<=16'd1736;
      119335:data<=16'd5054;
      119336:data<=16'd5949;
      119337:data<=16'd6537;
      119338:data<=16'd5427;
      119339:data<=16'd5256;
      119340:data<=16'd5982;
      119341:data<=16'd6120;
      119342:data<=16'd8040;
      119343:data<=16'd9317;
      119344:data<=16'd8604;
      119345:data<=16'd8548;
      119346:data<=16'd8422;
      119347:data<=16'd7991;
      119348:data<=16'd7856;
      119349:data<=16'd8680;
      119350:data<=16'd10422;
      119351:data<=16'd10114;
      119352:data<=16'd9097;
      119353:data<=16'd9367;
      119354:data<=16'd9130;
      119355:data<=16'd9925;
      119356:data<=16'd11083;
      119357:data<=16'd10624;
      119358:data<=16'd10956;
      119359:data<=16'd10944;
      119360:data<=16'd9941;
      119361:data<=16'd10419;
      119362:data<=16'd11841;
      119363:data<=16'd13256;
      119364:data<=16'd12527;
      119365:data<=16'd12736;
      119366:data<=16'd20168;
      119367:data<=16'd26597;
      119368:data<=16'd26200;
      119369:data<=16'd26488;
      119370:data<=16'd26520;
      119371:data<=16'd24256;
      119372:data<=16'd23848;
      119373:data<=16'd23253;
      119374:data<=16'd21930;
      119375:data<=16'd22189;
      119376:data<=16'd22014;
      119377:data<=16'd20742;
      119378:data<=16'd19761;
      119379:data<=16'd19887;
      119380:data<=16'd19748;
      119381:data<=16'd18807;
      119382:data<=16'd19849;
      119383:data<=16'd18862;
      119384:data<=16'd12948;
      119385:data<=16'd10328;
      119386:data<=16'd11304;
      119387:data<=16'd10146;
      119388:data<=16'd9870;
      119389:data<=16'd11232;
      119390:data<=16'd11203;
      119391:data<=16'd10269;
      119392:data<=16'd9054;
      119393:data<=16'd8244;
      119394:data<=16'd8332;
      119395:data<=16'd8916;
      119396:data<=16'd9253;
      119397:data<=16'd8733;
      119398:data<=16'd8907;
      119399:data<=16'd8818;
      119400:data<=16'd7065;
      119401:data<=16'd7333;
      119402:data<=16'd8904;
      119403:data<=16'd8499;
      119404:data<=16'd7551;
      119405:data<=16'd6404;
      119406:data<=16'd6642;
      119407:data<=16'd6778;
      119408:data<=-16'd64;
      119409:data<=-16'd8017;
      119410:data<=-16'd8537;
      119411:data<=-16'd7421;
      119412:data<=-16'd7574;
      119413:data<=-16'd6983;
      119414:data<=-16'd7635;
      119415:data<=-16'd8153;
      119416:data<=-16'd7342;
      119417:data<=-16'd7216;
      119418:data<=-16'd7004;
      119419:data<=-16'd6536;
      119420:data<=-16'd6696;
      119421:data<=-16'd7192;
      119422:data<=-16'd8228;
      119423:data<=-16'd8718;
      119424:data<=-16'd8038;
      119425:data<=-16'd7832;
      119426:data<=-16'd7758;
      119427:data<=-16'd6924;
      119428:data<=-16'd7511;
      119429:data<=-16'd9859;
      119430:data<=-16'd10140;
      119431:data<=-16'd8780;
      119432:data<=-16'd9294;
      119433:data<=-16'd8252;
      119434:data<=-16'd4264;
      119435:data<=-16'd3128;
      119436:data<=-16'd3926;
      119437:data<=-16'd3354;
      119438:data<=-16'd3372;
      119439:data<=-16'd3421;
      119440:data<=-16'd3378;
      119441:data<=-16'd4316;
      119442:data<=-16'd4675;
      119443:data<=-16'd5178;
      119444:data<=-16'd5271;
      119445:data<=-16'd4353;
      119446:data<=-16'd4578;
      119447:data<=-16'd3876;
      119448:data<=-16'd4790;
      119449:data<=-16'd8161;
      119450:data<=-16'd1911;
      119451:data<=16'd8994;
      119452:data<=16'd9500;
      119453:data<=16'd7595;
      119454:data<=16'd8269;
      119455:data<=16'd5586;
      119456:data<=16'd4316;
      119457:data<=16'd5090;
      119458:data<=16'd4106;
      119459:data<=16'd4128;
      119460:data<=16'd4179;
      119461:data<=16'd3018;
      119462:data<=16'd1768;
      119463:data<=16'd353;
      119464:data<=16'd725;
      119465:data<=16'd1286;
      119466:data<=16'd461;
      119467:data<=16'd490;
      119468:data<=-16'd945;
      119469:data<=-16'd3483;
      119470:data<=-16'd3415;
      119471:data<=-16'd3034;
      119472:data<=-16'd3369;
      119473:data<=-16'd3189;
      119474:data<=-16'd3603;
      119475:data<=-16'd4645;
      119476:data<=-16'd5163;
      119477:data<=-16'd4795;
      119478:data<=-16'd5212;
      119479:data<=-16'd5733;
      119480:data<=-16'd4485;
      119481:data<=-16'd5285;
      119482:data<=-16'd7050;
      119483:data<=-16'd6748;
      119484:data<=-16'd9908;
      119485:data<=-16'd13852;
      119486:data<=-16'd13230;
      119487:data<=-16'd13041;
      119488:data<=-16'd13729;
      119489:data<=-16'd14298;
      119490:data<=-16'd14149;
      119491:data<=-16'd11884;
      119492:data<=-16'd16950;
      119493:data<=-16'd27102;
      119494:data<=-16'd28368;
      119495:data<=-16'd27076;
      119496:data<=-16'd28127;
      119497:data<=-16'd25919;
      119498:data<=-16'd24905;
      119499:data<=-16'd24748;
      119500:data<=-16'd22583;
      119501:data<=-16'd22776;
      119502:data<=-16'd22967;
      119503:data<=-16'd21601;
      119504:data<=-16'd21171;
      119505:data<=-16'd20052;
      119506:data<=-16'd19143;
      119507:data<=-16'd19397;
      119508:data<=-16'd19637;
      119509:data<=-16'd19637;
      119510:data<=-16'd18363;
      119511:data<=-16'd17286;
      119512:data<=-16'd16774;
      119513:data<=-16'd15614;
      119514:data<=-16'd15960;
      119515:data<=-16'd16389;
      119516:data<=-16'd15352;
      119517:data<=-16'd14913;
      119518:data<=-16'd14189;
      119519:data<=-16'd13367;
      119520:data<=-16'd12584;
      119521:data<=-16'd10827;
      119522:data<=-16'd9746;
      119523:data<=-16'd8660;
      119524:data<=-16'd8222;
      119525:data<=-16'd8827;
      119526:data<=-16'd6872;
      119527:data<=-16'd4717;
      119528:data<=-16'd2886;
      119529:data<=-16'd334;
      119530:data<=-16'd1284;
      119531:data<=-16'd540;
      119532:data<=16'd1133;
      119533:data<=-16'd2358;
      119534:data<=16'd4796;
      119535:data<=16'd21376;
      119536:data<=16'd24438;
      119537:data<=16'd21188;
      119538:data<=16'd22465;
      119539:data<=16'd21033;
      119540:data<=16'd19902;
      119541:data<=16'd21349;
      119542:data<=16'd21317;
      119543:data<=16'd21090;
      119544:data<=16'd20439;
      119545:data<=16'd19590;
      119546:data<=16'd19403;
      119547:data<=16'd19326;
      119548:data<=16'd20360;
      119549:data<=16'd20290;
      119550:data<=16'd18998;
      119551:data<=16'd19147;
      119552:data<=16'd18522;
      119553:data<=16'd17340;
      119554:data<=16'd17529;
      119555:data<=16'd18216;
      119556:data<=16'd18923;
      119557:data<=16'd18148;
      119558:data<=16'd17136;
      119559:data<=16'd16982;
      119560:data<=16'd15703;
      119561:data<=16'd16161;
      119562:data<=16'd17585;
      119563:data<=16'd16245;
      119564:data<=16'd15656;
      119565:data<=16'd15391;
      119566:data<=16'd14025;
      119567:data<=16'd14527;
      119568:data<=16'd15086;
      119569:data<=16'd15145;
      119570:data<=16'd14694;
      119571:data<=16'd13082;
      119572:data<=16'd13126;
      119573:data<=16'd11523;
      119574:data<=16'd10596;
      119575:data<=16'd15133;
      119576:data<=16'd10803;
      119577:data<=-16'd1798;
      119578:data<=-16'd4128;
      119579:data<=-16'd2018;
      119580:data<=-16'd2913;
      119581:data<=-16'd1403;
      119582:data<=-16'd728;
      119583:data<=-16'd913;
      119584:data<=-16'd789;
      119585:data<=-16'd3953;
      119586:data<=-16'd5351;
      119587:data<=-16'd3651;
      119588:data<=-16'd3283;
      119589:data<=-16'd2764;
      119590:data<=-16'd2649;
      119591:data<=-16'd2887;
      119592:data<=-16'd2009;
      119593:data<=-16'd2566;
      119594:data<=-16'd2573;
      119595:data<=-16'd309;
      119596:data<=16'd303;
      119597:data<=-16'd464;
      119598:data<=-16'd185;
      119599:data<=16'd428;
      119600:data<=16'd426;
      119601:data<=16'd649;
      119602:data<=16'd1507;
      119603:data<=16'd1278;
      119604:data<=16'd930;
      119605:data<=16'd1410;
      119606:data<=16'd884;
      119607:data<=16'd1357;
      119608:data<=16'd2761;
      119609:data<=16'd2645;
      119610:data<=16'd3121;
      119611:data<=16'd3095;
      119612:data<=16'd2596;
      119613:data<=16'd3891;
      119614:data<=16'd3559;
      119615:data<=16'd4026;
      119616:data<=16'd5477;
      119617:data<=16'd2839;
      119618:data<=16'd6912;
      119619:data<=16'd18337;
      119620:data<=16'd20401;
      119621:data<=16'd17960;
      119622:data<=16'd19218;
      119623:data<=16'd18328;
      119624:data<=16'd17346;
      119625:data<=16'd17428;
      119626:data<=16'd15722;
      119627:data<=16'd14766;
      119628:data<=16'd14099;
      119629:data<=16'd13167;
      119630:data<=16'd12665;
      119631:data<=16'd11838;
      119632:data<=16'd11885;
      119633:data<=16'd10928;
      119634:data<=16'd9344;
      119635:data<=16'd10551;
      119636:data<=16'd10816;
      119637:data<=16'd9444;
      119638:data<=16'd9547;
      119639:data<=16'd9056;
      119640:data<=16'd7723;
      119641:data<=16'd6175;
      119642:data<=16'd4564;
      119643:data<=16'd4373;
      119644:data<=16'd4056;
      119645:data<=16'd3629;
      119646:data<=16'd3741;
      119647:data<=16'd2576;
      119648:data<=16'd776;
      119649:data<=-16'd1010;
      119650:data<=-16'd1345;
      119651:data<=-16'd428;
      119652:data<=-16'd1632;
      119653:data<=-16'd2043;
      119654:data<=-16'd2394;
      119655:data<=-16'd5747;
      119656:data<=-16'd5510;
      119657:data<=-16'd4584;
      119658:data<=-16'd6384;
      119659:data<=-16'd4240;
      119660:data<=-16'd8037;
      119661:data<=-16'd20407;
      119662:data<=-16'd23658;
      119663:data<=-16'd21268;
      119664:data<=-16'd22419;
      119665:data<=-16'd21211;
      119666:data<=-16'd19620;
      119667:data<=-16'd20845;
      119668:data<=-16'd21651;
      119669:data<=-16'd21634;
      119670:data<=-16'd20821;
      119671:data<=-16'd20139;
      119672:data<=-16'd19470;
      119673:data<=-16'd18534;
      119674:data<=-16'd19685;
      119675:data<=-16'd20528;
      119676:data<=-16'd19405;
      119677:data<=-16'd18997;
      119678:data<=-16'd18741;
      119679:data<=-16'd17951;
      119680:data<=-16'd17054;
      119681:data<=-16'd17189;
      119682:data<=-16'd18236;
      119683:data<=-16'd17156;
      119684:data<=-16'd17696;
      119685:data<=-16'd21053;
      119686:data<=-16'd20475;
      119687:data<=-16'd19725;
      119688:data<=-16'd21693;
      119689:data<=-16'd20800;
      119690:data<=-16'd19328;
      119691:data<=-16'd18750;
      119692:data<=-16'd17561;
      119693:data<=-16'd17620;
      119694:data<=-16'd17479;
      119695:data<=-16'd17512;
      119696:data<=-16'd17411;
      119697:data<=-16'd15476;
      119698:data<=-16'd15358;
      119699:data<=-16'd14202;
      119700:data<=-16'd12536;
      119701:data<=-16'd15940;
      119702:data<=-16'd12105;
      119703:data<=16'd36;
      119704:data<=16'd2808;
      119705:data<=16'd1074;
      119706:data<=16'd3099;
      119707:data<=16'd2033;
      119708:data<=-16'd68;
      119709:data<=16'd394;
      119710:data<=16'd764;
      119711:data<=16'd867;
      119712:data<=16'd447;
      119713:data<=16'd82;
      119714:data<=-16'd197;
      119715:data<=-16'd1181;
      119716:data<=-16'd939;
      119717:data<=-16'd305;
      119718:data<=-16'd453;
      119719:data<=16'd153;
      119720:data<=16'd323;
      119721:data<=-16'd957;
      119722:data<=-16'd2168;
      119723:data<=-16'd2173;
      119724:data<=-16'd1897;
      119725:data<=-16'd2226;
      119726:data<=-16'd1528;
      119727:data<=-16'd1209;
      119728:data<=-16'd2229;
      119729:data<=-16'd1521;
      119730:data<=-16'd1636;
      119731:data<=-16'd2946;
      119732:data<=-16'd1851;
      119733:data<=-16'd1842;
      119734:data<=-16'd1086;
      119735:data<=16'd2966;
      119736:data<=16'd3635;
      119737:data<=16'd3015;
      119738:data<=16'd3674;
      119739:data<=16'd2165;
      119740:data<=16'd2966;
      119741:data<=16'd4755;
      119742:data<=16'd4275;
      119743:data<=16'd5879;
      119744:data<=16'd2302;
      119745:data<=-16'd8263;
      119746:data<=-16'd11617;
      119747:data<=-16'd8470;
      119748:data<=-16'd7304;
      119749:data<=-16'd7025;
      119750:data<=-16'd6728;
      119751:data<=-16'd6329;
      119752:data<=-16'd5914;
      119753:data<=-16'd5233;
      119754:data<=-16'd3213;
      119755:data<=-16'd2748;
      119756:data<=-16'd3157;
      119757:data<=-16'd1683;
      119758:data<=-16'd1717;
      119759:data<=-16'd2689;
      119760:data<=-16'd1551;
      119761:data<=-16'd241;
      119762:data<=16'd831;
      119763:data<=16'd1683;
      119764:data<=16'd1668;
      119765:data<=16'd1862;
      119766:data<=16'd2006;
      119767:data<=16'd2623;
      119768:data<=16'd4023;
      119769:data<=16'd4138;
      119770:data<=16'd3504;
      119771:data<=16'd3500;
      119772:data<=16'd3689;
      119773:data<=16'd3933;
      119774:data<=16'd4604;
      119775:data<=16'd5899;
      119776:data<=16'd6410;
      119777:data<=16'd6296;
      119778:data<=16'd6534;
      119779:data<=16'd5401;
      119780:data<=16'd6006;
      119781:data<=16'd9247;
      119782:data<=16'd8737;
      119783:data<=16'd8105;
      119784:data<=16'd8692;
      119785:data<=16'd3994;
      119786:data<=16'd5398;
      119787:data<=16'd17488;
      119788:data<=16'd22277;
      119789:data<=16'd19657;
      119790:data<=16'd20016;
      119791:data<=16'd19858;
      119792:data<=16'd18597;
      119793:data<=16'd18729;
      119794:data<=16'd19064;
      119795:data<=16'd19331;
      119796:data<=16'd18469;
      119797:data<=16'd17840;
      119798:data<=16'd17805;
      119799:data<=16'd16365;
      119800:data<=16'd16956;
      119801:data<=16'd19035;
      119802:data<=16'd18299;
      119803:data<=16'd17223;
      119804:data<=16'd16501;
      119805:data<=16'd15359;
      119806:data<=16'd15538;
      119807:data<=16'd15505;
      119808:data<=16'd14968;
      119809:data<=16'd14942;
      119810:data<=16'd14539;
      119811:data<=16'd14327;
      119812:data<=16'd13832;
      119813:data<=16'd13391;
      119814:data<=16'd14422;
      119815:data<=16'd14519;
      119816:data<=16'd13394;
      119817:data<=16'd12833;
      119818:data<=16'd12043;
      119819:data<=16'd11389;
      119820:data<=16'd11515;
      119821:data<=16'd12005;
      119822:data<=16'd11743;
      119823:data<=16'd10466;
      119824:data<=16'd10443;
      119825:data<=16'd9984;
      119826:data<=16'd8810;
      119827:data<=16'd10537;
      119828:data<=16'd8070;
      119829:data<=-16'd1413;
      119830:data<=-16'd5897;
      119831:data<=-16'd4742;
      119832:data<=-16'd5060;
      119833:data<=-16'd5109;
      119834:data<=-16'd3524;
      119835:data<=-16'd996;
      119836:data<=16'd970;
      119837:data<=16'd729;
      119838:data<=16'd678;
      119839:data<=16'd828;
      119840:data<=16'd133;
      119841:data<=-16'd259;
      119842:data<=-16'd1251;
      119843:data<=-16'd1488;
      119844:data<=-16'd500;
      119845:data<=-16'd949;
      119846:data<=-16'd1638;
      119847:data<=-16'd2663;
      119848:data<=-16'd3912;
      119849:data<=-16'd2820;
      119850:data<=-16'd2517;
      119851:data<=-16'd3535;
      119852:data<=-16'd3099;
      119853:data<=-16'd3815;
      119854:data<=-16'd5128;
      119855:data<=-16'd5304;
      119856:data<=-16'd5912;
      119857:data<=-16'd5762;
      119858:data<=-16'd5139;
      119859:data<=-16'd5212;
      119860:data<=-16'd5594;
      119861:data<=-16'd6863;
      119862:data<=-16'd7134;
      119863:data<=-16'd6516;
      119864:data<=-16'd6567;
      119865:data<=-16'd5843;
      119866:data<=-16'd6522;
      119867:data<=-16'd7759;
      119868:data<=-16'd7225;
      119869:data<=-16'd8795;
      119870:data<=-16'd6293;
      119871:data<=16'd4303;
      119872:data<=16'd9556;
      119873:data<=16'd7298;
      119874:data<=16'd5782;
      119875:data<=16'd4707;
      119876:data<=16'd4419;
      119877:data<=16'd4875;
      119878:data<=16'd4560;
      119879:data<=16'd4541;
      119880:data<=16'd3121;
      119881:data<=16'd1119;
      119882:data<=16'd779;
      119883:data<=16'd517;
      119884:data<=16'd608;
      119885:data<=-16'd588;
      119886:data<=-16'd3836;
      119887:data<=-16'd5096;
      119888:data<=-16'd5513;
      119889:data<=-16'd6302;
      119890:data<=-16'd5753;
      119891:data<=-16'd5582;
      119892:data<=-16'd5535;
      119893:data<=-16'd5950;
      119894:data<=-16'd8046;
      119895:data<=-16'd8313;
      119896:data<=-16'd7124;
      119897:data<=-16'd6904;
      119898:data<=-16'd6449;
      119899:data<=-16'd6616;
      119900:data<=-16'd7612;
      119901:data<=-16'd8009;
      119902:data<=-16'd7667;
      119903:data<=-16'd7089;
      119904:data<=-16'd7550;
      119905:data<=-16'd7503;
      119906:data<=-16'd7210;
      119907:data<=-16'd9213;
      119908:data<=-16'd9559;
      119909:data<=-16'd8575;
      119910:data<=-16'd9360;
      119911:data<=-16'd7635;
      119912:data<=-16'd8978;
      119913:data<=-16'd18944;
      119914:data<=-16'd25205;
      119915:data<=-16'd23605;
      119916:data<=-16'd22231;
      119917:data<=-16'd21936;
      119918:data<=-16'd21121;
      119919:data<=-16'd20384;
      119920:data<=-16'd20456;
      119921:data<=-16'd20794;
      119922:data<=-16'd19892;
      119923:data<=-16'd19276;
      119924:data<=-16'd18804;
      119925:data<=-16'd17473;
      119926:data<=-16'd17587;
      119927:data<=-16'd18043;
      119928:data<=-16'd17717;
      119929:data<=-16'd17500;
      119930:data<=-16'd15995;
      119931:data<=-16'd14853;
      119932:data<=-16'd14653;
      119933:data<=-16'd13931;
      119934:data<=-16'd14528;
      119935:data<=-16'd13397;
      119936:data<=-16'd9450;
      119937:data<=-16'd8470;
      119938:data<=-16'd8680;
      119939:data<=-16'd7824;
      119940:data<=-16'd8420;
      119941:data<=-16'd8725;
      119942:data<=-16'd8501;
      119943:data<=-16'd8419;
      119944:data<=-16'd7228;
      119945:data<=-16'd6554;
      119946:data<=-16'd6213;
      119947:data<=-16'd5344;
      119948:data<=-16'd4751;
      119949:data<=-16'd3959;
      119950:data<=-16'd3976;
      119951:data<=-16'd3751;
      119952:data<=-16'd2775;
      119953:data<=-16'd3456;
      119954:data<=16'd284;
      119955:data<=16'd10299;
      119956:data<=16'd15570;
      119957:data<=16'd14803;
      119958:data<=16'd14196;
      119959:data<=16'd14478;
      119960:data<=16'd15829;
      119961:data<=16'd16330;
      119962:data<=16'd15085;
      119963:data<=16'd14982;
      119964:data<=16'd15029;
      119965:data<=16'd14328;
      119966:data<=16'd14590;
      119967:data<=16'd15464;
      119968:data<=16'd15960;
      119969:data<=16'd15271;
      119970:data<=16'd14572;
      119971:data<=16'd14698;
      119972:data<=16'd13681;
      119973:data<=16'd13549;
      119974:data<=16'd15362;
      119975:data<=16'd15006;
      119976:data<=16'd13702;
      119977:data<=16'd13788;
      119978:data<=16'd13098;
      119979:data<=16'd12501;
      119980:data<=16'd13433;
      119981:data<=16'd14099;
      119982:data<=16'd13691;
      119983:data<=16'd13383;
      119984:data<=16'd13136;
      119985:data<=16'd10654;
      119986:data<=16'd7953;
      119987:data<=16'd8725;
      119988:data<=16'd9141;
      119989:data<=16'd7611;
      119990:data<=16'd7486;
      119991:data<=16'd7168;
      119992:data<=16'd6833;
      119993:data<=16'd7918;
      119994:data<=16'd7905;
      119995:data<=16'd8316;
      119996:data<=16'd7148;
      119997:data<=-16'd1127;
      119998:data<=-16'd8302;
      119999:data<=-16'd7148;
      120000:data<=-16'd4807;
      120001:data<=-16'd4805;
      120002:data<=-16'd4678;
      120003:data<=-16'd4476;
      120004:data<=-16'd4305;
      120005:data<=-16'd4262;
      120006:data<=-16'd3818;
      120007:data<=-16'd2237;
      120008:data<=-16'd1498;
      120009:data<=-16'd2170;
      120010:data<=-16'd2441;
      120011:data<=-16'd2202;
      120012:data<=-16'd1861;
      120013:data<=-16'd898;
      120014:data<=16'd405;
      120015:data<=16'd725;
      120016:data<=16'd472;
      120017:data<=16'd820;
      120018:data<=16'd607;
      120019:data<=16'd391;
      120020:data<=16'd1780;
      120021:data<=16'd2414;
      120022:data<=16'd1870;
      120023:data<=16'd2032;
      120024:data<=16'd1548;
      120025:data<=16'd846;
      120026:data<=16'd1974;
      120027:data<=16'd3416;
      120028:data<=16'd3422;
      120029:data<=16'd2766;
      120030:data<=16'd2775;
      120031:data<=16'd2963;
      120032:data<=16'd3248;
      120033:data<=16'd4476;
      120034:data<=16'd4646;
      120035:data<=16'd5372;
      120036:data<=16'd9054;
      120037:data<=16'd9345;
      120038:data<=16'd8762;
      120039:data<=16'd16695;
      120040:data<=16'd24700;
      120041:data<=16'd24614;
      120042:data<=16'd22768;
      120043:data<=16'd21784;
      120044:data<=16'd21214;
      120045:data<=16'd20989;
      120046:data<=16'd19858;
      120047:data<=16'd19939;
      120048:data<=16'd20110;
      120049:data<=16'd18324;
      120050:data<=16'd17455;
      120051:data<=16'd16976;
      120052:data<=16'd15998;
      120053:data<=16'd15564;
      120054:data<=16'd14537;
      120055:data<=16'd13947;
      120056:data<=16'd13373;
      120057:data<=16'd11618;
      120058:data<=16'd11445;
      120059:data<=16'd11191;
      120060:data<=16'd8980;
      120061:data<=16'd7952;
      120062:data<=16'd7436;
      120063:data<=16'd6307;
      120064:data<=16'd6003;
      120065:data<=16'd5990;
      120066:data<=16'd5377;
      120067:data<=16'd3709;
      120068:data<=16'd2228;
      120069:data<=16'd1920;
      120070:data<=16'd1374;
      120071:data<=16'd1365;
      120072:data<=16'd1152;
      120073:data<=-16'd854;
      120074:data<=-16'd1709;
      120075:data<=-16'd2003;
      120076:data<=-16'd3134;
      120077:data<=-16'd2855;
      120078:data<=-16'd3040;
      120079:data<=-16'd3829;
      120080:data<=-16'd5072;
      120081:data<=-16'd12123;
      120082:data<=-16'd20604;
      120083:data<=-16'd21485;
      120084:data<=-16'd18630;
      120085:data<=-16'd18929;
      120086:data<=-16'd22410;
      120087:data<=-16'd25000;
      120088:data<=-16'd24278;
      120089:data<=-16'd23178;
      120090:data<=-16'd22773;
      120091:data<=-16'd21579;
      120092:data<=-16'd21244;
      120093:data<=-16'd22025;
      120094:data<=-16'd22121;
      120095:data<=-16'd21271;
      120096:data<=-16'd20274;
      120097:data<=-16'd20057;
      120098:data<=-16'd19499;
      120099:data<=-16'd18531;
      120100:data<=-16'd19193;
      120101:data<=-16'd19481;
      120102:data<=-16'd18016;
      120103:data<=-16'd17370;
      120104:data<=-16'd17171;
      120105:data<=-16'd16648;
      120106:data<=-16'd17127;
      120107:data<=-16'd17670;
      120108:data<=-16'd17208;
      120109:data<=-16'd16775;
      120110:data<=-16'd16665;
      120111:data<=-16'd15632;
      120112:data<=-16'd14457;
      120113:data<=-16'd15446;
      120114:data<=-16'd16205;
      120115:data<=-16'd14871;
      120116:data<=-16'd14566;
      120117:data<=-16'd13976;
      120118:data<=-16'd12128;
      120119:data<=-16'd12718;
      120120:data<=-16'd12994;
      120121:data<=-16'd12055;
      120122:data<=-16'd12639;
      120123:data<=-16'd7259;
      120124:data<=16'd3200;
      120125:data<=16'd5303;
      120126:data<=16'd1882;
      120127:data<=16'd1785;
      120128:data<=16'd2173;
      120129:data<=16'd2188;
      120130:data<=16'd2682;
      120131:data<=16'd2070;
      120132:data<=16'd1853;
      120133:data<=16'd1384;
      120134:data<=-16'd200;
      120135:data<=16'd738;
      120136:data<=16'd3836;
      120137:data<=16'd5348;
      120138:data<=16'd5171;
      120139:data<=16'd4384;
      120140:data<=16'd3107;
      120141:data<=16'd2332;
      120142:data<=16'd2928;
      120143:data<=16'd3450;
      120144:data<=16'd2854;
      120145:data<=16'd2161;
      120146:data<=16'd1306;
      120147:data<=16'd509;
      120148:data<=16'd822;
      120149:data<=16'd1304;
      120150:data<=16'd1457;
      120151:data<=16'd1434;
      120152:data<=16'd644;
      120153:data<=-16'd540;
      120154:data<=-16'd1287;
      120155:data<=-16'd704;
      120156:data<=16'd20;
      120157:data<=-16'd767;
      120158:data<=-16'd764;
      120159:data<=-16'd428;
      120160:data<=-16'd963;
      120161:data<=16'd290;
      120162:data<=16'd147;
      120163:data<=-16'd1256;
      120164:data<=16'd405;
      120165:data<=-16'd3698;
      120166:data<=-16'd13118;
      120167:data<=-16'd13926;
      120168:data<=-16'd11095;
      120169:data<=-16'd11670;
      120170:data<=-16'd10657;
      120171:data<=-16'd10199;
      120172:data<=-16'd10292;
      120173:data<=-16'd7733;
      120174:data<=-16'd6774;
      120175:data<=-16'd6739;
      120176:data<=-16'd5479;
      120177:data<=-16'd5761;
      120178:data<=-16'd5973;
      120179:data<=-16'd4519;
      120180:data<=-16'd2986;
      120181:data<=-16'd1961;
      120182:data<=-16'd1950;
      120183:data<=-16'd2020;
      120184:data<=-16'd1475;
      120185:data<=-16'd1513;
      120186:data<=-16'd2428;
      120187:data<=-16'd3433;
      120188:data<=-16'd3268;
      120189:data<=-16'd2582;
      120190:data<=-16'd2880;
      120191:data<=-16'd3134;
      120192:data<=-16'd2473;
      120193:data<=-16'd879;
      120194:data<=16'd443;
      120195:data<=16'd450;
      120196:data<=16'd1057;
      120197:data<=16'd1289;
      120198:data<=16'd782;
      120199:data<=16'd2529;
      120200:data<=16'd3689;
      120201:data<=16'd3688;
      120202:data<=16'd4667;
      120203:data<=16'd3650;
      120204:data<=16'd4055;
      120205:data<=16'd5934;
      120206:data<=16'd4237;
      120207:data<=16'd9012;
      120208:data<=16'd19843;
      120209:data<=16'd21416;
      120210:data<=16'd18638;
      120211:data<=16'd18864;
      120212:data<=16'd18636;
      120213:data<=16'd19973;
      120214:data<=16'd20609;
      120215:data<=16'd18395;
      120216:data<=16'd18161;
      120217:data<=16'd17864;
      120218:data<=16'd16741;
      120219:data<=16'd18011;
      120220:data<=16'd18595;
      120221:data<=16'd17453;
      120222:data<=16'd17020;
      120223:data<=16'd16792;
      120224:data<=16'd15823;
      120225:data<=16'd15009;
      120226:data<=16'd15887;
      120227:data<=16'd16722;
      120228:data<=16'd15961;
      120229:data<=16'd15556;
      120230:data<=16'd14918;
      120231:data<=16'd13770;
      120232:data<=16'd14284;
      120233:data<=16'd15470;
      120234:data<=16'd15283;
      120235:data<=16'd14176;
      120236:data<=16'd15189;
      120237:data<=16'd17493;
      120238:data<=16'd16522;
      120239:data<=16'd15847;
      120240:data<=16'd17161;
      120241:data<=16'd15649;
      120242:data<=16'd14765;
      120243:data<=16'd14615;
      120244:data<=16'd12163;
      120245:data<=16'd12980;
      120246:data<=16'd13908;
      120247:data<=16'd12568;
      120248:data<=16'd14439;
      120249:data<=16'd9976;
      120250:data<=-16'd1804;
      120251:data<=-16'd4811;
      120252:data<=-16'd1700;
      120253:data<=-16'd1048;
      120254:data<=-16'd876;
      120255:data<=-16'd1585;
      120256:data<=-16'd1991;
      120257:data<=-16'd1513;
      120258:data<=-16'd1820;
      120259:data<=-16'd587;
      120260:data<=16'd490;
      120261:data<=-16'd284;
      120262:data<=-16'd309;
      120263:data<=-16'd628;
      120264:data<=-16'd943;
      120265:data<=-16'd381;
      120266:data<=-16'd726;
      120267:data<=-16'd764;
      120268:data<=-16'd816;
      120269:data<=-16'd1868;
      120270:data<=-16'd1750;
      120271:data<=-16'd1413;
      120272:data<=-16'd2378;
      120273:data<=-16'd3664;
      120274:data<=-16'd4426;
      120275:data<=-16'd4358;
      120276:data<=-16'd4540;
      120277:data<=-16'd4552;
      120278:data<=-16'd4464;
      120279:data<=-16'd5817;
      120280:data<=-16'd5887;
      120281:data<=-16'd5101;
      120282:data<=-16'd6146;
      120283:data<=-16'd5817;
      120284:data<=-16'd4730;
      120285:data<=-16'd4998;
      120286:data<=-16'd6429;
      120287:data<=-16'd10411;
      120288:data<=-16'd10910;
      120289:data<=-16'd8294;
      120290:data<=-16'd10722;
      120291:data<=-16'd7386;
      120292:data<=16'd3923;
      120293:data<=16'd5794;
      120294:data<=16'd2849;
      120295:data<=16'd4272;
      120296:data<=16'd3818;
      120297:data<=16'd3303;
      120298:data<=16'd3641;
      120299:data<=16'd1533;
      120300:data<=16'd957;
      120301:data<=16'd1345;
      120302:data<=16'd870;
      120303:data<=16'd1192;
      120304:data<=16'd751;
      120305:data<=16'd15;
      120306:data<=-16'd734;
      120307:data<=-16'd1753;
      120308:data<=-16'd936;
      120309:data<=-16'd752;
      120310:data<=-16'd1650;
      120311:data<=-16'd1221;
      120312:data<=-16'd2108;
      120313:data<=-16'd3303;
      120314:data<=-16'd2566;
      120315:data<=-16'd2490;
      120316:data<=-16'd2713;
      120317:data<=-16'd2300;
      120318:data<=-16'd2375;
      120319:data<=-16'd3134;
      120320:data<=-16'd3997;
      120321:data<=-16'd3812;
      120322:data<=-16'd3894;
      120323:data<=-16'd4197;
      120324:data<=-16'd3127;
      120325:data<=-16'd3877;
      120326:data<=-16'd5703;
      120327:data<=-16'd5756;
      120328:data<=-16'd6199;
      120329:data<=-16'd5714;
      120330:data<=-16'd5172;
      120331:data<=-16'd5997;
      120332:data<=-16'd4716;
      120333:data<=-16'd8812;
      120334:data<=-16'd20131;
      120335:data<=-16'd23479;
      120336:data<=-16'd18933;
      120337:data<=-16'd15954;
      120338:data<=-16'd14551;
      120339:data<=-16'd15585;
      120340:data<=-16'd16792;
      120341:data<=-16'd15259;
      120342:data<=-16'd14319;
      120343:data<=-16'd13729;
      120344:data<=-16'd13327;
      120345:data<=-16'd14317;
      120346:data<=-16'd14386;
      120347:data<=-16'd13735;
      120348:data<=-16'd12979;
      120349:data<=-16'd12193;
      120350:data<=-16'd12163;
      120351:data<=-16'd11571;
      120352:data<=-16'd11837;
      120353:data<=-16'd12875;
      120354:data<=-16'd11647;
      120355:data<=-16'd10778;
      120356:data<=-16'd10818;
      120357:data<=-16'd9784;
      120358:data<=-16'd10058;
      120359:data<=-16'd11189;
      120360:data<=-16'd11342;
      120361:data<=-16'd10739;
      120362:data<=-16'd9777;
      120363:data<=-16'd9565;
      120364:data<=-16'd8910;
      120365:data<=-16'd8686;
      120366:data<=-16'd10052;
      120367:data<=-16'd9121;
      120368:data<=-16'd7867;
      120369:data<=-16'd8108;
      120370:data<=-16'd6730;
      120371:data<=-16'd6769;
      120372:data<=-16'd6661;
      120373:data<=-16'd5025;
      120374:data<=-16'd6858;
      120375:data<=-16'd2716;
      120376:data<=16'd9192;
      120377:data<=16'd12193;
      120378:data<=16'd9817;
      120379:data<=16'd11708;
      120380:data<=16'd12044;
      120381:data<=16'd11447;
      120382:data<=16'd12383;
      120383:data<=16'd11612;
      120384:data<=16'd10980;
      120385:data<=16'd11952;
      120386:data<=16'd11937;
      120387:data<=16'd9752;
      120388:data<=16'd7847;
      120389:data<=16'd8022;
      120390:data<=16'd7956;
      120391:data<=16'd8275;
      120392:data<=16'd9633;
      120393:data<=16'd9094;
      120394:data<=16'd8839;
      120395:data<=16'd9899;
      120396:data<=16'd9310;
      120397:data<=16'd8523;
      120398:data<=16'd8566;
      120399:data<=16'd9250;
      120400:data<=16'd10322;
      120401:data<=16'd9943;
      120402:data<=16'd9715;
      120403:data<=16'd9696;
      120404:data<=16'd8702;
      120405:data<=16'd9476;
      120406:data<=16'd10147;
      120407:data<=16'd9085;
      120408:data<=16'd8971;
      120409:data<=16'd8637;
      120410:data<=16'd8241;
      120411:data<=16'd8338;
      120412:data<=16'd8170;
      120413:data<=16'd9436;
      120414:data<=16'd9091;
      120415:data<=16'd7949;
      120416:data<=16'd9853;
      120417:data<=16'd5369;
      120418:data<=-16'd5028;
      120419:data<=-16'd7097;
      120420:data<=-16'd4394;
      120421:data<=-16'd4901;
      120422:data<=-16'd5080;
      120423:data<=-16'd4582;
      120424:data<=-16'd4676;
      120425:data<=-16'd3900;
      120426:data<=-16'd2504;
      120427:data<=-16'd1706;
      120428:data<=-16'd1923;
      120429:data<=-16'd1970;
      120430:data<=-16'd1812;
      120431:data<=-16'd1501;
      120432:data<=16'd14;
      120433:data<=16'd561;
      120434:data<=16'd2;
      120435:data<=16'd578;
      120436:data<=16'd1122;
      120437:data<=16'd2563;
      120438:data<=16'd5184;
      120439:data<=16'd6296;
      120440:data<=16'd6649;
      120441:data<=16'd6050;
      120442:data<=16'd4755;
      120443:data<=16'd5074;
      120444:data<=16'd5145;
      120445:data<=16'd5316;
      120446:data<=16'd6378;
      120447:data<=16'd5800;
      120448:data<=16'd6020;
      120449:data<=16'd6843;
      120450:data<=16'd5624;
      120451:data<=16'd5985;
      120452:data<=16'd7215;
      120453:data<=16'd7368;
      120454:data<=16'd7796;
      120455:data<=16'd6228;
      120456:data<=16'd5482;
      120457:data<=16'd6708;
      120458:data<=16'd5380;
      120459:data<=16'd9222;
      120460:data<=16'd19572;
      120461:data<=16'd22789;
      120462:data<=16'd20494;
      120463:data<=16'd20016;
      120464:data<=16'd18900;
      120465:data<=16'd18683;
      120466:data<=16'd19848;
      120467:data<=16'd19085;
      120468:data<=16'd17858;
      120469:data<=16'd16715;
      120470:data<=16'd15420;
      120471:data<=16'd15643;
      120472:data<=16'd16498;
      120473:data<=16'd16190;
      120474:data<=16'd14690;
      120475:data<=16'd13738;
      120476:data<=16'd13715;
      120477:data<=16'd12778;
      120478:data<=16'd11947;
      120479:data<=16'd11621;
      120480:data<=16'd10173;
      120481:data<=16'd9371;
      120482:data<=16'd9412;
      120483:data<=16'd8789;
      120484:data<=16'd8305;
      120485:data<=16'd6963;
      120486:data<=16'd4541;
      120487:data<=16'd2203;
      120488:data<=-16'd297;
      120489:data<=-16'd1151;
      120490:data<=-16'd790;
      120491:data<=-16'd1873;
      120492:data<=-16'd3004;
      120493:data<=-16'd3685;
      120494:data<=-16'd4537;
      120495:data<=-16'd4930;
      120496:data<=-16'd4984;
      120497:data<=-16'd4408;
      120498:data<=-16'd5530;
      120499:data<=-16'd7650;
      120500:data<=-16'd6420;
      120501:data<=-16'd9200;
      120502:data<=-16'd18895;
      120503:data<=-16'd22920;
      120504:data<=-16'd21538;
      120505:data<=-16'd22344;
      120506:data<=-16'd22143;
      120507:data<=-16'd21187;
      120508:data<=-16'd21688;
      120509:data<=-16'd21141;
      120510:data<=-16'd20007;
      120511:data<=-16'd19707;
      120512:data<=-16'd20454;
      120513:data<=-16'd20982;
      120514:data<=-16'd19854;
      120515:data<=-16'd19047;
      120516:data<=-16'd18258;
      120517:data<=-16'd17167;
      120518:data<=-16'd18277;
      120519:data<=-16'd18945;
      120520:data<=-16'd17644;
      120521:data<=-16'd17161;
      120522:data<=-16'd16780;
      120523:data<=-16'd15949;
      120524:data<=-16'd15702;
      120525:data<=-16'd16390;
      120526:data<=-16'd17223;
      120527:data<=-16'd16214;
      120528:data<=-16'd15274;
      120529:data<=-16'd14997;
      120530:data<=-16'd13309;
      120531:data<=-16'd13749;
      120532:data<=-16'd15568;
      120533:data<=-16'd14604;
      120534:data<=-16'd13903;
      120535:data<=-16'd13449;
      120536:data<=-16'd11359;
      120537:data<=-16'd9273;
      120538:data<=-16'd7577;
      120539:data<=-16'd8019;
      120540:data<=-16'd8301;
      120541:data<=-16'd6939;
      120542:data<=-16'd8507;
      120543:data<=-16'd5580;
      120544:data<=16'd4631;
      120545:data<=16'd7808;
      120546:data<=16'd5369;
      120547:data<=16'd5883;
      120548:data<=16'd5635;
      120549:data<=16'd5359;
      120550:data<=16'd6044;
      120551:data<=16'd5024;
      120552:data<=16'd4014;
      120553:data<=16'd3125;
      120554:data<=16'd2886;
      120555:data<=16'd3600;
      120556:data<=16'd3072;
      120557:data<=16'd2564;
      120558:data<=16'd1269;
      120559:data<=-16'd687;
      120560:data<=16'd262;
      120561:data<=16'd1019;
      120562:data<=16'd532;
      120563:data<=16'd1219;
      120564:data<=16'd370;
      120565:data<=-16'd1172;
      120566:data<=-16'd1333;
      120567:data<=-16'd1363;
      120568:data<=-16'd848;
      120569:data<=-16'd684;
      120570:data<=-16'd966;
      120571:data<=-16'd1343;
      120572:data<=-16'd2877;
      120573:data<=-16'd3033;
      120574:data<=-16'd2649;
      120575:data<=-16'd3676;
      120576:data<=-16'd2867;
      120577:data<=-16'd2355;
      120578:data<=-16'd4018;
      120579:data<=-16'd4708;
      120580:data<=-16'd4936;
      120581:data<=-16'd4308;
      120582:data<=-16'd3579;
      120583:data<=-16'd4120;
      120584:data<=-16'd2939;
      120585:data<=-16'd5125;
      120586:data<=-16'd14123;
      120587:data<=-16'd20231;
      120588:data<=-16'd20918;
      120589:data<=-16'd20609;
      120590:data<=-16'd19575;
      120591:data<=-16'd18187;
      120592:data<=-16'd16081;
      120593:data<=-16'd14631;
      120594:data<=-16'd14998;
      120595:data<=-16'd13917;
      120596:data<=-16'd12326;
      120597:data<=-16'd11761;
      120598:data<=-16'd10149;
      120599:data<=-16'd8733;
      120600:data<=-16'd7975;
      120601:data<=-16'd6998;
      120602:data<=-16'd6730;
      120603:data<=-16'd6393;
      120604:data<=-16'd5412;
      120605:data<=-16'd3994;
      120606:data<=-16'd2863;
      120607:data<=-16'd2911;
      120608:data<=-16'd2328;
      120609:data<=-16'd1610;
      120610:data<=-16'd1765;
      120611:data<=-16'd607;
      120612:data<=16'd291;
      120613:data<=16'd294;
      120614:data<=16'd1242;
      120615:data<=16'd1172;
      120616:data<=16'd1022;
      120617:data<=16'd2255;
      120618:data<=16'd2974;
      120619:data<=16'd3894;
      120620:data<=16'd4460;
      120621:data<=16'd4589;
      120622:data<=16'd5363;
      120623:data<=16'd4420;
      120624:data<=16'd4928;
      120625:data<=16'd7738;
      120626:data<=16'd6438;
      120627:data<=16'd7671;
      120628:data<=16'd16763;
      120629:data<=16'd21983;
      120630:data<=16'd20776;
      120631:data<=16'd20862;
      120632:data<=16'd21667;
      120633:data<=16'd20783;
      120634:data<=16'd19787;
      120635:data<=16'd19420;
      120636:data<=16'd18921;
      120637:data<=16'd19923;
      120638:data<=16'd23309;
      120639:data<=16'd24310;
      120640:data<=16'd22598;
      120641:data<=16'd22319;
      120642:data<=16'd21279;
      120643:data<=16'd19484;
      120644:data<=16'd20096;
      120645:data<=16'd20466;
      120646:data<=16'd19425;
      120647:data<=16'd18548;
      120648:data<=16'd17770;
      120649:data<=16'd17356;
      120650:data<=16'd16909;
      120651:data<=16'd17139;
      120652:data<=16'd17946;
      120653:data<=16'd16901;
      120654:data<=16'd15938;
      120655:data<=16'd15867;
      120656:data<=16'd14449;
      120657:data<=16'd14075;
      120658:data<=16'd14906;
      120659:data<=16'd14402;
      120660:data<=16'd13555;
      120661:data<=16'd12646;
      120662:data<=16'd12108;
      120663:data<=16'd11846;
      120664:data<=16'd11045;
      120665:data<=16'd11896;
      120666:data<=16'd11958;
      120667:data<=16'd9846;
      120668:data<=16'd10962;
      120669:data<=16'd9815;
      120670:data<=16'd848;
      120671:data<=-16'd4886;
      120672:data<=-16'd3677;
      120673:data<=-16'd3212;
      120674:data<=-16'd3574;
      120675:data<=-16'd3021;
      120676:data<=-16'd3110;
      120677:data<=-16'd2989;
      120678:data<=-16'd1947;
      120679:data<=-16'd1398;
      120680:data<=-16'd1613;
      120681:data<=-16'd1366;
      120682:data<=-16'd1034;
      120683:data<=-16'd1245;
      120684:data<=-16'd693;
      120685:data<=16'd444;
      120686:data<=16'd945;
      120687:data<=16'd12;
      120688:data<=-16'd2754;
      120689:data<=-16'd4303;
      120690:data<=-16'd3562;
      120691:data<=-16'd3644;
      120692:data<=-16'd3861;
      120693:data<=-16'd3682;
      120694:data<=-16'd4454;
      120695:data<=-16'd4429;
      120696:data<=-16'd4137;
      120697:data<=-16'd4610;
      120698:data<=-16'd4761;
      120699:data<=-16'd5600;
      120700:data<=-16'd5702;
      120701:data<=-16'd4669;
      120702:data<=-16'd5248;
      120703:data<=-16'd5046;
      120704:data<=-16'd4743;
      120705:data<=-16'd6910;
      120706:data<=-16'd6863;
      120707:data<=-16'd5726;
      120708:data<=-16'd6429;
      120709:data<=-16'd5688;
      120710:data<=-16'd6488;
      120711:data<=-16'd7216;
      120712:data<=-16'd52;
      120713:data<=16'd7253;
      120714:data<=16'd7006;
      120715:data<=16'd5909;
      120716:data<=16'd6511;
      120717:data<=16'd5730;
      120718:data<=16'd3914;
      120719:data<=16'd2878;
      120720:data<=16'd3106;
      120721:data<=16'd3112;
      120722:data<=16'd3043;
      120723:data<=16'd3310;
      120724:data<=16'd1809;
      120725:data<=-16'd121;
      120726:data<=-16'd182;
      120727:data<=-16'd94;
      120728:data<=-16'd358;
      120729:data<=-16'd273;
      120730:data<=-16'd623;
      120731:data<=-16'd1560;
      120732:data<=-16'd2228;
      120733:data<=-16'd2202;
      120734:data<=-16'd2375;
      120735:data<=-16'd2739;
      120736:data<=-16'd2209;
      120737:data<=-16'd1438;
      120738:data<=-16'd569;
      120739:data<=16'd209;
      120740:data<=-16'd277;
      120741:data<=-16'd435;
      120742:data<=-16'd49;
      120743:data<=-16'd1027;
      120744:data<=-16'd2206;
      120745:data<=-16'd3113;
      120746:data<=-16'd3603;
      120747:data<=-16'd3110;
      120748:data<=-16'd3676;
      120749:data<=-16'd3938;
      120750:data<=-16'd3321;
      120751:data<=-16'd5288;
      120752:data<=-16'd5723;
      120753:data<=-16'd4699;
      120754:data<=-16'd11435;
      120755:data<=-16'd19511;
      120756:data<=-16'd19233;
      120757:data<=-16'd18475;
      120758:data<=-16'd20295;
      120759:data<=-16'd19299;
      120760:data<=-16'd18042;
      120761:data<=-16'd18154;
      120762:data<=-16'd17094;
      120763:data<=-16'd16143;
      120764:data<=-16'd16587;
      120765:data<=-16'd17183;
      120766:data<=-16'd16600;
      120767:data<=-16'd15500;
      120768:data<=-16'd15341;
      120769:data<=-16'd14531;
      120770:data<=-16'd13277;
      120771:data<=-16'd14098;
      120772:data<=-16'd14698;
      120773:data<=-16'd13926;
      120774:data<=-16'd13869;
      120775:data<=-16'd12945;
      120776:data<=-16'd11273;
      120777:data<=-16'd11831;
      120778:data<=-16'd13244;
      120779:data<=-16'd12966;
      120780:data<=-16'd11803;
      120781:data<=-16'd11403;
      120782:data<=-16'd11083;
      120783:data<=-16'd10348;
      120784:data<=-16'd10845;
      120785:data<=-16'd10904;
      120786:data<=-16'd9439;
      120787:data<=-16'd10373;
      120788:data<=-16'd12568;
      120789:data<=-16'd12361;
      120790:data<=-16'd11694;
      120791:data<=-16'd12138;
      120792:data<=-16'd12625;
      120793:data<=-16'd11491;
      120794:data<=-16'd10320;
      120795:data<=-16'd10631;
      120796:data<=-16'd5002;
      120797:data<=16'd5145;
      120798:data<=16'd7080;
      120799:data<=16'd4986;
      120800:data<=16'd6337;
      120801:data<=16'd6070;
      120802:data<=16'd5661;
      120803:data<=16'd7175;
      120804:data<=16'd7423;
      120805:data<=16'd7874;
      120806:data<=16'd8088;
      120807:data<=16'd7808;
      120808:data<=16'd8608;
      120809:data<=16'd8140;
      120810:data<=16'd8084;
      120811:data<=16'd9652;
      120812:data<=16'd9442;
      120813:data<=16'd8942;
      120814:data<=16'd9216;
      120815:data<=16'd9115;
      120816:data<=16'd9411;
      120817:data<=16'd9615;
      120818:data<=16'd10261;
      120819:data<=16'd10877;
      120820:data<=16'd10326;
      120821:data<=16'd10618;
      120822:data<=16'd10633;
      120823:data<=16'd10072;
      120824:data<=16'd11110;
      120825:data<=16'd11455;
      120826:data<=16'd10922;
      120827:data<=16'd10739;
      120828:data<=16'd10008;
      120829:data<=16'd9831;
      120830:data<=16'd9774;
      120831:data<=16'd10285;
      120832:data<=16'd11200;
      120833:data<=16'd9982;
      120834:data<=16'd10103;
      120835:data<=16'd10128;
      120836:data<=16'd8035;
      120837:data<=16'd11221;
      120838:data<=16'd11121;
      120839:data<=16'd1119;
      120840:data<=-16'd1898;
      120841:data<=16'd1371;
      120842:data<=16'd32;
      120843:data<=16'd344;
      120844:data<=16'd1924;
      120845:data<=16'd1392;
      120846:data<=16'd2036;
      120847:data<=16'd2029;
      120848:data<=16'd1685;
      120849:data<=16'd1879;
      120850:data<=16'd1754;
      120851:data<=16'd3668;
      120852:data<=16'd4693;
      120853:data<=16'd3636;
      120854:data<=16'd3991;
      120855:data<=16'd3711;
      120856:data<=16'd3280;
      120857:data<=16'd4363;
      120858:data<=16'd4514;
      120859:data<=16'd4499;
      120860:data<=16'd4745;
      120861:data<=16'd4378;
      120862:data<=16'd4056;
      120863:data<=16'd4306;
      120864:data<=16'd5830;
      120865:data<=16'd6175;
      120866:data<=16'd5127;
      120867:data<=16'd5574;
      120868:data<=16'd4951;
      120869:data<=16'd4481;
      120870:data<=16'd6572;
      120871:data<=16'd7028;
      120872:data<=16'd6711;
      120873:data<=16'd6643;
      120874:data<=16'd6023;
      120875:data<=16'd6895;
      120876:data<=16'd6391;
      120877:data<=16'd6673;
      120878:data<=16'd8795;
      120879:data<=16'd6217;
      120880:data<=16'd9414;
      120881:data<=16'd20709;
      120882:data<=16'd21713;
      120883:data<=16'd18448;
      120884:data<=16'd21082;
      120885:data<=16'd20697;
      120886:data<=16'd19324;
      120887:data<=16'd19015;
      120888:data<=16'd15212;
      120889:data<=16'd12766;
      120890:data<=16'd13150;
      120891:data<=16'd13709;
      120892:data<=16'd13678;
      120893:data<=16'd12220;
      120894:data<=16'd11952;
      120895:data<=16'd11706;
      120896:data<=16'd10527;
      120897:data<=16'd11668;
      120898:data<=16'd11743;
      120899:data<=16'd10430;
      120900:data<=16'd10983;
      120901:data<=16'd10158;
      120902:data<=16'd8815;
      120903:data<=16'd9039;
      120904:data<=16'd8780;
      120905:data<=16'd8387;
      120906:data<=16'd7565;
      120907:data<=16'd6775;
      120908:data<=16'd6786;
      120909:data<=16'd6240;
      120910:data<=16'd5650;
      120911:data<=16'd3723;
      120912:data<=16'd1503;
      120913:data<=16'd1780;
      120914:data<=16'd1089;
      120915:data<=16'd400;
      120916:data<=16'd367;
      120917:data<=-16'd2261;
      120918:data<=-16'd2514;
      120919:data<=-16'd2457;
      120920:data<=-16'd4981;
      120921:data<=-16'd2819;
      120922:data<=-16'd5332;
      120923:data<=-16'd16948;
      120924:data<=-16'd20572;
      120925:data<=-16'd18299;
      120926:data<=-16'd19558;
      120927:data<=-16'd19528;
      120928:data<=-16'd18672;
      120929:data<=-16'd18120;
      120930:data<=-16'd17515;
      120931:data<=-16'd18801;
      120932:data<=-16'd18528;
      120933:data<=-16'd17652;
      120934:data<=-16'd18265;
      120935:data<=-16'd17089;
      120936:data<=-16'd16756;
      120937:data<=-16'd17529;
      120938:data<=-16'd15523;
      120939:data<=-16'd13349;
      120940:data<=-16'd12686;
      120941:data<=-16'd12422;
      120942:data<=-16'd11993;
      120943:data<=-16'd11743;
      120944:data<=-16'd13279;
      120945:data<=-16'd13894;
      120946:data<=-16'd12798;
      120947:data<=-16'd12924;
      120948:data<=-16'd11938;
      120949:data<=-16'd10845;
      120950:data<=-16'd12652;
      120951:data<=-16'd13549;
      120952:data<=-16'd12652;
      120953:data<=-16'd11765;
      120954:data<=-16'd11119;
      120955:data<=-16'd11312;
      120956:data<=-16'd11342;
      120957:data<=-16'd12029;
      120958:data<=-16'd12525;
      120959:data<=-16'd11092;
      120960:data<=-16'd11682;
      120961:data<=-16'd11576;
      120962:data<=-16'd9172;
      120963:data<=-16'd11166;
      120964:data<=-16'd8866;
      120965:data<=16'd1903;
      120966:data<=16'd4861;
      120967:data<=16'd1642;
      120968:data<=16'd3075;
      120969:data<=16'd3697;
      120970:data<=16'd2196;
      120971:data<=16'd2011;
      120972:data<=16'd1528;
      120973:data<=16'd1078;
      120974:data<=16'd1002;
      120975:data<=16'd1384;
      120976:data<=16'd1501;
      120977:data<=-16'd209;
      120978:data<=-16'd895;
      120979:data<=-16'd540;
      120980:data<=-16'd1113;
      120981:data<=-16'd381;
      120982:data<=-16'd35;
      120983:data<=-16'd1471;
      120984:data<=-16'd2030;
      120985:data<=-16'd2479;
      120986:data<=-16'd2552;
      120987:data<=-16'd2059;
      120988:data<=-16'd3718;
      120989:data<=-16'd6041;
      120990:data<=-16'd7241;
      120991:data<=-16'd7752;
      120992:data<=-16'd7166;
      120993:data<=-16'd6772;
      120994:data<=-16'd6833;
      120995:data<=-16'd6542;
      120996:data<=-16'd6868;
      120997:data<=-16'd7888;
      120998:data<=-16'd8645;
      120999:data<=-16'd8046;
      121000:data<=-16'd7553;
      121001:data<=-16'd8093;
      121002:data<=-16'd6857;
      121003:data<=-16'd7321;
      121004:data<=-16'd9809;
      121005:data<=-16'd7559;
      121006:data<=-16'd9867;
      121007:data<=-16'd20550;
      121008:data<=-16'd22959;
      121009:data<=-16'd19423;
      121010:data<=-16'd20237;
      121011:data<=-16'd19167;
      121012:data<=-16'd17338;
      121013:data<=-16'd18008;
      121014:data<=-16'd16732;
      121015:data<=-16'd15535;
      121016:data<=-16'd14912;
      121017:data<=-16'd12760;
      121018:data<=-16'd11400;
      121019:data<=-16'd10652;
      121020:data<=-16'd10140;
      121021:data<=-16'd9981;
      121022:data<=-16'd9048;
      121023:data<=-16'd7820;
      121024:data<=-16'd5874;
      121025:data<=-16'd4766;
      121026:data<=-16'd5521;
      121027:data<=-16'd4954;
      121028:data<=-16'd4062;
      121029:data<=-16'd3404;
      121030:data<=-16'd1350;
      121031:data<=-16'd584;
      121032:data<=-16'd446;
      121033:data<=16'd235;
      121034:data<=-16'd553;
      121035:data<=-16'd678;
      121036:data<=16'd509;
      121037:data<=16'd2026;
      121038:data<=16'd4792;
      121039:data<=16'd7368;
      121040:data<=16'd8862;
      121041:data<=16'd8384;
      121042:data<=16'd7407;
      121043:data<=16'd9321;
      121044:data<=16'd10043;
      121045:data<=16'd9539;
      121046:data<=16'd10616;
      121047:data<=16'd9138;
      121048:data<=16'd12304;
      121049:data<=16'd23132;
      121050:data<=16'd26621;
      121051:data<=16'd24065;
      121052:data<=16'd24400;
      121053:data<=16'd23962;
      121054:data<=16'd23329;
      121055:data<=16'd23044;
      121056:data<=16'd22231;
      121057:data<=16'd23375;
      121058:data<=16'd22795;
      121059:data<=16'd21124;
      121060:data<=16'd21696;
      121061:data<=16'd20447;
      121062:data<=16'd19359;
      121063:data<=16'd20724;
      121064:data<=16'd20909;
      121065:data<=16'd20735;
      121066:data<=16'd20202;
      121067:data<=16'd18844;
      121068:data<=16'd18316;
      121069:data<=16'd17741;
      121070:data<=16'd18037;
      121071:data<=16'd18776;
      121072:data<=16'd17987;
      121073:data<=16'd17518;
      121074:data<=16'd16724;
      121075:data<=16'd15458;
      121076:data<=16'd16067;
      121077:data<=16'd16906;
      121078:data<=16'd16466;
      121079:data<=16'd15089;
      121080:data<=16'd14160;
      121081:data<=16'd13793;
      121082:data<=16'd12063;
      121083:data<=16'd12536;
      121084:data<=16'd14357;
      121085:data<=16'd12307;
      121086:data<=16'd12114;
      121087:data<=16'd12913;
      121088:data<=16'd9321;
      121089:data<=16'd8011;
      121090:data<=16'd4805;
      121091:data<=-16'd4883;
      121092:data<=-16'd8351;
      121093:data<=-16'd6288;
      121094:data<=-16'd7122;
      121095:data<=-16'd7227;
      121096:data<=-16'd5994;
      121097:data<=-16'd5046;
      121098:data<=-16'd4355;
      121099:data<=-16'd4695;
      121100:data<=-16'd3905;
      121101:data<=-16'd3336;
      121102:data<=-16'd4088;
      121103:data<=-16'd3178;
      121104:data<=-16'd2608;
      121105:data<=-16'd3062;
      121106:data<=-16'd2734;
      121107:data<=-16'd3368;
      121108:data<=-16'd3667;
      121109:data<=-16'd2120;
      121110:data<=-16'd760;
      121111:data<=-16'd382;
      121112:data<=-16'd701;
      121113:data<=-16'd632;
      121114:data<=-16'd679;
      121115:data<=-16'd1512;
      121116:data<=-16'd1334;
      121117:data<=-16'd1545;
      121118:data<=-16'd2300;
      121119:data<=-16'd1199;
      121120:data<=-16'd816;
      121121:data<=-16'd1521;
      121122:data<=-16'd1569;
      121123:data<=-16'd2522;
      121124:data<=-16'd3133;
      121125:data<=-16'd2996;
      121126:data<=-16'd3207;
      121127:data<=-16'd2849;
      121128:data<=-16'd3347;
      121129:data<=-16'd3767;
      121130:data<=-16'd4344;
      121131:data<=-16'd6977;
      121132:data<=-16'd2817;
      121133:data<=16'd7685;
      121134:data<=16'd10545;
      121135:data<=16'd8849;
      121136:data<=16'd8593;
      121137:data<=16'd5994;
      121138:data<=16'd6273;
      121139:data<=16'd9875;
      121140:data<=16'd9580;
      121141:data<=16'd8786;
      121142:data<=16'd8634;
      121143:data<=16'd6388;
      121144:data<=16'd5927;
      121145:data<=16'd6540;
      121146:data<=16'd5109;
      121147:data<=16'd4419;
      121148:data<=16'd5142;
      121149:data<=16'd4622;
      121150:data<=16'd2493;
      121151:data<=16'd1125;
      121152:data<=16'd1368;
      121153:data<=16'd1406;
      121154:data<=16'd1556;
      121155:data<=16'd1677;
      121156:data<=16'd5;
      121157:data<=-16'd1221;
      121158:data<=-16'd666;
      121159:data<=-16'd569;
      121160:data<=-16'd1024;
      121161:data<=-16'd1240;
      121162:data<=-16'd1653;
      121163:data<=-16'd2740;
      121164:data<=-16'd3680;
      121165:data<=-16'd3842;
      121166:data<=-16'd4705;
      121167:data<=-16'd4780;
      121168:data<=-16'd3268;
      121169:data<=-16'd4328;
      121170:data<=-16'd6423;
      121171:data<=-16'd6675;
      121172:data<=-16'd6754;
      121173:data<=-16'd5823;
      121174:data<=-16'd8577;
      121175:data<=-16'd17976;
      121176:data<=-16'd22944;
      121177:data<=-16'd21505;
      121178:data<=-16'd21391;
      121179:data<=-16'd21268;
      121180:data<=-16'd20002;
      121181:data<=-16'd18806;
      121182:data<=-16'd18016;
      121183:data<=-16'd19059;
      121184:data<=-16'd18998;
      121185:data<=-16'd17814;
      121186:data<=-16'd18124;
      121187:data<=-16'd16866;
      121188:data<=-16'd16354;
      121189:data<=-16'd19672;
      121190:data<=-16'd21792;
      121191:data<=-16'd21441;
      121192:data<=-16'd20316;
      121193:data<=-16'd18989;
      121194:data<=-16'd18513;
      121195:data<=-16'd18061;
      121196:data<=-16'd18211;
      121197:data<=-16'd18310;
      121198:data<=-16'd16824;
      121199:data<=-16'd16615;
      121200:data<=-16'd16536;
      121201:data<=-16'd14839;
      121202:data<=-16'd14727;
      121203:data<=-16'd15167;
      121204:data<=-16'd15013;
      121205:data<=-16'd15036;
      121206:data<=-16'd13903;
      121207:data<=-16'd12498;
      121208:data<=-16'd11244;
      121209:data<=-16'd11045;
      121210:data<=-16'd12381;
      121211:data<=-16'd11664;
      121212:data<=-16'd10862;
      121213:data<=-16'd10956;
      121214:data<=-16'd9245;
      121215:data<=-16'd9791;
      121216:data<=-16'd7715;
      121217:data<=16'd1933;
      121218:data<=16'd6340;
      121219:data<=16'd4648;
      121220:data<=16'd5915;
      121221:data<=16'd6278;
      121222:data<=16'd5315;
      121223:data<=16'd5797;
      121224:data<=16'd5739;
      121225:data<=16'd6067;
      121226:data<=16'd6141;
      121227:data<=16'd5491;
      121228:data<=16'd5856;
      121229:data<=16'd6578;
      121230:data<=16'd7943;
      121231:data<=16'd8633;
      121232:data<=16'd8143;
      121233:data<=16'd8818;
      121234:data<=16'd8677;
      121235:data<=16'd8792;
      121236:data<=16'd10787;
      121237:data<=16'd10428;
      121238:data<=16'd10473;
      121239:data<=16'd13154;
      121240:data<=16'd13526;
      121241:data<=16'd13186;
      121242:data<=16'd14314;
      121243:data<=16'd14938;
      121244:data<=16'd14804;
      121245:data<=16'd13635;
      121246:data<=16'd13189;
      121247:data<=16'd13517;
      121248:data<=16'd12581;
      121249:data<=16'd13019;
      121250:data<=16'd14013;
      121251:data<=16'd12948;
      121252:data<=16'd12431;
      121253:data<=16'd12245;
      121254:data<=16'd11550;
      121255:data<=16'd11461;
      121256:data<=16'd11953;
      121257:data<=16'd13265;
      121258:data<=16'd10323;
      121259:data<=16'd1354;
      121260:data<=-16'd3970;
      121261:data<=-16'd3735;
      121262:data<=-16'd3062;
      121263:data<=-16'd1497;
      121264:data<=-16'd566;
      121265:data<=-16'd1081;
      121266:data<=-16'd836;
      121267:data<=-16'd1040;
      121268:data<=-16'd870;
      121269:data<=16'd622;
      121270:data<=16'd1078;
      121271:data<=16'd1328;
      121272:data<=16'd1880;
      121273:data<=16'd1454;
      121274:data<=16'd1051;
      121275:data<=16'd1209;
      121276:data<=16'd2270;
      121277:data<=16'd3583;
      121278:data<=16'd3465;
      121279:data<=16'd3424;
      121280:data<=16'd3397;
      121281:data<=16'd2267;
      121282:data<=16'd3102;
      121283:data<=16'd5128;
      121284:data<=16'd4737;
      121285:data<=16'd3765;
      121286:data<=16'd3751;
      121287:data<=16'd3600;
      121288:data<=16'd3115;
      121289:data<=16'd2126;
      121290:data<=16'd1146;
      121291:data<=16'd1046;
      121292:data<=16'd1606;
      121293:data<=16'd1694;
      121294:data<=16'd1034;
      121295:data<=16'd1668;
      121296:data<=16'd3248;
      121297:data<=16'd3827;
      121298:data<=16'd4046;
      121299:data<=16'd3121;
      121300:data<=16'd4416;
      121301:data<=16'd12930;
      121302:data<=16'd19837;
      121303:data<=16'd19103;
      121304:data<=16'd18325;
      121305:data<=16'd18201;
      121306:data<=16'd16803;
      121307:data<=16'd16754;
      121308:data<=16'd16239;
      121309:data<=16'd15690;
      121310:data<=16'd16202;
      121311:data<=16'd15355;
      121312:data<=16'd15097;
      121313:data<=16'd14904;
      121314:data<=16'd13019;
      121315:data<=16'd13397;
      121316:data<=16'd14821;
      121317:data<=16'd14277;
      121318:data<=16'd13778;
      121319:data<=16'd13418;
      121320:data<=16'd12683;
      121321:data<=16'd11576;
      121322:data<=16'd11092;
      121323:data<=16'd12604;
      121324:data<=16'd12486;
      121325:data<=16'd10819;
      121326:data<=16'd11326;
      121327:data<=16'd10892;
      121328:data<=16'd9066;
      121329:data<=16'd8587;
      121330:data<=16'd7903;
      121331:data<=16'd7700;
      121332:data<=16'd7926;
      121333:data<=16'd6496;
      121334:data<=16'd5485;
      121335:data<=16'd5316;
      121336:data<=16'd3844;
      121337:data<=16'd1767;
      121338:data<=16'd1431;
      121339:data<=16'd3142;
      121340:data<=16'd4701;
      121341:data<=16'd5733;
      121342:data<=16'd3156;
      121343:data<=-16'd6643;
      121344:data<=-16'd14038;
      121345:data<=-16'd13030;
      121346:data<=-16'd12440;
      121347:data<=-16'd13254;
      121348:data<=-16'd12446;
      121349:data<=-16'd13318;
      121350:data<=-16'd14170;
      121351:data<=-16'd13415;
      121352:data<=-16'd13142;
      121353:data<=-16'd12649;
      121354:data<=-16'd12192;
      121355:data<=-16'd12402;
      121356:data<=-16'd13253;
      121357:data<=-16'd14396;
      121358:data<=-16'd13931;
      121359:data<=-16'd13432;
      121360:data<=-16'd13758;
      121361:data<=-16'd13026;
      121362:data<=-16'd13585;
      121363:data<=-16'd14771;
      121364:data<=-16'd13632;
      121365:data<=-16'd13123;
      121366:data<=-16'd13280;
      121367:data<=-16'd12013;
      121368:data<=-16'd11979;
      121369:data<=-16'd13658;
      121370:data<=-16'd14151;
      121371:data<=-16'd13059;
      121372:data<=-16'd12622;
      121373:data<=-16'd12659;
      121374:data<=-16'd11341;
      121375:data<=-16'd11100;
      121376:data<=-16'd12578;
      121377:data<=-16'd12671;
      121378:data<=-16'd11973;
      121379:data<=-16'd11101;
      121380:data<=-16'd10452;
      121381:data<=-16'd10910;
      121382:data<=-16'd10578;
      121383:data<=-16'd11429;
      121384:data<=-16'd11658;
      121385:data<=-16'd3953;
      121386:data<=16'd4093;
      121387:data<=16'd4585;
      121388:data<=16'd3921;
      121389:data<=16'd1945;
      121390:data<=-16'd2455;
      121391:data<=-16'd3287;
      121392:data<=-16'd2420;
      121393:data<=-16'd2532;
      121394:data<=-16'd1986;
      121395:data<=-16'd2734;
      121396:data<=-16'd4309;
      121397:data<=-16'd4394;
      121398:data<=-16'd4294;
      121399:data<=-16'd4317;
      121400:data<=-16'd3539;
      121401:data<=-16'd3040;
      121402:data<=-16'd4128;
      121403:data<=-16'd4980;
      121404:data<=-16'd4347;
      121405:data<=-16'd4830;
      121406:data<=-16'd5348;
      121407:data<=-16'd3800;
      121408:data<=-16'd3991;
      121409:data<=-16'd6068;
      121410:data<=-16'd6114;
      121411:data<=-16'd4983;
      121412:data<=-16'd4864;
      121413:data<=-16'd5600;
      121414:data<=-16'd5533;
      121415:data<=-16'd4992;
      121416:data<=-16'd5935;
      121417:data<=-16'd6311;
      121418:data<=-16'd5802;
      121419:data<=-16'd6499;
      121420:data<=-16'd6090;
      121421:data<=-16'd5647;
      121422:data<=-16'd7042;
      121423:data<=-16'd7291;
      121424:data<=-16'd7871;
      121425:data<=-16'd8372;
      121426:data<=-16'd7304;
      121427:data<=-16'd12323;
      121428:data<=-16'd21244;
      121429:data<=-16'd23141;
      121430:data<=-16'd21406;
      121431:data<=-16'd21197;
      121432:data<=-16'd20016;
      121433:data<=-16'd18600;
      121434:data<=-16'd17907;
      121435:data<=-16'd16736;
      121436:data<=-16'd15320;
      121437:data<=-16'd14942;
      121438:data<=-16'd15514;
      121439:data<=-16'd13602;
      121440:data<=-16'd9641;
      121441:data<=-16'd7928;
      121442:data<=-16'd6866;
      121443:data<=-16'd5100;
      121444:data<=-16'd4901;
      121445:data<=-16'd4936;
      121446:data<=-16'd4426;
      121447:data<=-16'd4534;
      121448:data<=-16'd3753;
      121449:data<=-16'd1572;
      121450:data<=-16'd183;
      121451:data<=-16'd120;
      121452:data<=16'd227;
      121453:data<=16'd97;
      121454:data<=-16'd869;
      121455:data<=16'd905;
      121456:data<=16'd3324;
      121457:data<=16'd2250;
      121458:data<=16'd2097;
      121459:data<=16'd3474;
      121460:data<=16'd2766;
      121461:data<=16'd2972;
      121462:data<=16'd4845;
      121463:data<=16'd6040;
      121464:data<=16'd6159;
      121465:data<=16'd5379;
      121466:data<=16'd6252;
      121467:data<=16'd6264;
      121468:data<=16'd4849;
      121469:data<=16'd12137;
      121470:data<=16'd22621;
      121471:data<=16'd22833;
      121472:data<=16'd20550;
      121473:data<=16'd20985;
      121474:data<=16'd19364;
      121475:data<=16'd19669;
      121476:data<=16'd21231;
      121477:data<=16'd19667;
      121478:data<=16'd18760;
      121479:data<=16'd18868;
      121480:data<=16'd17854;
      121481:data<=16'd17455;
      121482:data<=16'd17996;
      121483:data<=16'd18186;
      121484:data<=16'd17317;
      121485:data<=16'd16483;
      121486:data<=16'd15923;
      121487:data<=16'd14974;
      121488:data<=16'd15808;
      121489:data<=16'd16280;
      121490:data<=16'd13176;
      121491:data<=16'd11148;
      121492:data<=16'd10988;
      121493:data<=16'd9705;
      121494:data<=16'd9583;
      121495:data<=16'd10825;
      121496:data<=16'd11558;
      121497:data<=16'd11389;
      121498:data<=16'd10481;
      121499:data<=16'd10243;
      121500:data<=16'd9359;
      121501:data<=16'd8329;
      121502:data<=16'd9847;
      121503:data<=16'd10208;
      121504:data<=16'd8881;
      121505:data<=16'd8846;
      121506:data<=16'd8076;
      121507:data<=16'd7548;
      121508:data<=16'd7730;
      121509:data<=16'd7970;
      121510:data<=16'd9794;
      121511:data<=16'd5451;
      121512:data<=-16'd5286;
      121513:data<=-16'd8467;
      121514:data<=-16'd6147;
      121515:data<=-16'd5865;
      121516:data<=-16'd4504;
      121517:data<=-16'd3820;
      121518:data<=-16'd4458;
      121519:data<=-16'd3554;
      121520:data<=-16'd3392;
      121521:data<=-16'd3324;
      121522:data<=-16'd2120;
      121523:data<=-16'd1580;
      121524:data<=-16'd1444;
      121525:data<=-16'd1729;
      121526:data<=-16'd1886;
      121527:data<=-16'd1665;
      121528:data<=-16'd1647;
      121529:data<=-16'd432;
      121530:data<=16'd464;
      121531:data<=16'd83;
      121532:data<=16'd484;
      121533:data<=16'd447;
      121534:data<=16'd390;
      121535:data<=16'd1671;
      121536:data<=16'd2643;
      121537:data<=16'd2798;
      121538:data<=16'd1798;
      121539:data<=16'd2331;
      121540:data<=16'd5489;
      121541:data<=16'd5827;
      121542:data<=16'd5068;
      121543:data<=16'd5924;
      121544:data<=16'd4869;
      121545:data<=16'd4223;
      121546:data<=16'd4599;
      121547:data<=16'd4199;
      121548:data<=16'd4112;
      121549:data<=16'd2023;
      121550:data<=16'd1760;
      121551:data<=16'd3504;
      121552:data<=16'd414;
      121553:data<=16'd3962;
      121554:data<=16'd15534;
      121555:data<=16'd16578;
      121556:data<=16'd12786;
      121557:data<=16'd13458;
      121558:data<=16'd11735;
      121559:data<=16'd10602;
      121560:data<=16'd11333;
      121561:data<=16'd9303;
      121562:data<=16'd7228;
      121563:data<=16'd6229;
      121564:data<=16'd6396;
      121565:data<=16'd6849;
      121566:data<=16'd5788;
      121567:data<=16'd5841;
      121568:data<=16'd4946;
      121569:data<=16'd2413;
      121570:data<=16'd2748;
      121571:data<=16'd2902;
      121572:data<=16'd1817;
      121573:data<=16'd2215;
      121574:data<=16'd1741;
      121575:data<=16'd485;
      121576:data<=-16'd555;
      121577:data<=-16'd1096;
      121578:data<=-16'd281;
      121579:data<=-16'd220;
      121580:data<=-16'd252;
      121581:data<=-16'd655;
      121582:data<=-16'd2999;
      121583:data<=-16'd3218;
      121584:data<=-16'd2678;
      121585:data<=-16'd3694;
      121586:data<=-16'd3040;
      121587:data<=-16'd2975;
      121588:data<=-16'd3900;
      121589:data<=-16'd5090;
      121590:data<=-16'd8146;
      121591:data<=-16'd8505;
      121592:data<=-16'd8687;
      121593:data<=-16'd10537;
      121594:data<=-16'd7632;
      121595:data<=-16'd10308;
      121596:data<=-16'd21220;
      121597:data<=-16'd23033;
      121598:data<=-16'd19804;
      121599:data<=-16'd20477;
      121600:data<=-16'd19297;
      121601:data<=-16'd18953;
      121602:data<=-16'd20683;
      121603:data<=-16'd19826;
      121604:data<=-16'd18487;
      121605:data<=-16'd17685;
      121606:data<=-16'd17333;
      121607:data<=-16'd17384;
      121608:data<=-16'd16675;
      121609:data<=-16'd16918;
      121610:data<=-16'd16822;
      121611:data<=-16'd15603;
      121612:data<=-16'd15380;
      121613:data<=-16'd14104;
      121614:data<=-16'd13295;
      121615:data<=-16'd15236;
      121616:data<=-16'd15606;
      121617:data<=-16'd14302;
      121618:data<=-16'd13835;
      121619:data<=-16'd13292;
      121620:data<=-16'd12548;
      121621:data<=-16'd12334;
      121622:data<=-16'd13139;
      121623:data<=-16'd13235;
      121624:data<=-16'd12061;
      121625:data<=-16'd12145;
      121626:data<=-16'd11582;
      121627:data<=-16'd10226;
      121628:data<=-16'd11191;
      121629:data<=-16'd11611;
      121630:data<=-16'd10818;
      121631:data<=-16'd10417;
      121632:data<=-16'd9505;
      121633:data<=-16'd9749;
      121634:data<=-16'd9283;
      121635:data<=-16'd8558;
      121636:data<=-16'd10910;
      121637:data<=-16'd6749;
      121638:data<=16'd3970;
      121639:data<=16'd6792;
      121640:data<=16'd5489;
      121641:data<=16'd6649;
      121642:data<=16'd5771;
      121643:data<=16'd5650;
      121644:data<=16'd6670;
      121645:data<=16'd5292;
      121646:data<=16'd4830;
      121647:data<=16'd5072;
      121648:data<=16'd4884;
      121649:data<=16'd5665;
      121650:data<=16'd5203;
      121651:data<=16'd4649;
      121652:data<=16'd5485;
      121653:data<=16'd5175;
      121654:data<=16'd5436;
      121655:data<=16'd7294;
      121656:data<=16'd7908;
      121657:data<=16'd7656;
      121658:data<=16'd7691;
      121659:data<=16'd7248;
      121660:data<=16'd6537;
      121661:data<=16'd7104;
      121662:data<=16'd8575;
      121663:data<=16'd8604;
      121664:data<=16'd8372;
      121665:data<=16'd9292;
      121666:data<=16'd8853;
      121667:data<=16'd7700;
      121668:data<=16'd8343;
      121669:data<=16'd9356;
      121670:data<=16'd9213;
      121671:data<=16'd8793;
      121672:data<=16'd8953;
      121673:data<=16'd8311;
      121674:data<=16'd7600;
      121675:data<=16'd9492;
      121676:data<=16'd9762;
      121677:data<=16'd7868;
      121678:data<=16'd9538;
      121679:data<=16'd6777;
      121680:data<=-16'd3595;
      121681:data<=-16'd6196;
      121682:data<=-16'd1797;
      121683:data<=-16'd2115;
      121684:data<=-16'd3030;
      121685:data<=-16'd2035;
      121686:data<=-16'd2772;
      121687:data<=-16'd2504;
      121688:data<=-16'd332;
      121689:data<=16'd754;
      121690:data<=16'd58;
      121691:data<=-16'd1178;
      121692:data<=-16'd1856;
      121693:data<=-16'd2205;
      121694:data<=-16'd1155;
      121695:data<=16'd1014;
      121696:data<=16'd1095;
      121697:data<=16'd368;
      121698:data<=16'd925;
      121699:data<=16'd907;
      121700:data<=16'd790;
      121701:data<=16'd1874;
      121702:data<=16'd2901;
      121703:data<=16'd2983;
      121704:data<=16'd2855;
      121705:data<=16'd3193;
      121706:data<=16'd2770;
      121707:data<=16'd2296;
      121708:data<=16'd3645;
      121709:data<=16'd4552;
      121710:data<=16'd4396;
      121711:data<=16'd4742;
      121712:data<=16'd4711;
      121713:data<=16'd4683;
      121714:data<=16'd4840;
      121715:data<=16'd5310;
      121716:data<=16'd6445;
      121717:data<=16'd5970;
      121718:data<=16'd6213;
      121719:data<=16'd7178;
      121720:data<=16'd4778;
      121721:data<=16'd8395;
      121722:data<=16'd19317;
      121723:data<=16'd21735;
      121724:data<=16'd18704;
      121725:data<=16'd19053;
      121726:data<=16'd17719;
      121727:data<=16'd17009;
      121728:data<=16'd18842;
      121729:data<=16'd18031;
      121730:data<=16'd16738;
      121731:data<=16'd16365;
      121732:data<=16'd15327;
      121733:data<=16'd14712;
      121734:data<=16'd14509;
      121735:data<=16'd15103;
      121736:data<=16'd15286;
      121737:data<=16'd14220;
      121738:data<=16'd14172;
      121739:data<=16'd13509;
      121740:data<=16'd12745;
      121741:data<=16'd14906;
      121742:data<=16'd16131;
      121743:data<=16'd14954;
      121744:data<=16'd14176;
      121745:data<=16'd13444;
      121746:data<=16'd12839;
      121747:data<=16'd12777;
      121748:data<=16'd13259;
      121749:data<=16'd13667;
      121750:data<=16'd12437;
      121751:data<=16'd11367;
      121752:data<=16'd11280;
      121753:data<=16'd10686;
      121754:data<=16'd10058;
      121755:data<=16'd8966;
      121756:data<=16'd8337;
      121757:data<=16'd8379;
      121758:data<=16'd6965;
      121759:data<=16'd6616;
      121760:data<=16'd6129;
      121761:data<=16'd3491;
      121762:data<=16'd3718;
      121763:data<=16'd878;
      121764:data<=-16'd9142;
      121765:data<=-16'd12859;
      121766:data<=-16'd10090;
      121767:data<=-16'd11142;
      121768:data<=-16'd12871;
      121769:data<=-16'd12754;
      121770:data<=-16'd12965;
      121771:data<=-16'd12427;
      121772:data<=-16'd11244;
      121773:data<=-16'd10745;
      121774:data<=-16'd11761;
      121775:data<=-16'd12818;
      121776:data<=-16'd12507;
      121777:data<=-16'd12721;
      121778:data<=-16'd12420;
      121779:data<=-16'd11030;
      121780:data<=-16'd11500;
      121781:data<=-16'd12692;
      121782:data<=-16'd12982;
      121783:data<=-16'd12748;
      121784:data<=-16'd11960;
      121785:data<=-16'd11743;
      121786:data<=-16'd11629;
      121787:data<=-16'd11994;
      121788:data<=-16'd13443;
      121789:data<=-16'd12957;
      121790:data<=-16'd12383;
      121791:data<=-16'd13998;
      121792:data<=-16'd14154;
      121793:data<=-16'd13564;
      121794:data<=-16'd14105;
      121795:data<=-16'd14395;
      121796:data<=-16'd14058;
      121797:data<=-16'd12854;
      121798:data<=-16'd12725;
      121799:data<=-16'd13032;
      121800:data<=-16'd11761;
      121801:data<=-16'd12860;
      121802:data<=-16'd13468;
      121803:data<=-16'd11292;
      121804:data<=-16'd13042;
      121805:data<=-16'd10677;
      121806:data<=16'd273;
      121807:data<=16'd3221;
      121808:data<=-16'd1081;
      121809:data<=-16'd506;
      121810:data<=16'd358;
      121811:data<=-16'd698;
      121812:data<=16'd74;
      121813:data<=16'd212;
      121814:data<=-16'd1528;
      121815:data<=-16'd2783;
      121816:data<=-16'd2388;
      121817:data<=-16'd2302;
      121818:data<=-16'd3010;
      121819:data<=-16'd2073;
      121820:data<=-16'd2059;
      121821:data<=-16'd4390;
      121822:data<=-16'd4731;
      121823:data<=-16'd3932;
      121824:data<=-16'd4173;
      121825:data<=-16'd3706;
      121826:data<=-16'd3256;
      121827:data<=-16'd4109;
      121828:data<=-16'd5351;
      121829:data<=-16'd5526;
      121830:data<=-16'd4672;
      121831:data<=-16'd4619;
      121832:data<=-16'd4684;
      121833:data<=-16'd4434;
      121834:data<=-16'd5495;
      121835:data<=-16'd6405;
      121836:data<=-16'd6115;
      121837:data<=-16'd5486;
      121838:data<=-16'd4974;
      121839:data<=-16'd5441;
      121840:data<=-16'd5257;
      121841:data<=-16'd4485;
      121842:data<=-16'd5134;
      121843:data<=-16'd4657;
      121844:data<=-16'd4314;
      121845:data<=-16'd5435;
      121846:data<=-16'd4043;
      121847:data<=-16'd6792;
      121848:data<=-16'd16645;
      121849:data<=-16'd20196;
      121850:data<=-16'd17258;
      121851:data<=-16'd17283;
      121852:data<=-16'd17441;
      121853:data<=-16'd16463;
      121854:data<=-16'd17200;
      121855:data<=-16'd17270;
      121856:data<=-16'd15884;
      121857:data<=-16'd14750;
      121858:data<=-16'd14192;
      121859:data<=-16'd13809;
      121860:data<=-16'd13317;
      121861:data<=-16'd13106;
      121862:data<=-16'd12492;
      121863:data<=-16'd11185;
      121864:data<=-16'd10325;
      121865:data<=-16'd9926;
      121866:data<=-16'd9705;
      121867:data<=-16'd8457;
      121868:data<=-16'd6178;
      121869:data<=-16'd5653;
      121870:data<=-16'd5739;
      121871:data<=-16'd5031;
      121872:data<=-16'd5360;
      121873:data<=-16'd4687;
      121874:data<=-16'd2485;
      121875:data<=-16'd1773;
      121876:data<=-16'd1580;
      121877:data<=-16'd1025;
      121878:data<=-16'd954;
      121879:data<=-16'd1140;
      121880:data<=-16'd673;
      121881:data<=16'd1425;
      121882:data<=16'd2470;
      121883:data<=16'd1785;
      121884:data<=16'd2399;
      121885:data<=16'd2050;
      121886:data<=16'd1720;
      121887:data<=16'd3947;
      121888:data<=16'd3921;
      121889:data<=16'd6028;
      121890:data<=16'd14211;
      121891:data<=16'd17191;
      121892:data<=16'd14715;
      121893:data<=16'd15167;
      121894:data<=16'd15969;
      121895:data<=16'd15876;
      121896:data<=16'd16184;
      121897:data<=16'd15696;
      121898:data<=16'd15097;
      121899:data<=16'd14073;
      121900:data<=16'd13753;
      121901:data<=16'd14980;
      121902:data<=16'd14821;
      121903:data<=16'd14199;
      121904:data<=16'd14025;
      121905:data<=16'd12888;
      121906:data<=16'd12715;
      121907:data<=16'd13461;
      121908:data<=16'd13731;
      121909:data<=16'd13696;
      121910:data<=16'd12880;
      121911:data<=16'd12615;
      121912:data<=16'd12587;
      121913:data<=16'd11952;
      121914:data<=16'd13110;
      121915:data<=16'd14041;
      121916:data<=16'd12809;
      121917:data<=16'd12355;
      121918:data<=16'd11882;
      121919:data<=16'd10587;
      121920:data<=16'd10762;
      121921:data<=16'd11990;
      121922:data<=16'd12217;
      121923:data<=16'd10880;
      121924:data<=16'd10364;
      121925:data<=16'd10968;
      121926:data<=16'd10219;
      121927:data<=16'd10433;
      121928:data<=16'd11248;
      121929:data<=16'd9888;
      121930:data<=16'd9978;
      121931:data<=16'd8128;
      121932:data<=-16'd276;
      121933:data<=-16'd4993;
      121934:data<=-16'd2523;
      121935:data<=-16'd1689;
      121936:data<=-16'd2799;
      121937:data<=-16'd2464;
      121938:data<=-16'd2240;
      121939:data<=-16'd2340;
      121940:data<=-16'd1039;
      121941:data<=16'd1219;
      121942:data<=16'd2205;
      121943:data<=16'd1942;
      121944:data<=16'd1955;
      121945:data<=16'd1994;
      121946:data<=16'd1968;
      121947:data<=16'd2417;
      121948:data<=16'd3074;
      121949:data<=16'd3294;
      121950:data<=16'd3072;
      121951:data<=16'd3149;
      121952:data<=16'd2825;
      121953:data<=16'd2566;
      121954:data<=16'd4300;
      121955:data<=16'd5022;
      121956:data<=16'd3432;
      121957:data<=16'd3491;
      121958:data<=16'd4058;
      121959:data<=16'd3601;
      121960:data<=16'd4485;
      121961:data<=16'd5159;
      121962:data<=16'd4438;
      121963:data<=16'd4187;
      121964:data<=16'd4353;
      121965:data<=16'd4385;
      121966:data<=16'd3802;
      121967:data<=16'd3110;
      121968:data<=16'd3128;
      121969:data<=16'd2491;
      121970:data<=16'd2179;
      121971:data<=16'd2857;
      121972:data<=16'd2155;
      121973:data<=16'd3422;
      121974:data<=16'd9201;
      121975:data<=16'd12836;
      121976:data<=16'd12000;
      121977:data<=16'd11405;
      121978:data<=16'd11562;
      121979:data<=16'd10847;
      121980:data<=16'd9424;
      121981:data<=16'd7412;
      121982:data<=16'd6176;
      121983:data<=16'd6385;
      121984:data<=16'd6123;
      121985:data<=16'd5506;
      121986:data<=16'd5081;
      121987:data<=16'd3115;
      121988:data<=16'd1286;
      121989:data<=16'd1627;
      121990:data<=16'd1354;
      121991:data<=16'd238;
      121992:data<=16'd62;
      121993:data<=-16'd958;
      121994:data<=-16'd2757;
      121995:data<=-16'd3245;
      121996:data<=-16'd3018;
      121997:data<=-16'd2886;
      121998:data<=-16'd2786;
      121999:data<=-16'd2946;
      122000:data<=-16'd3782;
      122001:data<=-16'd5148;
      122002:data<=-16'd5435;
      122003:data<=-16'd4804;
      122004:data<=-16'd5169;
      122005:data<=-16'd5436;
      122006:data<=-16'd5147;
      122007:data<=-16'd6211;
      122008:data<=-16'd7122;
      122009:data<=-16'd6657;
      122010:data<=-16'd6790;
      122011:data<=-16'd6476;
      122012:data<=-16'd5375;
      122013:data<=-16'd6488;
      122014:data<=-16'd8114;
      122015:data<=-16'd9567;
      122016:data<=-16'd15220;
      122017:data<=-16'd21055;
      122018:data<=-16'd20729;
      122019:data<=-16'd19284;
      122020:data<=-16'd20477;
      122021:data<=-16'd20848;
      122022:data<=-16'd20011;
      122023:data<=-16'd19300;
      122024:data<=-16'd18360;
      122025:data<=-16'd17238;
      122026:data<=-16'd16683;
      122027:data<=-16'd17376;
      122028:data<=-16'd17708;
      122029:data<=-16'd16468;
      122030:data<=-16'd15666;
      122031:data<=-16'd15283;
      122032:data<=-16'd14184;
      122033:data<=-16'd14098;
      122034:data<=-16'd15082;
      122035:data<=-16'd14944;
      122036:data<=-16'd13861;
      122037:data<=-16'd13224;
      122038:data<=-16'd12756;
      122039:data<=-16'd12322;
      122040:data<=-16'd12615;
      122041:data<=-16'd12307;
      122042:data<=-16'd10712;
      122043:data<=-16'd9734;
      122044:data<=-16'd9072;
      122045:data<=-16'd8135;
      122046:data<=-16'd8439;
      122047:data<=-16'd9462;
      122048:data<=-16'd9691;
      122049:data<=-16'd8689;
      122050:data<=-16'd7536;
      122051:data<=-16'd7606;
      122052:data<=-16'd7363;
      122053:data<=-16'd7256;
      122054:data<=-16'd8419;
      122055:data<=-16'd7639;
      122056:data<=-16'd6596;
      122057:data<=-16'd6122;
      122058:data<=16'd229;
      122059:data<=16'd7473;
      122060:data<=16'd7162;
      122061:data<=16'd5547;
      122062:data<=16'd6237;
      122063:data<=16'd5729;
      122064:data<=16'd5375;
      122065:data<=16'd5655;
      122066:data<=16'd4692;
      122067:data<=16'd3284;
      122068:data<=16'd2984;
      122069:data<=16'd3659;
      122070:data<=16'd3495;
      122071:data<=16'd2646;
      122072:data<=16'd2670;
      122073:data<=16'd3051;
      122074:data<=16'd3403;
      122075:data<=16'd3469;
      122076:data<=16'd3303;
      122077:data<=16'd3668;
      122078:data<=16'd3436;
      122079:data<=16'd3465;
      122080:data<=16'd5368;
      122081:data<=16'd6296;
      122082:data<=16'd5785;
      122083:data<=16'd6015;
      122084:data<=16'd6096;
      122085:data<=16'd5741;
      122086:data<=16'd5937;
      122087:data<=16'd6804;
      122088:data<=16'd7445;
      122089:data<=16'd7048;
      122090:data<=16'd6980;
      122091:data<=16'd6375;
      122092:data<=16'd4361;
      122093:data<=16'd4948;
      122094:data<=16'd6986;
      122095:data<=16'd6652;
      122096:data<=16'd6445;
      122097:data<=16'd6516;
      122098:data<=16'd6141;
      122099:data<=16'd6114;
      122100:data<=16'd1897;
      122101:data<=-16'd4898;
      122102:data<=-16'd6275;
      122103:data<=-16'd4672;
      122104:data<=-16'd4845;
      122105:data<=-16'd4992;
      122106:data<=-16'd4250;
      122107:data<=-16'd2886;
      122108:data<=-16'd1583;
      122109:data<=-16'd1419;
      122110:data<=-16'd1268;
      122111:data<=-16'd870;
      122112:data<=-16'd694;
      122113:data<=16'd256;
      122114:data<=16'd1457;
      122115:data<=16'd1656;
      122116:data<=16'd1340;
      122117:data<=16'd1334;
      122118:data<=16'd1425;
      122119:data<=16'd1516;
      122120:data<=16'd2717;
      122121:data<=16'd4153;
      122122:data<=16'd3803;
      122123:data<=16'd3263;
      122124:data<=16'd3453;
      122125:data<=16'd3128;
      122126:data<=16'd3742;
      122127:data<=16'd5498;
      122128:data<=16'd6044;
      122129:data<=16'd5659;
      122130:data<=16'd5612;
      122131:data<=16'd5560;
      122132:data<=16'd5113;
      122133:data<=16'd5529;
      122134:data<=16'd7081;
      122135:data<=16'd7151;
      122136:data<=16'd6479;
      122137:data<=16'd6830;
      122138:data<=16'd6194;
      122139:data<=16'd6464;
      122140:data<=16'd8041;
      122141:data<=16'd8123;
      122142:data<=16'd13076;
      122143:data<=16'd22010;
      122144:data<=16'd22952;
      122145:data<=16'd20121;
      122146:data<=16'd21456;
      122147:data<=16'd21855;
      122148:data<=16'd20622;
      122149:data<=16'd20169;
      122150:data<=16'd19156;
      122151:data<=16'd18439;
      122152:data<=16'd17958;
      122153:data<=16'd17482;
      122154:data<=16'd17696;
      122155:data<=16'd17202;
      122156:data<=16'd16336;
      122157:data<=16'd15738;
      122158:data<=16'd15076;
      122159:data<=16'd15394;
      122160:data<=16'd16002;
      122161:data<=16'd15594;
      122162:data<=16'd14260;
      122163:data<=16'd13167;
      122164:data<=16'd13452;
      122165:data<=16'd13129;
      122166:data<=16'd12530;
      122167:data<=16'd13470;
      122168:data<=16'd12995;
      122169:data<=16'd11881;
      122170:data<=16'd12120;
      122171:data<=16'd10962;
      122172:data<=16'd10129;
      122173:data<=16'd10988;
      122174:data<=16'd11066;
      122175:data<=16'd10718;
      122176:data<=16'd9464;
      122177:data<=16'd8343;
      122178:data<=16'd8690;
      122179:data<=16'd7915;
      122180:data<=16'd7230;
      122181:data<=16'd6649;
      122182:data<=16'd5356;
      122183:data<=16'd6143;
      122184:data<=16'd2334;
      122185:data<=-16'd7441;
      122186:data<=-16'd10889;
      122187:data<=-16'd9937;
      122188:data<=-16'd11042;
      122189:data<=-16'd10605;
      122190:data<=-16'd10417;
      122191:data<=-16'd11524;
      122192:data<=-16'd11949;
      122193:data<=-16'd13417;
      122194:data<=-16'd13691;
      122195:data<=-16'd12753;
      122196:data<=-16'd13524;
      122197:data<=-16'd13279;
      122198:data<=-16'd12111;
      122199:data<=-16'd12610;
      122200:data<=-16'd13947;
      122201:data<=-16'd14832;
      122202:data<=-16'd14057;
      122203:data<=-16'd13112;
      122204:data<=-16'd13173;
      122205:data<=-16'd12797;
      122206:data<=-16'd13471;
      122207:data<=-16'd14631;
      122208:data<=-16'd13919;
      122209:data<=-16'd13361;
      122210:data<=-16'd13497;
      122211:data<=-16'd13176;
      122212:data<=-16'd12748;
      122213:data<=-16'd12927;
      122214:data<=-16'd14008;
      122215:data<=-16'd13756;
      122216:data<=-16'd12851;
      122217:data<=-16'd13147;
      122218:data<=-16'd11841;
      122219:data<=-16'd11176;
      122220:data<=-16'd12837;
      122221:data<=-16'd12443;
      122222:data<=-16'd11879;
      122223:data<=-16'd11426;
      122224:data<=-16'd10034;
      122225:data<=-16'd11351;
      122226:data<=-16'd8160;
      122227:data<=16'd1001;
      122228:data<=16'd2996;
      122229:data<=16'd917;
      122230:data<=16'd2080;
      122231:data<=16'd1859;
      122232:data<=16'd1143;
      122233:data<=16'd431;
      122234:data<=-16'd1688;
      122235:data<=-16'd1451;
      122236:data<=-16'd731;
      122237:data<=-16'd1198;
      122238:data<=-16'd520;
      122239:data<=-16'd1283;
      122240:data<=-16'd3148;
      122241:data<=-16'd2467;
      122242:data<=-16'd534;
      122243:data<=16'd126;
      122244:data<=-16'd538;
      122245:data<=-16'd834;
      122246:data<=-16'd1115;
      122247:data<=-16'd2296;
      122248:data<=-16'd2472;
      122249:data<=-16'd2311;
      122250:data<=-16'd2613;
      122251:data<=-16'd2065;
      122252:data<=-16'd2604;
      122253:data<=-16'd4087;
      122254:data<=-16'd4217;
      122255:data<=-16'd3651;
      122256:data<=-16'd2969;
      122257:data<=-16'd3254;
      122258:data<=-16'd3850;
      122259:data<=-16'd3683;
      122260:data<=-16'd5007;
      122261:data<=-16'd5557;
      122262:data<=-16'd4447;
      122263:data<=-16'd5209;
      122264:data<=-16'd5221;
      122265:data<=-16'd5338;
      122266:data<=-16'd6924;
      122267:data<=-16'd5604;
      122268:data<=-16'd8710;
      122269:data<=-16'd18077;
      122270:data<=-16'd20295;
      122271:data<=-16'd17832;
      122272:data<=-16'd18460;
      122273:data<=-16'd18554;
      122274:data<=-16'd18240;
      122275:data<=-16'd17693;
      122276:data<=-16'd16380;
      122277:data<=-16'd16486;
      122278:data<=-16'd15784;
      122279:data<=-16'd15177;
      122280:data<=-16'd16128;
      122281:data<=-16'd15250;
      122282:data<=-16'd14545;
      122283:data<=-16'd14818;
      122284:data<=-16'd13694;
      122285:data<=-16'd13217;
      122286:data<=-16'd12704;
      122287:data<=-16'd11656;
      122288:data<=-16'd11752;
      122289:data<=-16'd10702;
      122290:data<=-16'd9401;
      122291:data<=-16'd9982;
      122292:data<=-16'd10043;
      122293:data<=-16'd9024;
      122294:data<=-16'd7978;
      122295:data<=-16'd7395;
      122296:data<=-16'd7039;
      122297:data<=-16'd6485;
      122298:data<=-16'd6448;
      122299:data<=-16'd5077;
      122300:data<=-16'd2734;
      122301:data<=-16'd2707;
      122302:data<=-16'd2361;
      122303:data<=-16'd1084;
      122304:data<=-16'd1134;
      122305:data<=-16'd349;
      122306:data<=16'd789;
      122307:data<=16'd2052;
      122308:data<=16'd3104;
      122309:data<=16'd1606;
      122310:data<=16'd4989;
      122311:data<=16'd13938;
      122312:data<=16'd16728;
      122313:data<=16'd16333;
      122314:data<=16'd17687;
      122315:data<=16'd16192;
      122316:data<=16'd15109;
      122317:data<=16'd15465;
      122318:data<=16'd14142;
      122319:data<=16'd14634;
      122320:data<=16'd15963;
      122321:data<=16'd15444;
      122322:data<=16'd15050;
      122323:data<=16'd14333;
      122324:data<=16'd13562;
      122325:data<=16'd13978;
      122326:data<=16'd14904;
      122327:data<=16'd15593;
      122328:data<=16'd14862;
      122329:data<=16'd13896;
      122330:data<=16'd13493;
      122331:data<=16'd12302;
      122332:data<=16'd12436;
      122333:data<=16'd13825;
      122334:data<=16'd13577;
      122335:data<=16'd12885;
      122336:data<=16'd12486;
      122337:data<=16'd11996;
      122338:data<=16'd12044;
      122339:data<=16'd12477;
      122340:data<=16'd13080;
      122341:data<=16'd12954;
      122342:data<=16'd12986;
      122343:data<=16'd13740;
      122344:data<=16'd12631;
      122345:data<=16'd12090;
      122346:data<=16'd13396;
      122347:data<=16'd12756;
      122348:data<=16'd12111;
      122349:data<=16'd11432;
      122350:data<=16'd9897;
      122351:data<=16'd11188;
      122352:data<=16'd8537;
      122353:data<=-16'd140;
      122354:data<=-16'd3148;
      122355:data<=-16'd1930;
      122356:data<=-16'd2303;
      122357:data<=-16'd1613;
      122358:data<=-16'd1404;
      122359:data<=-16'd1228;
      122360:data<=16'd224;
      122361:data<=16'd109;
      122362:data<=16'd346;
      122363:data<=16'd698;
      122364:data<=-16'd420;
      122365:data<=16'd475;
      122366:data<=16'd1754;
      122367:data<=16'd1248;
      122368:data<=16'd1074;
      122369:data<=16'd1002;
      122370:data<=16'd1322;
      122371:data<=16'd1594;
      122372:data<=16'd1340;
      122373:data<=16'd2523;
      122374:data<=16'd3219;
      122375:data<=16'd2684;
      122376:data<=16'd2921;
      122377:data<=16'd2473;
      122378:data<=16'd2303;
      122379:data<=16'd3706;
      122380:data<=16'd4316;
      122381:data<=16'd3933;
      122382:data<=16'd3441;
      122383:data<=16'd3324;
      122384:data<=16'd3124;
      122385:data<=16'd2820;
      122386:data<=16'd4366;
      122387:data<=16'd4987;
      122388:data<=16'd3798;
      122389:data<=16'd4463;
      122390:data<=16'd4331;
      122391:data<=16'd3706;
      122392:data<=16'd3472;
      122393:data<=16'd140;
      122394:data<=16'd3092;
      122395:data<=16'd13397;
      122396:data<=16'd15255;
      122397:data<=16'd12504;
      122398:data<=16'd13032;
      122399:data<=16'd11142;
      122400:data<=16'd9784;
      122401:data<=16'd10131;
      122402:data<=16'd8214;
      122403:data<=16'd7711;
      122404:data<=16'd7794;
      122405:data<=16'd6322;
      122406:data<=16'd5275;
      122407:data<=16'd3723;
      122408:data<=16'd3266;
      122409:data<=16'd4100;
      122410:data<=16'd3656;
      122411:data<=16'd3345;
      122412:data<=16'd2147;
      122413:data<=16'd293;
      122414:data<=16'd557;
      122415:data<=16'd214;
      122416:data<=-16'd761;
      122417:data<=-16'd277;
      122418:data<=-16'd676;
      122419:data<=-16'd1886;
      122420:data<=-16'd2590;
      122421:data<=-16'd3031;
      122422:data<=-16'd3069;
      122423:data<=-16'd2878;
      122424:data<=-16'd2541;
      122425:data<=-16'd3472;
      122426:data<=-16'd5137;
      122427:data<=-16'd4905;
      122428:data<=-16'd4543;
      122429:data<=-16'd4742;
      122430:data<=-16'd4551;
      122431:data<=-16'd5109;
      122432:data<=-16'd5335;
      122433:data<=-16'd6334;
      122434:data<=-16'd7412;
      122435:data<=-16'd5448;
      122436:data<=-16'd8332;
      122437:data<=-16'd17026;
      122438:data<=-16'd19822;
      122439:data<=-16'd19079;
      122440:data<=-16'd20074;
      122441:data<=-16'd19112;
      122442:data<=-16'd17388;
      122443:data<=-16'd15782;
      122444:data<=-16'd14452;
      122445:data<=-16'd15662;
      122446:data<=-16'd16154;
      122447:data<=-16'd15006;
      122448:data<=-16'd14665;
      122449:data<=-16'd14208;
      122450:data<=-16'd14031;
      122451:data<=-16'd14099;
      122452:data<=-16'd13896;
      122453:data<=-16'd14073;
      122454:data<=-16'd13426;
      122455:data<=-16'd13039;
      122456:data<=-16'd13274;
      122457:data<=-16'd12010;
      122458:data<=-16'd11597;
      122459:data<=-16'd12443;
      122460:data<=-16'd11985;
      122461:data<=-16'd11400;
      122462:data<=-16'd11115;
      122463:data<=-16'd10508;
      122464:data<=-16'd9941;
      122465:data<=-16'd10037;
      122466:data<=-16'd10907;
      122467:data<=-16'd10131;
      122468:data<=-16'd9101;
      122469:data<=-16'd10064;
      122470:data<=-16'd9318;
      122471:data<=-16'd8275;
      122472:data<=-16'd9135;
      122473:data<=-16'd8708;
      122474:data<=-16'd8752;
      122475:data<=-16'd8490;
      122476:data<=-16'd6740;
      122477:data<=-16'd7853;
      122478:data<=-16'd5310;
      122479:data<=16'd3262;
      122480:data<=16'd6175;
      122481:data<=16'd5084;
      122482:data<=16'd5762;
      122483:data<=16'd5019;
      122484:data<=16'd4796;
      122485:data<=16'd5040;
      122486:data<=16'd3498;
      122487:data<=16'd3277;
      122488:data<=16'd3177;
      122489:data<=16'd2464;
      122490:data<=16'd3303;
      122491:data<=16'd3018;
      122492:data<=16'd1172;
      122493:data<=-16'd140;
      122494:data<=-16'd807;
      122495:data<=-16'd388;
      122496:data<=-16'd105;
      122497:data<=-16'd382;
      122498:data<=-16'd103;
      122499:data<=-16'd53;
      122500:data<=16'd112;
      122501:data<=16'd531;
      122502:data<=16'd472;
      122503:data<=16'd587;
      122504:data<=16'd560;
      122505:data<=16'd1284;
      122506:data<=16'd3051;
      122507:data<=16'd3156;
      122508:data<=16'd2740;
      122509:data<=16'd3339;
      122510:data<=16'd3397;
      122511:data<=16'd3744;
      122512:data<=16'd4772;
      122513:data<=16'd5430;
      122514:data<=16'd5482;
      122515:data<=16'd5131;
      122516:data<=16'd5541;
      122517:data<=16'd5154;
      122518:data<=16'd4639;
      122519:data<=16'd7310;
      122520:data<=16'd5604;
      122521:data<=-16'd3427;
      122522:data<=-16'd7329;
      122523:data<=-16'd5526;
      122524:data<=-16'd5606;
      122525:data<=-16'd4499;
      122526:data<=-16'd2264;
      122527:data<=-16'd2387;
      122528:data<=-16'd2373;
      122529:data<=-16'd1712;
      122530:data<=-16'd1677;
      122531:data<=-16'd1240;
      122532:data<=16'd118;
      122533:data<=16'd1463;
      122534:data<=16'd1275;
      122535:data<=16'd666;
      122536:data<=16'd1154;
      122537:data<=16'd1201;
      122538:data<=16'd1671;
      122539:data<=16'd3733;
      122540:data<=16'd4347;
      122541:data<=16'd3521;
      122542:data<=16'd4317;
      122543:data<=16'd5574;
      122544:data<=16'd5588;
      122545:data<=16'd6372;
      122546:data<=16'd7941;
      122547:data<=16'd7914;
      122548:data<=16'd7580;
      122549:data<=16'd7806;
      122550:data<=16'd7163;
      122551:data<=16'd7494;
      122552:data<=16'd8824;
      122553:data<=16'd8843;
      122554:data<=16'd8830;
      122555:data<=16'd8584;
      122556:data<=16'd7935;
      122557:data<=16'd8502;
      122558:data<=16'd8605;
      122559:data<=16'd9119;
      122560:data<=16'd10028;
      122561:data<=16'd8431;
      122562:data<=16'd11071;
      122563:data<=16'd19382;
      122564:data<=16'd22501;
      122565:data<=16'd21510;
      122566:data<=16'd21875;
      122567:data<=16'd20988;
      122568:data<=16'd20225;
      122569:data<=16'd20222;
      122570:data<=16'd18901;
      122571:data<=16'd18477;
      122572:data<=16'd18744;
      122573:data<=16'd18243;
      122574:data<=16'd17625;
      122575:data<=16'd16656;
      122576:data<=16'd16117;
      122577:data<=16'd15708;
      122578:data<=16'd15123;
      122579:data<=16'd15667;
      122580:data<=16'd15324;
      122581:data<=16'd14129;
      122582:data<=16'd14082;
      122583:data<=16'd12969;
      122584:data<=16'd11853;
      122585:data<=16'd12857;
      122586:data<=16'd13100;
      122587:data<=16'd12281;
      122588:data<=16'd11561;
      122589:data<=16'd10225;
      122590:data<=16'd9502;
      122591:data<=16'd10113;
      122592:data<=16'd10258;
      122593:data<=16'd8702;
      122594:data<=16'd7241;
      122595:data<=16'd7301;
      122596:data<=16'd6781;
      122597:data<=16'd6188;
      122598:data<=16'd6942;
      122599:data<=16'd6901;
      122600:data<=16'd6848;
      122601:data<=16'd6796;
      122602:data<=16'd5206;
      122603:data<=16'd5236;
      122604:data<=16'd3515;
      122605:data<=-16'd4422;
      122606:data<=-16'd9602;
      122607:data<=-16'd8681;
      122608:data<=-16'd8678;
      122609:data<=-16'd9057;
      122610:data<=-16'd8049;
      122611:data<=-16'd8617;
      122612:data<=-16'd10428;
      122613:data<=-16'd10915;
      122614:data<=-16'd9859;
      122615:data<=-16'd9327;
      122616:data<=-16'd9480;
      122617:data<=-16'd8931;
      122618:data<=-16'd9617;
      122619:data<=-16'd11348;
      122620:data<=-16'd10978;
      122621:data<=-16'd10147;
      122622:data<=-16'd10107;
      122623:data<=-16'd9310;
      122624:data<=-16'd9559;
      122625:data<=-16'd11045;
      122626:data<=-16'd10894;
      122627:data<=-16'd10313;
      122628:data<=-16'd10783;
      122629:data<=-16'd10063;
      122630:data<=-16'd8795;
      122631:data<=-16'd9735;
      122632:data<=-16'd11153;
      122633:data<=-16'd10933;
      122634:data<=-16'd10305;
      122635:data<=-16'd9864;
      122636:data<=-16'd9680;
      122637:data<=-16'd9917;
      122638:data<=-16'd10131;
      122639:data<=-16'd10766;
      122640:data<=-16'd10992;
      122641:data<=-16'd10302;
      122642:data<=-16'd10102;
      122643:data<=-16'd8429;
      122644:data<=-16'd6416;
      122645:data<=-16'd8536;
      122646:data<=-16'd8015;
      122647:data<=-16'd127;
      122648:data<=16'd5068;
      122649:data<=16'd4552;
      122650:data<=16'd4322;
      122651:data<=16'd3576;
      122652:data<=16'd1650;
      122653:data<=16'd1280;
      122654:data<=16'd1536;
      122655:data<=16'd961;
      122656:data<=16'd473;
      122657:data<=16'd490;
      122658:data<=-16'd285;
      122659:data<=-16'd1735;
      122660:data<=-16'd1754;
      122661:data<=-16'd1409;
      122662:data<=-16'd1891;
      122663:data<=-16'd1371;
      122664:data<=-16'd1556;
      122665:data<=-16'd3636;
      122666:data<=-16'd4050;
      122667:data<=-16'd3529;
      122668:data<=-16'd4420;
      122669:data<=-16'd4407;
      122670:data<=-16'd3735;
      122671:data<=-16'd4875;
      122672:data<=-16'd6137;
      122673:data<=-16'd5879;
      122674:data<=-16'd5735;
      122675:data<=-16'd6181;
      122676:data<=-16'd5897;
      122677:data<=-16'd5570;
      122678:data<=-16'd6358;
      122679:data<=-16'd7142;
      122680:data<=-16'd7141;
      122681:data<=-16'd6728;
      122682:data<=-16'd6206;
      122683:data<=-16'd5970;
      122684:data<=-16'd6178;
      122685:data<=-16'd7633;
      122686:data<=-16'd8989;
      122687:data<=-16'd7247;
      122688:data<=-16'd7521;
      122689:data<=-16'd14543;
      122690:data<=-16'd19905;
      122691:data<=-16'd19456;
      122692:data<=-16'd19751;
      122693:data<=-16'd20936;
      122694:data<=-16'd20354;
      122695:data<=-16'd19776;
      122696:data<=-16'd19017;
      122697:data<=-16'd18271;
      122698:data<=-16'd18771;
      122699:data<=-16'd18616;
      122700:data<=-16'd17305;
      122701:data<=-16'd16421;
      122702:data<=-16'd15816;
      122703:data<=-16'd15223;
      122704:data<=-16'd15329;
      122705:data<=-16'd15982;
      122706:data<=-16'd15690;
      122707:data<=-16'd14509;
      122708:data<=-16'd14046;
      122709:data<=-16'd13465;
      122710:data<=-16'd12345;
      122711:data<=-16'd12091;
      122712:data<=-16'd11529;
      122713:data<=-16'd10366;
      122714:data<=-16'd10016;
      122715:data<=-16'd9219;
      122716:data<=-16'd8147;
      122717:data<=-16'd7861;
      122718:data<=-16'd6663;
      122719:data<=-16'd5319;
      122720:data<=-16'd5407;
      122721:data<=-16'd4830;
      122722:data<=-16'd3515;
      122723:data<=-16'd3653;
      122724:data<=-16'd3563;
      122725:data<=-16'd1281;
      122726:data<=16'd206;
      122727:data<=-16'd247;
      122728:data<=16'd284;
      122729:data<=16'd358;
      122730:data<=16'd702;
      122731:data<=16'd7774;
      122732:data<=16'd16186;
      122733:data<=16'd16475;
      122734:data<=16'd14507;
      122735:data<=16'd15311;
      122736:data<=16'd14800;
      122737:data<=16'd13905;
      122738:data<=16'd14775;
      122739:data<=16'd15186;
      122740:data<=16'd14525;
      122741:data<=16'd13920;
      122742:data<=16'd13665;
      122743:data<=16'd13541;
      122744:data<=16'd14302;
      122745:data<=16'd15861;
      122746:data<=16'd15758;
      122747:data<=16'd14690;
      122748:data<=16'd14818;
      122749:data<=16'd14586;
      122750:data<=16'd13684;
      122751:data<=16'd13396;
      122752:data<=16'd13558;
      122753:data<=16'd14075;
      122754:data<=16'd13926;
      122755:data<=16'd12844;
      122756:data<=16'd12075;
      122757:data<=16'd11712;
      122758:data<=16'd12239;
      122759:data<=16'd12980;
      122760:data<=16'd12534;
      122761:data<=16'd12240;
      122762:data<=16'd11849;
      122763:data<=16'd10796;
      122764:data<=16'd11212;
      122765:data<=16'd12260;
      122766:data<=16'd12125;
      122767:data<=16'd11605;
      122768:data<=16'd11203;
      122769:data<=16'd10558;
      122770:data<=16'd9471;
      122771:data<=16'd10023;
      122772:data<=16'd10807;
      122773:data<=16'd5124;
      122774:data<=-16'd2540;
      122775:data<=-16'd3272;
      122776:data<=-16'd2320;
      122777:data<=-16'd3052;
      122778:data<=-16'd1491;
      122779:data<=-16'd484;
      122780:data<=-16'd1216;
      122781:data<=-16'd760;
      122782:data<=-16'd746;
      122783:data<=-16'd1001;
      122784:data<=16'd469;
      122785:data<=16'd1698;
      122786:data<=16'd1471;
      122787:data<=16'd1233;
      122788:data<=16'd1475;
      122789:data<=16'd1154;
      122790:data<=16'd717;
      122791:data<=16'd1659;
      122792:data<=16'd2549;
      122793:data<=16'd1964;
      122794:data<=16'd1013;
      122795:data<=16'd127;
      122796:data<=-16'd331;
      122797:data<=16'd461;
      122798:data<=16'd1962;
      122799:data<=16'd2593;
      122800:data<=16'd1870;
      122801:data<=16'd1848;
      122802:data<=16'd2434;
      122803:data<=16'd1707;
      122804:data<=16'd2011;
      122805:data<=16'd3668;
      122806:data<=16'd3573;
      122807:data<=16'd2974;
      122808:data<=16'd2955;
      122809:data<=16'd2793;
      122810:data<=16'd3054;
      122811:data<=16'd3516;
      122812:data<=16'd4781;
      122813:data<=16'd5034;
      122814:data<=16'd3550;
      122815:data<=16'd8049;
      122816:data<=16'd16377;
      122817:data<=16'd17144;
      122818:data<=16'd14211;
      122819:data<=16'd14114;
      122820:data<=16'd13825;
      122821:data<=16'd13480;
      122822:data<=16'd13494;
      122823:data<=16'd12284;
      122824:data<=16'd10464;
      122825:data<=16'd8445;
      122826:data<=16'd8053;
      122827:data<=16'd8578;
      122828:data<=16'd7175;
      122829:data<=16'd6354;
      122830:data<=16'd6132;
      122831:data<=16'd4223;
      122832:data<=16'd3441;
      122833:data<=16'd3805;
      122834:data<=16'd3136;
      122835:data<=16'd2340;
      122836:data<=16'd1767;
      122837:data<=16'd1175;
      122838:data<=-16'd328;
      122839:data<=-16'd1700;
      122840:data<=-16'd610;
      122841:data<=-16'd309;
      122842:data<=-16'd1615;
      122843:data<=-16'd741;
      122844:data<=-16'd99;
      122845:data<=-16'd1342;
      122846:data<=-16'd1445;
      122847:data<=-16'd1113;
      122848:data<=-16'd1676;
      122849:data<=-16'd1971;
      122850:data<=-16'd2071;
      122851:data<=-16'd3410;
      122852:data<=-16'd4827;
      122853:data<=-16'd4123;
      122854:data<=-16'd4331;
      122855:data<=-16'd5203;
      122856:data<=-16'd3268;
      122857:data<=-16'd6904;
      122858:data<=-16'd17403;
      122859:data<=-16'd20172;
      122860:data<=-16'd16804;
      122861:data<=-16'd17211;
      122862:data<=-16'd17059;
      122863:data<=-16'd15414;
      122864:data<=-16'd16261;
      122865:data<=-16'd16907;
      122866:data<=-16'd16267;
      122867:data<=-16'd15775;
      122868:data<=-16'd15091;
      122869:data<=-16'd14187;
      122870:data<=-16'd13888;
      122871:data<=-16'd14953;
      122872:data<=-16'd15675;
      122873:data<=-16'd14769;
      122874:data<=-16'd13913;
      122875:data<=-16'd13159;
      122876:data<=-16'd12474;
      122877:data<=-16'd12895;
      122878:data<=-16'd13402;
      122879:data<=-16'd13162;
      122880:data<=-16'd12481;
      122881:data<=-16'd11972;
      122882:data<=-16'd11629;
      122883:data<=-16'd10898;
      122884:data<=-16'd11230;
      122885:data<=-16'd11931;
      122886:data<=-16'd11154;
      122887:data<=-16'd11006;
      122888:data<=-16'd10511;
      122889:data<=-16'd8812;
      122890:data<=-16'd9579;
      122891:data<=-16'd10859;
      122892:data<=-16'd10363;
      122893:data<=-16'd10423;
      122894:data<=-16'd10772;
      122895:data<=-16'd10959;
      122896:data<=-16'd10114;
      122897:data<=-16'd9800;
      122898:data<=-16'd12290;
      122899:data<=-16'd8387;
      122900:data<=16'd1970;
      122901:data<=16'd4350;
      122902:data<=16'd2457;
      122903:data<=16'd3738;
      122904:data<=16'd2314;
      122905:data<=16'd688;
      122906:data<=16'd1642;
      122907:data<=16'd1037;
      122908:data<=16'd901;
      122909:data<=16'd1330;
      122910:data<=16'd187;
      122911:data<=-16'd694;
      122912:data<=-16'd934;
      122913:data<=-16'd376;
      122914:data<=-16'd138;
      122915:data<=-16'd772;
      122916:data<=16'd115;
      122917:data<=16'd100;
      122918:data<=-16'd1818;
      122919:data<=-16'd2190;
      122920:data<=-16'd1980;
      122921:data<=-16'd1559;
      122922:data<=-16'd705;
      122923:data<=-16'd975;
      122924:data<=-16'd828;
      122925:data<=-16'd688;
      122926:data<=-16'd1236;
      122927:data<=-16'd497;
      122928:data<=-16'd36;
      122929:data<=-16'd182;
      122930:data<=16'd590;
      122931:data<=16'd1532;
      122932:data<=16'd2358;
      122933:data<=16'd2083;
      122934:data<=16'd1809;
      122935:data<=16'd2572;
      122936:data<=16'd2159;
      122937:data<=16'd3098;
      122938:data<=16'd4655;
      122939:data<=16'd3647;
      122940:data<=16'd4684;
      122941:data<=16'd2355;
      122942:data<=-16'd7136;
      122943:data<=-16'd8796;
      122944:data<=-16'd3586;
      122945:data<=-16'd3595;
      122946:data<=-16'd3568;
      122947:data<=-16'd1809;
      122948:data<=-16'd2469;
      122949:data<=-16'd2478;
      122950:data<=-16'd1563;
      122951:data<=-16'd325;
      122952:data<=16'd1027;
      122953:data<=16'd593;
      122954:data<=16'd701;
      122955:data<=16'd1513;
      122956:data<=16'd1248;
      122957:data<=16'd2161;
      122958:data<=16'd3557;
      122959:data<=16'd3597;
      122960:data<=16'd3870;
      122961:data<=16'd4689;
      122962:data<=16'd4593;
      122963:data<=16'd3896;
      122964:data<=16'd4877;
      122965:data<=16'd6360;
      122966:data<=16'd5844;
      122967:data<=16'd5670;
      122968:data<=16'd5971;
      122969:data<=16'd5198;
      122970:data<=16'd5630;
      122971:data<=16'd6804;
      122972:data<=16'd7316;
      122973:data<=16'd7636;
      122974:data<=16'd7379;
      122975:data<=16'd7413;
      122976:data<=16'd6984;
      122977:data<=16'd6702;
      122978:data<=16'd8572;
      122979:data<=16'd8522;
      122980:data<=16'd7732;
      122981:data<=16'd8425;
      122982:data<=16'd6028;
      122983:data<=16'd8957;
      122984:data<=16'd20145;
      122985:data<=16'd23175;
      122986:data<=16'd20019;
      122987:data<=16'd20597;
      122988:data<=16'd19399;
      122989:data<=16'd17823;
      122990:data<=16'd18888;
      122991:data<=16'd18534;
      122992:data<=16'd18133;
      122993:data<=16'd17297;
      122994:data<=16'd15068;
      122995:data<=16'd14213;
      122996:data<=16'd13581;
      122997:data<=16'd13376;
      122998:data<=16'd14022;
      122999:data<=16'd13456;
      123000:data<=16'd13207;
      123001:data<=16'd12859;
      123002:data<=16'd11427;
      123003:data<=16'd11506;
      123004:data<=16'd12252;
      123005:data<=16'd12038;
      123006:data<=16'd11485;
      123007:data<=16'd11138;
      123008:data<=16'd11082;
      123009:data<=16'd10047;
      123010:data<=16'd9691;
      123011:data<=16'd11039;
      123012:data<=16'd10651;
      123013:data<=16'd9814;
      123014:data<=16'd9896;
      123015:data<=16'd8596;
      123016:data<=16'd7958;
      123017:data<=16'd8718;
      123018:data<=16'd9197;
      123019:data<=16'd9182;
      123020:data<=16'd8022;
      123021:data<=16'd7444;
      123022:data<=16'd6910;
      123023:data<=16'd6367;
      123024:data<=16'd8775;
      123025:data<=16'd5702;
      123026:data<=-16'd4387;
      123027:data<=-16'd6849;
      123028:data<=-16'd4848;
      123029:data<=-16'd6887;
      123030:data<=-16'd6660;
      123031:data<=-16'd5695;
      123032:data<=-16'd6581;
      123033:data<=-16'd5442;
      123034:data<=-16'd5342;
      123035:data<=-16'd6132;
      123036:data<=-16'd5676;
      123037:data<=-16'd6846;
      123038:data<=-16'd7553;
      123039:data<=-16'd6922;
      123040:data<=-16'd7418;
      123041:data<=-16'd7453;
      123042:data<=-16'd7021;
      123043:data<=-16'd7033;
      123044:data<=-16'd6957;
      123045:data<=-16'd6977;
      123046:data<=-16'd6422;
      123047:data<=-16'd5923;
      123048:data<=-16'd5839;
      123049:data<=-16'd5586;
      123050:data<=-16'd6683;
      123051:data<=-16'd7952;
      123052:data<=-16'd7708;
      123053:data<=-16'd7517;
      123054:data<=-16'd7271;
      123055:data<=-16'd6790;
      123056:data<=-16'd6878;
      123057:data<=-16'd7682;
      123058:data<=-16'd8498;
      123059:data<=-16'd7747;
      123060:data<=-16'd7424;
      123061:data<=-16'd7790;
      123062:data<=-16'd6305;
      123063:data<=-16'd6916;
      123064:data<=-16'd8721;
      123065:data<=-16'd7961;
      123066:data<=-16'd9068;
      123067:data<=-16'd6495;
      123068:data<=16'd3222;
      123069:data<=16'd6354;
      123070:data<=16'd3419;
      123071:data<=16'd3298;
      123072:data<=16'd2552;
      123073:data<=16'd2021;
      123074:data<=16'd2977;
      123075:data<=16'd2481;
      123076:data<=16'd2256;
      123077:data<=16'd878;
      123078:data<=-16'd1356;
      123079:data<=-16'd820;
      123080:data<=-16'd538;
      123081:data<=-16'd884;
      123082:data<=-16'd391;
      123083:data<=-16'd1568;
      123084:data<=-16'd3083;
      123085:data<=-16'd3597;
      123086:data<=-16'd3814;
      123087:data<=-16'd3375;
      123088:data<=-16'd3260;
      123089:data<=-16'd3347;
      123090:data<=-16'd3991;
      123091:data<=-16'd5269;
      123092:data<=-16'd4842;
      123093:data<=-16'd4851;
      123094:data<=-16'd6364;
      123095:data<=-16'd6479;
      123096:data<=-16'd6975;
      123097:data<=-16'd8511;
      123098:data<=-16'd8804;
      123099:data<=-16'd8352;
      123100:data<=-16'd8028;
      123101:data<=-16'd8102;
      123102:data<=-16'd7580;
      123103:data<=-16'd7539;
      123104:data<=-16'd9439;
      123105:data<=-16'd9229;
      123106:data<=-16'd8490;
      123107:data<=-16'd9400;
      123108:data<=-16'd7169;
      123109:data<=-16'd9185;
      123110:data<=-16'd19035;
      123111:data<=-16'd22615;
      123112:data<=-16'd20583;
      123113:data<=-16'd21137;
      123114:data<=-16'd20259;
      123115:data<=-16'd18707;
      123116:data<=-16'd18964;
      123117:data<=-16'd19039;
      123118:data<=-16'd19296;
      123119:data<=-16'd18559;
      123120:data<=-16'd17397;
      123121:data<=-16'd16830;
      123122:data<=-16'd15130;
      123123:data<=-16'd15121;
      123124:data<=-16'd16574;
      123125:data<=-16'd15717;
      123126:data<=-16'd14750;
      123127:data<=-16'd14052;
      123128:data<=-16'd12659;
      123129:data<=-16'd12605;
      123130:data<=-16'd13285;
      123131:data<=-16'd13653;
      123132:data<=-16'd13207;
      123133:data<=-16'd11935;
      123134:data<=-16'd11304;
      123135:data<=-16'd10545;
      123136:data<=-16'd9882;
      123137:data<=-16'd9785;
      123138:data<=-16'd8724;
      123139:data<=-16'd8332;
      123140:data<=-16'd8329;
      123141:data<=-16'd7242;
      123142:data<=-16'd6953;
      123143:data<=-16'd5418;
      123144:data<=-16'd2605;
      123145:data<=-16'd1874;
      123146:data<=-16'd1086;
      123147:data<=-16'd133;
      123148:data<=16'd402;
      123149:data<=16'd1542;
      123150:data<=16'd1066;
      123151:data<=16'd4235;
      123152:data<=16'd13186;
      123153:data<=16'd16487;
      123154:data<=16'd14252;
      123155:data<=16'd14184;
      123156:data<=16'd14609;
      123157:data<=16'd15523;
      123158:data<=16'd16366;
      123159:data<=16'd14897;
      123160:data<=16'd14516;
      123161:data<=16'd14821;
      123162:data<=16'd13850;
      123163:data<=16'd14264;
      123164:data<=16'd15183;
      123165:data<=16'd14671;
      123166:data<=16'd13940;
      123167:data<=16'd13590;
      123168:data<=16'd13192;
      123169:data<=16'd12690;
      123170:data<=16'd13250;
      123171:data<=16'd14173;
      123172:data<=16'd13600;
      123173:data<=16'd13068;
      123174:data<=16'd12813;
      123175:data<=16'd11879;
      123176:data<=16'd12063;
      123177:data<=16'd12798;
      123178:data<=16'd12433;
      123179:data<=16'd11781;
      123180:data<=16'd11327;
      123181:data<=16'd10933;
      123182:data<=16'd10446;
      123183:data<=16'd10769;
      123184:data<=16'd11526;
      123185:data<=16'd10645;
      123186:data<=16'd10225;
      123187:data<=16'd10477;
      123188:data<=16'd8912;
      123189:data<=16'd8868;
      123190:data<=16'd9838;
      123191:data<=16'd9453;
      123192:data<=16'd10983;
      123193:data<=16'd8539;
      123194:data<=-16'd1375;
      123195:data<=-16'd6490;
      123196:data<=-16'd4570;
      123197:data<=-16'd3594;
      123198:data<=-16'd3609;
      123199:data<=-16'd3701;
      123200:data<=-16'd3791;
      123201:data<=-16'd3237;
      123202:data<=-16'd3313;
      123203:data<=-16'd2667;
      123204:data<=-16'd1158;
      123205:data<=-16'd908;
      123206:data<=-16'd769;
      123207:data<=-16'd560;
      123208:data<=-16'd913;
      123209:data<=-16'd508;
      123210:data<=16'd714;
      123211:data<=16'd1873;
      123212:data<=16'd1838;
      123213:data<=16'd1078;
      123214:data<=16'd1104;
      123215:data<=16'd647;
      123216:data<=16'd619;
      123217:data<=16'd2540;
      123218:data<=16'd3078;
      123219:data<=16'd2458;
      123220:data<=16'd3031;
      123221:data<=16'd2631;
      123222:data<=16'd1962;
      123223:data<=16'd3265;
      123224:data<=16'd4451;
      123225:data<=16'd4211;
      123226:data<=16'd3991;
      123227:data<=16'd4150;
      123228:data<=16'd3237;
      123229:data<=16'd2783;
      123230:data<=16'd4837;
      123231:data<=16'd5533;
      123232:data<=16'd4789;
      123233:data<=16'd5503;
      123234:data<=16'd3970;
      123235:data<=16'd4645;
      123236:data<=16'd13400;
      123237:data<=16'd18838;
      123238:data<=16'd16979;
      123239:data<=16'd16348;
      123240:data<=16'd15835;
      123241:data<=16'd14666;
      123242:data<=16'd14897;
      123243:data<=16'd13728;
      123244:data<=16'd13251;
      123245:data<=16'd14672;
      123246:data<=16'd14252;
      123247:data<=16'd13335;
      123248:data<=16'd12938;
      123249:data<=16'd11347;
      123250:data<=16'd9323;
      123251:data<=16'd8204;
      123252:data<=16'd8302;
      123253:data<=16'd7638;
      123254:data<=16'd6199;
      123255:data<=16'd6542;
      123256:data<=16'd6017;
      123257:data<=16'd3833;
      123258:data<=16'd3747;
      123259:data<=16'd3927;
      123260:data<=16'd2816;
      123261:data<=16'd2555;
      123262:data<=16'd2050;
      123263:data<=16'd388;
      123264:data<=-16'd778;
      123265:data<=-16'd864;
      123266:data<=-16'd875;
      123267:data<=-16'd1075;
      123268:data<=-16'd930;
      123269:data<=-16'd1850;
      123270:data<=-16'd3442;
      123271:data<=-16'd3500;
      123272:data<=-16'd3509;
      123273:data<=-16'd3751;
      123274:data<=-16'd3597;
      123275:data<=-16'd3959;
      123276:data<=-16'd3706;
      123277:data<=-16'd6589;
      123278:data<=-16'd14451;
      123279:data<=-16'd18298;
      123280:data<=-16'd17141;
      123281:data<=-16'd16804;
      123282:data<=-16'd16641;
      123283:data<=-16'd17471;
      123284:data<=-16'd18359;
      123285:data<=-16'd16873;
      123286:data<=-16'd16483;
      123287:data<=-16'd16480;
      123288:data<=-16'd15233;
      123289:data<=-16'd15678;
      123290:data<=-16'd16358;
      123291:data<=-16'd15916;
      123292:data<=-16'd15095;
      123293:data<=-16'd13809;
      123294:data<=-16'd13967;
      123295:data<=-16'd14722;
      123296:data<=-16'd15050;
      123297:data<=-16'd16263;
      123298:data<=-16'd16267;
      123299:data<=-16'd15634;
      123300:data<=-16'd15860;
      123301:data<=-16'd14556;
      123302:data<=-16'd13637;
      123303:data<=-16'd14483;
      123304:data<=-16'd14404;
      123305:data<=-16'd13858;
      123306:data<=-16'd13203;
      123307:data<=-16'd12079;
      123308:data<=-16'd11517;
      123309:data<=-16'd11729;
      123310:data<=-16'd12390;
      123311:data<=-16'd12134;
      123312:data<=-16'd11541;
      123313:data<=-16'd11627;
      123314:data<=-16'd10399;
      123315:data<=-16'd9797;
      123316:data<=-16'd10812;
      123317:data<=-16'd10756;
      123318:data<=-16'd11499;
      123319:data<=-16'd9592;
      123320:data<=-16'd1155;
      123321:data<=16'd4431;
      123322:data<=16'd3570;
      123323:data<=16'd2083;
      123324:data<=16'd1337;
      123325:data<=16'd2123;
      123326:data<=16'd2870;
      123327:data<=16'd2055;
      123328:data<=16'd2729;
      123329:data<=16'd2728;
      123330:data<=16'd795;
      123331:data<=16'd799;
      123332:data<=16'd1075;
      123333:data<=16'd540;
      123334:data<=16'd1101;
      123335:data<=16'd1007;
      123336:data<=-16'd284;
      123337:data<=-16'd1409;
      123338:data<=-16'd1795;
      123339:data<=-16'd1316;
      123340:data<=-16'd679;
      123341:data<=16'd325;
      123342:data<=16'd318;
      123343:data<=-16'd1768;
      123344:data<=-16'd2052;
      123345:data<=-16'd206;
      123346:data<=16'd397;
      123347:data<=16'd581;
      123348:data<=16'd707;
      123349:data<=16'd429;
      123350:data<=16'd1102;
      123351:data<=16'd1448;
      123352:data<=16'd657;
      123353:data<=16'd647;
      123354:data<=16'd1306;
      123355:data<=16'd1485;
      123356:data<=16'd2065;
      123357:data<=16'd3483;
      123358:data<=16'd3773;
      123359:data<=16'd3297;
      123360:data<=16'd4284;
      123361:data<=16'd2822;
      123362:data<=-16'd3488;
      123363:data<=-16'd7283;
      123364:data<=-16'd6090;
      123365:data<=-16'd5550;
      123366:data<=-16'd6024;
      123367:data<=-16'd5749;
      123368:data<=-16'd5623;
      123369:data<=-16'd4526;
      123370:data<=-16'd2541;
      123371:data<=-16'd2076;
      123372:data<=-16'd2458;
      123373:data<=-16'd2185;
      123374:data<=-16'd1945;
      123375:data<=-16'd1466;
      123376:data<=16'd390;
      123377:data<=16'd2164;
      123378:data<=16'd2170;
      123379:data<=16'd1953;
      123380:data<=16'd2088;
      123381:data<=16'd1592;
      123382:data<=16'd2319;
      123383:data<=16'd4209;
      123384:data<=16'd4328;
      123385:data<=16'd3894;
      123386:data<=16'd4464;
      123387:data<=16'd4531;
      123388:data<=16'd4384;
      123389:data<=16'd4984;
      123390:data<=16'd5867;
      123391:data<=16'd6169;
      123392:data<=16'd5873;
      123393:data<=16'd6178;
      123394:data<=16'd6070;
      123395:data<=16'd5053;
      123396:data<=16'd5483;
      123397:data<=16'd6138;
      123398:data<=16'd5647;
      123399:data<=16'd5439;
      123400:data<=16'd4939;
      123401:data<=16'd4977;
      123402:data<=16'd5999;
      123403:data<=16'd7705;
      123404:data<=16'd13605;
      123405:data<=16'd19973;
      123406:data<=16'd20118;
      123407:data<=16'd18434;
      123408:data<=16'd17996;
      123409:data<=16'd17761;
      123410:data<=16'd18942;
      123411:data<=16'd19055;
      123412:data<=16'd17707;
      123413:data<=16'd17285;
      123414:data<=16'd16537;
      123415:data<=16'd16606;
      123416:data<=16'd17547;
      123417:data<=16'd16757;
      123418:data<=16'd15737;
      123419:data<=16'd14973;
      123420:data<=16'd13947;
      123421:data<=16'd13662;
      123422:data<=16'd13761;
      123423:data<=16'd14480;
      123424:data<=16'd14590;
      123425:data<=16'd13485;
      123426:data<=16'd13377;
      123427:data<=16'd12590;
      123428:data<=16'd11285;
      123429:data<=16'd12275;
      123430:data<=16'd12848;
      123431:data<=16'd12225;
      123432:data<=16'd12002;
      123433:data<=16'd11223;
      123434:data<=16'd10519;
      123435:data<=16'd10378;
      123436:data<=16'd11001;
      123437:data<=16'd11515;
      123438:data<=16'd9990;
      123439:data<=16'd9215;
      123440:data<=16'd9163;
      123441:data<=16'd7993;
      123442:data<=16'd8869;
      123443:data<=16'd9280;
      123444:data<=16'd8445;
      123445:data<=16'd9427;
      123446:data<=16'd4696;
      123447:data<=-16'd4093;
      123448:data<=-16'd5013;
      123449:data<=-16'd2446;
      123450:data<=-16'd2481;
      123451:data<=-16'd2437;
      123452:data<=-16'd2914;
      123453:data<=-16'd3319;
      123454:data<=-16'd2529;
      123455:data<=-16'd2102;
      123456:data<=-16'd2428;
      123457:data<=-16'd3436;
      123458:data<=-16'd3227;
      123459:data<=-16'd2082;
      123460:data<=-16'd2520;
      123461:data<=-16'd2669;
      123462:data<=-16'd3080;
      123463:data<=-16'd5212;
      123464:data<=-16'd5668;
      123465:data<=-16'd4986;
      123466:data<=-16'd4962;
      123467:data<=-16'd4526;
      123468:data<=-16'd4937;
      123469:data<=-16'd6244;
      123470:data<=-16'd7121;
      123471:data<=-16'd7533;
      123472:data<=-16'd7194;
      123473:data<=-16'd6783;
      123474:data<=-16'd6496;
      123475:data<=-16'd6868;
      123476:data<=-16'd8561;
      123477:data<=-16'd8833;
      123478:data<=-16'd7853;
      123479:data<=-16'd7985;
      123480:data<=-16'd7705;
      123481:data<=-16'd7165;
      123482:data<=-16'd7500;
      123483:data<=-16'd8467;
      123484:data<=-16'd9467;
      123485:data<=-16'd8287;
      123486:data<=-16'd7821;
      123487:data<=-16'd9060;
      123488:data<=-16'd4006;
      123489:data<=16'd3548;
      123490:data<=16'd3894;
      123491:data<=16'd2261;
      123492:data<=16'd2425;
      123493:data<=16'd1992;
      123494:data<=16'd2507;
      123495:data<=16'd1562;
      123496:data<=-16'd1791;
      123497:data<=-16'd2526;
      123498:data<=-16'd1744;
      123499:data<=-16'd2326;
      123500:data<=-16'd2673;
      123501:data<=-16'd2629;
      123502:data<=-16'd3297;
      123503:data<=-16'd4484;
      123504:data<=-16'd5010;
      123505:data<=-16'd4814;
      123506:data<=-16'd4957;
      123507:data<=-16'd4670;
      123508:data<=-16'd4717;
      123509:data<=-16'd6398;
      123510:data<=-16'd6845;
      123511:data<=-16'd5938;
      123512:data<=-16'd6176;
      123513:data<=-16'd5914;
      123514:data<=-16'd4989;
      123515:data<=-16'd5800;
      123516:data<=-16'd7247;
      123517:data<=-16'd7086;
      123518:data<=-16'd6291;
      123519:data<=-16'd6714;
      123520:data<=-16'd6930;
      123521:data<=-16'd6363;
      123522:data<=-16'd7254;
      123523:data<=-16'd8305;
      123524:data<=-16'd8396;
      123525:data<=-16'd8364;
      123526:data<=-16'd7133;
      123527:data<=-16'd7127;
      123528:data<=-16'd8014;
      123529:data<=-16'd6931;
      123530:data<=-16'd11414;
      123531:data<=-16'd20269;
      123532:data<=-16'd21262;
      123533:data<=-16'd18639;
      123534:data<=-16'd18618;
      123535:data<=-16'd18142;
      123536:data<=-16'd18976;
      123537:data<=-16'd19355;
      123538:data<=-16'd17462;
      123539:data<=-16'd17370;
      123540:data<=-16'd16607;
      123541:data<=-16'd14986;
      123542:data<=-16'd15803;
      123543:data<=-16'd15969;
      123544:data<=-16'd15286;
      123545:data<=-16'd14172;
      123546:data<=-16'd11635;
      123547:data<=-16'd10939;
      123548:data<=-16'd11342;
      123549:data<=-16'd11121;
      123550:data<=-16'd11147;
      123551:data<=-16'd10181;
      123552:data<=-16'd9964;
      123553:data<=-16'd10223;
      123554:data<=-16'd8775;
      123555:data<=-16'd9042;
      123556:data<=-16'd9919;
      123557:data<=-16'd8953;
      123558:data<=-16'd8889;
      123559:data<=-16'd8608;
      123560:data<=-16'd7609;
      123561:data<=-16'd7326;
      123562:data<=-16'd6428;
      123563:data<=-16'd5494;
      123564:data<=-16'd4905;
      123565:data<=-16'd4438;
      123566:data<=-16'd4147;
      123567:data<=-16'd3548;
      123568:data<=-16'd3553;
      123569:data<=-16'd1384;
      123570:data<=16'd937;
      123571:data<=-16'd1917;
      123572:data<=16'd1286;
      123573:data<=16'd12035;
      123574:data<=16'd13969;
      123575:data<=16'd11961;
      123576:data<=16'd14280;
      123577:data<=16'd13979;
      123578:data<=16'd13191;
      123579:data<=16'd13882;
      123580:data<=16'd12828;
      123581:data<=16'd12868;
      123582:data<=16'd13377;
      123583:data<=16'd13127;
      123584:data<=16'd13265;
      123585:data<=16'd12622;
      123586:data<=16'd12176;
      123587:data<=16'd11426;
      123588:data<=16'd10824;
      123589:data<=16'd12718;
      123590:data<=16'd13106;
      123591:data<=16'd11556;
      123592:data<=16'd11529;
      123593:data<=16'd11336;
      123594:data<=16'd10950;
      123595:data<=16'd10598;
      123596:data<=16'd9919;
      123597:data<=16'd10358;
      123598:data<=16'd10088;
      123599:data<=16'd8989;
      123600:data<=16'd8536;
      123601:data<=16'd8258;
      123602:data<=16'd9347;
      123603:data<=16'd9812;
      123604:data<=16'd8672;
      123605:data<=16'd8581;
      123606:data<=16'd7674;
      123607:data<=16'd6848;
      123608:data<=16'd7817;
      123609:data<=16'd8094;
      123610:data<=16'd8586;
      123611:data<=16'd7688;
      123612:data<=16'd6451;
      123613:data<=16'd8627;
      123614:data<=16'd4733;
      123615:data<=-16'd4520;
      123616:data<=-16'd5332;
      123617:data<=-16'd2971;
      123618:data<=-16'd3864;
      123619:data<=-16'd3592;
      123620:data<=-16'd4011;
      123621:data<=-16'd4134;
      123622:data<=-16'd1988;
      123623:data<=-16'd1541;
      123624:data<=-16'd1704;
      123625:data<=-16'd1171;
      123626:data<=-16'd1453;
      123627:data<=-16'd1478;
      123628:data<=-16'd732;
      123629:data<=16'd696;
      123630:data<=16'd1386;
      123631:data<=16'd722;
      123632:data<=16'd1011;
      123633:data<=16'd1186;
      123634:data<=16'd761;
      123635:data<=16'd1824;
      123636:data<=16'd2817;
      123637:data<=16'd2914;
      123638:data<=16'd2632;
      123639:data<=16'd1660;
      123640:data<=16'd1319;
      123641:data<=16'd2061;
      123642:data<=16'd3563;
      123643:data<=16'd4294;
      123644:data<=16'd3239;
      123645:data<=16'd4055;
      123646:data<=16'd5821;
      123647:data<=16'd5239;
      123648:data<=16'd5844;
      123649:data<=16'd7251;
      123650:data<=16'd7065;
      123651:data<=16'd7222;
      123652:data<=16'd6502;
      123653:data<=16'd5832;
      123654:data<=16'd6196;
      123655:data<=16'd5412;
      123656:data<=16'd9615;
      123657:data<=16'd18354;
      123658:data<=16'd20124;
      123659:data<=16'd17720;
      123660:data<=16'd17770;
      123661:data<=16'd17444;
      123662:data<=16'd17452;
      123663:data<=16'd17638;
      123664:data<=16'd16164;
      123665:data<=16'd15723;
      123666:data<=16'd15245;
      123667:data<=16'd13584;
      123668:data<=16'd12998;
      123669:data<=16'd12179;
      123670:data<=16'd11030;
      123671:data<=16'd10660;
      123672:data<=16'd9721;
      123673:data<=16'd9053;
      123674:data<=16'd8648;
      123675:data<=16'd7068;
      123676:data<=16'd5715;
      123677:data<=16'd5059;
      123678:data<=16'd4490;
      123679:data<=16'd4238;
      123680:data<=16'd3941;
      123681:data<=16'd3228;
      123682:data<=16'd1621;
      123683:data<=16'd164;
      123684:data<=16'd256;
      123685:data<=16'd162;
      123686:data<=-16'd522;
      123687:data<=-16'd743;
      123688:data<=-16'd1601;
      123689:data<=-16'd2960;
      123690:data<=-16'd3689;
      123691:data<=-16'd3835;
      123692:data<=-16'd4053;
      123693:data<=-16'd4364;
      123694:data<=-16'd4020;
      123695:data<=-16'd5203;
      123696:data<=-16'd6901;
      123697:data<=-16'd5383;
      123698:data<=-16'd8304;
      123699:data<=-16'd17279;
      123700:data<=-16'd19408;
      123701:data<=-16'd17587;
      123702:data<=-16'd19881;
      123703:data<=-16'd19911;
      123704:data<=-16'd18460;
      123705:data<=-16'd19384;
      123706:data<=-16'd18478;
      123707:data<=-16'd17262;
      123708:data<=-16'd17879;
      123709:data<=-16'd18026;
      123710:data<=-16'd17841;
      123711:data<=-16'd17303;
      123712:data<=-16'd16425;
      123713:data<=-16'd15474;
      123714:data<=-16'd14997;
      123715:data<=-16'd16325;
      123716:data<=-16'd16782;
      123717:data<=-16'd15499;
      123718:data<=-16'd15100;
      123719:data<=-16'd14173;
      123720:data<=-16'd13050;
      123721:data<=-16'd13805;
      123722:data<=-16'd14963;
      123723:data<=-16'd15365;
      123724:data<=-16'd14387;
      123725:data<=-16'd13368;
      123726:data<=-16'd13408;
      123727:data<=-16'd12609;
      123728:data<=-16'd12831;
      123729:data<=-16'd14214;
      123730:data<=-16'd13420;
      123731:data<=-16'd12499;
      123732:data<=-16'd12040;
      123733:data<=-16'd10948;
      123734:data<=-16'd10945;
      123735:data<=-16'd11426;
      123736:data<=-16'd11970;
      123737:data<=-16'd11072;
      123738:data<=-16'd9323;
      123739:data<=-16'd10619;
      123740:data<=-16'd7315;
      123741:data<=16'd2014;
      123742:data<=16'd3633;
      123743:data<=16'd1328;
      123744:data<=16'd3086;
      123745:data<=16'd2552;
      123746:data<=16'd1939;
      123747:data<=16'd3450;
      123748:data<=16'd1812;
      123749:data<=16'd256;
      123750:data<=16'd823;
      123751:data<=16'd804;
      123752:data<=16'd981;
      123753:data<=16'd1327;
      123754:data<=16'd934;
      123755:data<=-16'd534;
      123756:data<=-16'd1468;
      123757:data<=-16'd456;
      123758:data<=-16'd546;
      123759:data<=-16'd1081;
      123760:data<=-16'd279;
      123761:data<=-16'd1216;
      123762:data<=-16'd2402;
      123763:data<=-16'd1999;
      123764:data<=-16'd2052;
      123765:data<=-16'd1677;
      123766:data<=-16'd1110;
      123767:data<=-16'd1428;
      123768:data<=-16'd1930;
      123769:data<=-16'd2487;
      123770:data<=-16'd1958;
      123771:data<=-16'd1480;
      123772:data<=-16'd2036;
      123773:data<=-16'd1592;
      123774:data<=-16'd1707;
      123775:data<=-16'd2067;
      123776:data<=-16'd958;
      123777:data<=-16'd970;
      123778:data<=-16'd779;
      123779:data<=-16'd293;
      123780:data<=-16'd1010;
      123781:data<=16'd919;
      123782:data<=-16'd65;
      123783:data<=-16'd8358;
      123784:data<=-16'd12010;
      123785:data<=-16'd9620;
      123786:data<=-16'd9738;
      123787:data<=-16'd9586;
      123788:data<=-16'd7509;
      123789:data<=-16'd6604;
      123790:data<=-16'd5750;
      123791:data<=-16'd4698;
      123792:data<=-16'd4566;
      123793:data<=-16'd4616;
      123794:data<=-16'd3755;
      123795:data<=-16'd2334;
      123796:data<=-16'd1636;
      123797:data<=-16'd1128;
      123798:data<=-16'd484;
      123799:data<=-16'd434;
      123800:data<=-16'd88;
      123801:data<=16'd731;
      123802:data<=16'd1541;
      123803:data<=16'd2478;
      123804:data<=16'd2892;
      123805:data<=16'd2820;
      123806:data<=16'd2473;
      123807:data<=16'd2476;
      123808:data<=16'd4077;
      123809:data<=16'd5422;
      123810:data<=16'd5353;
      123811:data<=16'd5379;
      123812:data<=16'd5042;
      123813:data<=16'd4770;
      123814:data<=16'd5799;
      123815:data<=16'd7110;
      123816:data<=16'd7803;
      123817:data<=16'd7274;
      123818:data<=16'd6775;
      123819:data<=16'd7003;
      123820:data<=16'd6061;
      123821:data<=16'd6830;
      123822:data<=16'd9106;
      123823:data<=16'd7827;
      123824:data<=16'd10213;
      123825:data<=16'd19047;
      123826:data<=16'd21704;
      123827:data<=16'd19767;
      123828:data<=16'd22016;
      123829:data<=16'd22891;
      123830:data<=16'd20903;
      123831:data<=16'd20686;
      123832:data<=16'd19983;
      123833:data<=16'd18571;
      123834:data<=16'd18915;
      123835:data<=16'd19314;
      123836:data<=16'd18707;
      123837:data<=16'd18290;
      123838:data<=16'd18116;
      123839:data<=16'd17177;
      123840:data<=16'd16114;
      123841:data<=16'd16433;
      123842:data<=16'd16904;
      123843:data<=16'd16369;
      123844:data<=16'd15929;
      123845:data<=16'd15352;
      123846:data<=16'd14261;
      123847:data<=16'd14183;
      123848:data<=16'd15249;
      123849:data<=16'd15238;
      123850:data<=16'd13797;
      123851:data<=16'd13267;
      123852:data<=16'd13345;
      123853:data<=16'd12578;
      123854:data<=16'd12622;
      123855:data<=16'd13309;
      123856:data<=16'd12789;
      123857:data<=16'd11926;
      123858:data<=16'd11124;
      123859:data<=16'd10164;
      123860:data<=16'd9641;
      123861:data<=16'd10085;
      123862:data<=16'd11442;
      123863:data<=16'd10921;
      123864:data<=16'd9336;
      123865:data<=16'd10373;
      123866:data<=16'd7711;
      123867:data<=-16'd1046;
      123868:data<=-16'd4854;
      123869:data<=-16'd3439;
      123870:data<=-16'd4175;
      123871:data<=-16'd4270;
      123872:data<=-16'd3162;
      123873:data<=-16'd3920;
      123874:data<=-16'd3692;
      123875:data<=-16'd2003;
      123876:data<=-16'd1494;
      123877:data<=-16'd1392;
      123878:data<=-16'd1196;
      123879:data<=-16'd1820;
      123880:data<=-16'd2455;
      123881:data<=-16'd2132;
      123882:data<=-16'd1974;
      123883:data<=-16'd2652;
      123884:data<=-16'd2993;
      123885:data<=-16'd2837;
      123886:data<=-16'd2880;
      123887:data<=-16'd3621;
      123888:data<=-16'd5090;
      123889:data<=-16'd5497;
      123890:data<=-16'd4786;
      123891:data<=-16'd5027;
      123892:data<=-16'd5494;
      123893:data<=-16'd5448;
      123894:data<=-16'd6028;
      123895:data<=-16'd7027;
      123896:data<=-16'd7570;
      123897:data<=-16'd7380;
      123898:data<=-16'd7177;
      123899:data<=-16'd7016;
      123900:data<=-16'd6467;
      123901:data<=-16'd7476;
      123902:data<=-16'd8924;
      123903:data<=-16'd8510;
      123904:data<=-16'd9207;
      123905:data<=-16'd9374;
      123906:data<=-16'd7456;
      123907:data<=-16'd9148;
      123908:data<=-16'd8692;
      123909:data<=16'd159;
      123910:data<=16'd5442;
      123911:data<=16'd3736;
      123912:data<=16'd3659;
      123913:data<=16'd3694;
      123914:data<=16'd2036;
      123915:data<=16'd1428;
      123916:data<=16'd699;
      123917:data<=-16'd123;
      123918:data<=16'd17;
      123919:data<=16'd205;
      123920:data<=-16'd291;
      123921:data<=-16'd2027;
      123922:data<=-16'd3439;
      123923:data<=-16'd3262;
      123924:data<=-16'd2969;
      123925:data<=-16'd2585;
      123926:data<=-16'd2199;
      123927:data<=-16'd3090;
      123928:data<=-16'd4435;
      123929:data<=-16'd4916;
      123930:data<=-16'd4731;
      123931:data<=-16'd4936;
      123932:data<=-16'd5181;
      123933:data<=-16'd4537;
      123934:data<=-16'd4805;
      123935:data<=-16'd6065;
      123936:data<=-16'd6223;
      123937:data<=-16'd6340;
      123938:data<=-16'd6566;
      123939:data<=-16'd6028;
      123940:data<=-16'd6361;
      123941:data<=-16'd7639;
      123942:data<=-16'd8508;
      123943:data<=-16'd8244;
      123944:data<=-16'd7385;
      123945:data<=-16'd7265;
      123946:data<=-16'd6677;
      123947:data<=-16'd6663;
      123948:data<=-16'd8578;
      123949:data<=-16'd8170;
      123950:data<=-16'd9121;
      123951:data<=-16'd16838;
      123952:data<=-16'd21728;
      123953:data<=-16'd20240;
      123954:data<=-16'd20221;
      123955:data<=-16'd20967;
      123956:data<=-16'd20307;
      123957:data<=-16'd19966;
      123958:data<=-16'd19106;
      123959:data<=-16'd18425;
      123960:data<=-16'd18680;
      123961:data<=-16'd18607;
      123962:data<=-16'd18037;
      123963:data<=-16'd17053;
      123964:data<=-16'd16340;
      123965:data<=-16'd15614;
      123966:data<=-16'd14354;
      123967:data<=-16'd14487;
      123968:data<=-16'd15402;
      123969:data<=-16'd15100;
      123970:data<=-16'd14352;
      123971:data<=-16'd13628;
      123972:data<=-16'd13044;
      123973:data<=-16'd12630;
      123974:data<=-16'd12642;
      123975:data<=-16'd13427;
      123976:data<=-16'd13044;
      123977:data<=-16'd11931;
      123978:data<=-16'd11779;
      123979:data<=-16'd11042;
      123980:data<=-16'd10804;
      123981:data<=-16'd11623;
      123982:data<=-16'd11168;
      123983:data<=-16'd10743;
      123984:data<=-16'd10458;
      123985:data<=-16'd9426;
      123986:data<=-16'd9154;
      123987:data<=-16'd8681;
      123988:data<=-16'd8370;
      123989:data<=-16'd8475;
      123990:data<=-16'd7200;
      123991:data<=-16'd6984;
      123992:data<=-16'd5071;
      123993:data<=16'd3145;
      123994:data<=16'd9636;
      123995:data<=16'd10146;
      123996:data<=16'd10270;
      123997:data<=16'd10439;
      123998:data<=16'd9696;
      123999:data<=16'd9612;
      124000:data<=16'd10499;
      124001:data<=16'd11935;
      124002:data<=16'd12258;
      124003:data<=16'd11486;
      124004:data<=16'd11153;
      124005:data<=16'd10610;
      124006:data<=16'd10061;
      124007:data<=16'd10583;
      124008:data<=16'd11433;
      124009:data<=16'd11577;
      124010:data<=16'd11430;
      124011:data<=16'd11803;
      124012:data<=16'd11573;
      124013:data<=16'd11151;
      124014:data<=16'd12349;
      124015:data<=16'd12739;
      124016:data<=16'd11634;
      124017:data<=16'd11473;
      124018:data<=16'd11016;
      124019:data<=16'd10445;
      124020:data<=16'd11394;
      124021:data<=16'd12107;
      124022:data<=16'd12135;
      124023:data<=16'd12052;
      124024:data<=16'd11590;
      124025:data<=16'd11174;
      124026:data<=16'd10766;
      124027:data<=16'd10897;
      124028:data<=16'd11204;
      124029:data<=16'd10818;
      124030:data<=16'd11479;
      124031:data<=16'd11840;
      124032:data<=16'd10302;
      124033:data<=16'd10756;
      124034:data<=16'd10856;
      124035:data<=16'd4548;
      124036:data<=-16'd2329;
      124037:data<=-16'd2996;
      124038:data<=-16'd2173;
      124039:data<=-16'd2819;
      124040:data<=-16'd1478;
      124041:data<=16'd682;
      124042:data<=16'd717;
      124043:data<=16'd381;
      124044:data<=16'd711;
      124045:data<=16'd864;
      124046:data<=16'd992;
      124047:data<=16'd1645;
      124048:data<=16'd3095;
      124049:data<=16'd3829;
      124050:data<=16'd3334;
      124051:data<=16'd3286;
      124052:data<=16'd3046;
      124053:data<=16'd3106;
      124054:data<=16'd4825;
      124055:data<=16'd5197;
      124056:data<=16'd4021;
      124057:data<=16'd4115;
      124058:data<=16'd4228;
      124059:data<=16'd3723;
      124060:data<=16'd4015;
      124061:data<=16'd4905;
      124062:data<=16'd5407;
      124063:data<=16'd5039;
      124064:data<=16'd4802;
      124065:data<=16'd4775;
      124066:data<=16'd4225;
      124067:data<=16'd4701;
      124068:data<=16'd5823;
      124069:data<=16'd5676;
      124070:data<=16'd5539;
      124071:data<=16'd5711;
      124072:data<=16'd4648;
      124073:data<=16'd4123;
      124074:data<=16'd5683;
      124075:data<=16'd5815;
      124076:data<=16'd5480;
      124077:data<=16'd11535;
      124078:data<=16'd18697;
      124079:data<=16'd18202;
      124080:data<=16'd16850;
      124081:data<=16'd18495;
      124082:data<=16'd18114;
      124083:data<=16'd17082;
      124084:data<=16'd16142;
      124085:data<=16'd14613;
      124086:data<=16'd14706;
      124087:data<=16'd14912;
      124088:data<=16'd14568;
      124089:data<=16'd13764;
      124090:data<=16'd11762;
      124091:data<=16'd11699;
      124092:data<=16'd12516;
      124093:data<=16'd11586;
      124094:data<=16'd11088;
      124095:data<=16'd9969;
      124096:data<=16'd8366;
      124097:data<=16'd8290;
      124098:data<=16'd7705;
      124099:data<=16'd6677;
      124100:data<=16'd5265;
      124101:data<=16'd3465;
      124102:data<=16'd3512;
      124103:data<=16'd2849;
      124104:data<=16'd1080;
      124105:data<=16'd1259;
      124106:data<=16'd1025;
      124107:data<=-16'd447;
      124108:data<=-16'd1660;
      124109:data<=-16'd2431;
      124110:data<=-16'd2056;
      124111:data<=-16'd1850;
      124112:data<=-16'd2000;
      124113:data<=-16'd2739;
      124114:data<=-16'd4939;
      124115:data<=-16'd5225;
      124116:data<=-16'd4790;
      124117:data<=-16'd5463;
      124118:data<=-16'd5218;
      124119:data<=-16'd10061;
      124120:data<=-16'd18607;
      124121:data<=-16'd20415;
      124122:data<=-16'd19420;
      124123:data<=-16'd19708;
      124124:data<=-16'd18468;
      124125:data<=-16'd18158;
      124126:data<=-16'd18296;
      124127:data<=-16'd18269;
      124128:data<=-16'd19159;
      124129:data<=-16'd17964;
      124130:data<=-16'd16669;
      124131:data<=-16'd16600;
      124132:data<=-16'd15226;
      124133:data<=-16'd15544;
      124134:data<=-16'd17083;
      124135:data<=-16'd16663;
      124136:data<=-16'd15910;
      124137:data<=-16'd14883;
      124138:data<=-16'd14155;
      124139:data<=-16'd14324;
      124140:data<=-16'd13900;
      124141:data<=-16'd14280;
      124142:data<=-16'd15120;
      124143:data<=-16'd14969;
      124144:data<=-16'd14528;
      124145:data<=-16'd12904;
      124146:data<=-16'd12135;
      124147:data<=-16'd14011;
      124148:data<=-16'd14807;
      124149:data<=-16'd14082;
      124150:data<=-16'd13809;
      124151:data<=-16'd13471;
      124152:data<=-16'd13039;
      124153:data<=-16'd13024;
      124154:data<=-16'd13379;
      124155:data<=-16'd12930;
      124156:data<=-16'd12460;
      124157:data<=-16'd13177;
      124158:data<=-16'd11819;
      124159:data<=-16'd10580;
      124160:data<=-16'd12225;
      124161:data<=-16'd7970;
      124162:data<=16'd731;
      124163:data<=16'd2405;
      124164:data<=16'd1337;
      124165:data<=16'd2763;
      124166:data<=16'd1970;
      124167:data<=16'd318;
      124168:data<=16'd408;
      124169:data<=16'd267;
      124170:data<=-16'd3;
      124171:data<=16'd190;
      124172:data<=16'd478;
      124173:data<=-16'd32;
      124174:data<=-16'd1386;
      124175:data<=-16'd1406;
      124176:data<=-16'd863;
      124177:data<=-16'd1439;
      124178:data<=-16'd1269;
      124179:data<=-16'd919;
      124180:data<=-16'd2052;
      124181:data<=-16'd2766;
      124182:data<=-16'd2517;
      124183:data<=-16'd2220;
      124184:data<=-16'd1645;
      124185:data<=-16'd1477;
      124186:data<=-16'd2258;
      124187:data<=-16'd3168;
      124188:data<=-16'd3383;
      124189:data<=-16'd2810;
      124190:data<=-16'd2505;
      124191:data<=-16'd2582;
      124192:data<=-16'd1900;
      124193:data<=-16'd1535;
      124194:data<=-16'd2778;
      124195:data<=-16'd3494;
      124196:data<=-16'd2460;
      124197:data<=-16'd1971;
      124198:data<=-16'd2036;
      124199:data<=-16'd1251;
      124200:data<=-16'd1798;
      124201:data<=-16'd2367;
      124202:data<=-16'd664;
      124203:data<=-16'd3961;
      124204:data<=-16'd12562;
      124205:data<=-16'd15041;
      124206:data<=-16'd12604;
      124207:data<=-16'd11975;
      124208:data<=-16'd10678;
      124209:data<=-16'd9415;
      124210:data<=-16'd9503;
      124211:data<=-16'd8486;
      124212:data<=-16'd7615;
      124213:data<=-16'd6167;
      124214:data<=-16'd3485;
      124215:data<=-16'd3010;
      124216:data<=-16'd3388;
      124217:data<=-16'd2914;
      124218:data<=-16'd2975;
      124219:data<=-16'd2303;
      124220:data<=-16'd849;
      124221:data<=16'd325;
      124222:data<=16'd1498;
      124223:data<=16'd1864;
      124224:data<=16'd1439;
      124225:data<=16'd1336;
      124226:data<=16'd2191;
      124227:data<=16'd3130;
      124228:data<=16'd2845;
      124229:data<=16'd3131;
      124230:data<=16'd4115;
      124231:data<=16'd3852;
      124232:data<=16'd4012;
      124233:data<=16'd4992;
      124234:data<=16'd5560;
      124235:data<=16'd6026;
      124236:data<=16'd6155;
      124237:data<=16'd6551;
      124238:data<=16'd6722;
      124239:data<=16'd6734;
      124240:data<=16'd8026;
      124241:data<=16'd7843;
      124242:data<=16'd7406;
      124243:data<=16'd8304;
      124244:data<=16'd6620;
      124245:data<=16'd9914;
      124246:data<=16'd20360;
      124247:data<=16'd23234;
      124248:data<=16'd20709;
      124249:data<=16'd21487;
      124250:data<=16'd20748;
      124251:data<=16'd19646;
      124252:data<=16'd19942;
      124253:data<=16'd19478;
      124254:data<=16'd20679;
      124255:data<=16'd20921;
      124256:data<=16'd19146;
      124257:data<=16'd18721;
      124258:data<=16'd17423;
      124259:data<=16'd16448;
      124260:data<=16'd17711;
      124261:data<=16'd18204;
      124262:data<=16'd18234;
      124263:data<=16'd17605;
      124264:data<=16'd15985;
      124265:data<=16'd15338;
      124266:data<=16'd15230;
      124267:data<=16'd15882;
      124268:data<=16'd16301;
      124269:data<=16'd15500;
      124270:data<=16'd15700;
      124271:data<=16'd14739;
      124272:data<=16'd12427;
      124273:data<=16'd12982;
      124274:data<=16'd14032;
      124275:data<=16'd13562;
      124276:data<=16'd13467;
      124277:data<=16'd13171;
      124278:data<=16'd12276;
      124279:data<=16'd11935;
      124280:data<=16'd12991;
      124281:data<=16'd12648;
      124282:data<=16'd10316;
      124283:data<=16'd11306;
      124284:data<=16'd12058;
      124285:data<=16'd10025;
      124286:data<=16'd11649;
      124287:data<=16'd8860;
      124288:data<=-16'd1729;
      124289:data<=-16'd4598;
      124290:data<=-16'd2231;
      124291:data<=-16'd4132;
      124292:data<=-16'd3882;
      124293:data<=-16'd1347;
      124294:data<=-16'd831;
      124295:data<=-16'd1040;
      124296:data<=-16'd2237;
      124297:data<=-16'd2690;
      124298:data<=-16'd1635;
      124299:data<=-16'd1005;
      124300:data<=16'd281;
      124301:data<=16'd1293;
      124302:data<=16'd704;
      124303:data<=16'd146;
      124304:data<=-16'd355;
      124305:data<=-16'd704;
      124306:data<=-16'd466;
      124307:data<=-16'd244;
      124308:data<=-16'd115;
      124309:data<=-16'd372;
      124310:data<=-16'd936;
      124311:data<=-16'd1474;
      124312:data<=-16'd1939;
      124313:data<=-16'd2399;
      124314:data<=-16'd3181;
      124315:data<=-16'd3321;
      124316:data<=-16'd3436;
      124317:data<=-16'd4432;
      124318:data<=-16'd4111;
      124319:data<=-16'd4358;
      124320:data<=-16'd6170;
      124321:data<=-16'd5782;
      124322:data<=-16'd5551;
      124323:data<=-16'd5827;
      124324:data<=-16'd4328;
      124325:data<=-16'd5582;
      124326:data<=-16'd6980;
      124327:data<=-16'd6155;
      124328:data<=-16'd8062;
      124329:data<=-16'd4892;
      124330:data<=16'd4613;
      124331:data<=16'd6572;
      124332:data<=16'd4074;
      124333:data<=16'd3980;
      124334:data<=16'd2507;
      124335:data<=16'd2152;
      124336:data<=16'd2922;
      124337:data<=16'd1779;
      124338:data<=16'd1933;
      124339:data<=16'd1513;
      124340:data<=-16'd804;
      124341:data<=-16'd826;
      124342:data<=-16'd193;
      124343:data<=-16'd678;
      124344:data<=-16'd1111;
      124345:data<=-16'd2118;
      124346:data<=-16'd2635;
      124347:data<=-16'd2819;
      124348:data<=-16'd4211;
      124349:data<=-16'd4681;
      124350:data<=-16'd3498;
      124351:data<=-16'd2884;
      124352:data<=-16'd3495;
      124353:data<=-16'd4552;
      124354:data<=-16'd4998;
      124355:data<=-16'd4842;
      124356:data<=-16'd5086;
      124357:data<=-16'd5439;
      124358:data<=-16'd5221;
      124359:data<=-16'd5328;
      124360:data<=-16'd6396;
      124361:data<=-16'd7370;
      124362:data<=-16'd7984;
      124363:data<=-16'd8325;
      124364:data<=-16'd7636;
      124365:data<=-16'd7456;
      124366:data<=-16'd8419;
      124367:data<=-16'd8405;
      124368:data<=-16'd8493;
      124369:data<=-16'd8284;
      124370:data<=-16'd6047;
      124371:data<=-16'd8190;
      124372:data<=-16'd16172;
      124373:data<=-16'd20158;
      124374:data<=-16'd18813;
      124375:data<=-16'd18205;
      124376:data<=-16'd18345;
      124377:data<=-16'd17719;
      124378:data<=-16'd16718;
      124379:data<=-16'd16378;
      124380:data<=-16'd17432;
      124381:data<=-16'd17572;
      124382:data<=-16'd16199;
      124383:data<=-16'd16134;
      124384:data<=-16'd16148;
      124385:data<=-16'd14176;
      124386:data<=-16'd13521;
      124387:data<=-16'd14783;
      124388:data<=-16'd13994;
      124389:data<=-16'd12592;
      124390:data<=-16'd12922;
      124391:data<=-16'd12298;
      124392:data<=-16'd12003;
      124393:data<=-16'd13418;
      124394:data<=-16'd12787;
      124395:data<=-16'd11779;
      124396:data<=-16'd12464;
      124397:data<=-16'd11984;
      124398:data<=-16'd11491;
      124399:data<=-16'd11573;
      124400:data<=-16'd11453;
      124401:data<=-16'd12182;
      124402:data<=-16'd11062;
      124403:data<=-16'd9520;
      124404:data<=-16'd10251;
      124405:data<=-16'd9254;
      124406:data<=-16'd9227;
      124407:data<=-16'd11004;
      124408:data<=-16'd8940;
      124409:data<=-16'd8025;
      124410:data<=-16'd9007;
      124411:data<=-16'd7881;
      124412:data<=-16'd8804;
      124413:data<=-16'd5507;
      124414:data<=16'd3472;
      124415:data<=16'd5018;
      124416:data<=16'd3698;
      124417:data<=16'd5315;
      124418:data<=16'd4032;
      124419:data<=16'd4787;
      124420:data<=16'd7373;
      124421:data<=16'd6267;
      124422:data<=16'd6910;
      124423:data<=16'd7834;
      124424:data<=16'd5832;
      124425:data<=16'd6247;
      124426:data<=16'd7893;
      124427:data<=16'd7785;
      124428:data<=16'd7670;
      124429:data<=16'd8035;
      124430:data<=16'd8061;
      124431:data<=16'd7295;
      124432:data<=16'd7929;
      124433:data<=16'd9462;
      124434:data<=16'd8856;
      124435:data<=16'd8772;
      124436:data<=16'd9435;
      124437:data<=16'd8583;
      124438:data<=16'd8458;
      124439:data<=16'd8940;
      124440:data<=16'd9905;
      124441:data<=16'd10930;
      124442:data<=16'd9565;
      124443:data<=16'd9078;
      124444:data<=16'd9473;
      124445:data<=16'd8337;
      124446:data<=16'd9582;
      124447:data<=16'd11274;
      124448:data<=16'd10989;
      124449:data<=16'd11207;
      124450:data<=16'd10103;
      124451:data<=16'd9536;
      124452:data<=16'd10351;
      124453:data<=16'd9846;
      124454:data<=16'd11210;
      124455:data<=16'd9159;
      124456:data<=16'd626;
      124457:data<=-16'd2593;
      124458:data<=-16'd1724;
      124459:data<=-16'd2352;
      124460:data<=-16'd340;
      124461:data<=16'd206;
      124462:data<=-16'd1315;
      124463:data<=16'd3;
      124464:data<=16'd183;
      124465:data<=-16'd6;
      124466:data<=16'd1933;
      124467:data<=16'd2560;
      124468:data<=16'd2637;
      124469:data<=16'd2460;
      124470:data<=16'd1842;
      124471:data<=16'd2786;
      124472:data<=16'd3083;
      124473:data<=16'd2734;
      124474:data<=16'd3557;
      124475:data<=16'd3427;
      124476:data<=16'd2913;
      124477:data<=16'd3566;
      124478:data<=16'd4249;
      124479:data<=16'd4443;
      124480:data<=16'd4353;
      124481:data<=16'd4528;
      124482:data<=16'd4648;
      124483:data<=16'd4470;
      124484:data<=16'd4660;
      124485:data<=16'd4746;
      124486:data<=16'd5429;
      124487:data<=16'd6326;
      124488:data<=16'd5509;
      124489:data<=16'd5083;
      124490:data<=16'd5280;
      124491:data<=16'd4273;
      124492:data<=16'd4400;
      124493:data<=16'd5703;
      124494:data<=16'd6528;
      124495:data<=16'd6701;
      124496:data<=16'd5891;
      124497:data<=16'd8420;
      124498:data<=16'd14851;
      124499:data<=16'd17471;
      124500:data<=16'd16536;
      124501:data<=16'd16601;
      124502:data<=16'd16052;
      124503:data<=16'd15145;
      124504:data<=16'd15197;
      124505:data<=16'd14995;
      124506:data<=16'd15064;
      124507:data<=16'd14962;
      124508:data<=16'd13558;
      124509:data<=16'd12777;
      124510:data<=16'd12592;
      124511:data<=16'd11113;
      124512:data<=16'd10619;
      124513:data<=16'd12152;
      124514:data<=16'd11973;
      124515:data<=16'd10293;
      124516:data<=16'd9818;
      124517:data<=16'd9312;
      124518:data<=16'd8825;
      124519:data<=16'd9104;
      124520:data<=16'd8442;
      124521:data<=16'd7685;
      124522:data<=16'd7471;
      124523:data<=16'd6401;
      124524:data<=16'd5706;
      124525:data<=16'd5521;
      124526:data<=16'd4087;
      124527:data<=16'd2191;
      124528:data<=16'd1365;
      124529:data<=16'd1764;
      124530:data<=16'd1817;
      124531:data<=16'd776;
      124532:data<=16'd61;
      124533:data<=-16'd837;
      124534:data<=-16'd1830;
      124535:data<=-16'd1663;
      124536:data<=-16'd2326;
      124537:data<=-16'd2826;
      124538:data<=-16'd2174;
      124539:data<=-16'd6435;
      124540:data<=-16'd13952;
      124541:data<=-16'd15923;
      124542:data<=-16'd14721;
      124543:data<=-16'd15039;
      124544:data<=-16'd14797;
      124545:data<=-16'd15094;
      124546:data<=-16'd16653;
      124547:data<=-16'd16302;
      124548:data<=-16'd15424;
      124549:data<=-16'd15402;
      124550:data<=-16'd14160;
      124551:data<=-16'd13571;
      124552:data<=-16'd14803;
      124553:data<=-16'd14903;
      124554:data<=-16'd14487;
      124555:data<=-16'd14838;
      124556:data<=-16'd14207;
      124557:data<=-16'd13168;
      124558:data<=-16'd13295;
      124559:data<=-16'd14107;
      124560:data<=-16'd14445;
      124561:data<=-16'd13518;
      124562:data<=-16'd12630;
      124563:data<=-16'd12502;
      124564:data<=-16'd11902;
      124565:data<=-16'd12034;
      124566:data<=-16'd13098;
      124567:data<=-16'd12769;
      124568:data<=-16'd12220;
      124569:data<=-16'd12273;
      124570:data<=-16'd11479;
      124571:data<=-16'd11335;
      124572:data<=-16'd12404;
      124573:data<=-16'd13229;
      124574:data<=-16'd13743;
      124575:data<=-16'd12710;
      124576:data<=-16'd10948;
      124577:data<=-16'd11106;
      124578:data<=-16'd10978;
      124579:data<=-16'd10628;
      124580:data<=-16'd11999;
      124581:data<=-16'd9045;
      124582:data<=-16'd1046;
      124583:data<=16'd2739;
      124584:data<=16'd1830;
      124585:data<=16'd1166;
      124586:data<=16'd218;
      124587:data<=-16'd610;
      124588:data<=-16'd488;
      124589:data<=-16'd690;
      124590:data<=-16'd872;
      124591:data<=-16'd1086;
      124592:data<=-16'd1882;
      124593:data<=-16'd2475;
      124594:data<=-16'd2848;
      124595:data<=-16'd3472;
      124596:data<=-16'd3918;
      124597:data<=-16'd3137;
      124598:data<=-16'd2027;
      124599:data<=-16'd2558;
      124600:data<=-16'd2889;
      124601:data<=-16'd2203;
      124602:data<=-16'd2772;
      124603:data<=-16'd2989;
      124604:data<=-16'd2299;
      124605:data<=-16'd3209;
      124606:data<=-16'd4255;
      124607:data<=-16'd4302;
      124608:data<=-16'd4672;
      124609:data<=-16'd4992;
      124610:data<=-16'd4526;
      124611:data<=-16'd3603;
      124612:data<=-16'd3642;
      124613:data<=-16'd3786;
      124614:data<=-16'd2787;
      124615:data<=-16'd3697;
      124616:data<=-16'd4866;
      124617:data<=-16'd3294;
      124618:data<=-16'd3498;
      124619:data<=-16'd4884;
      124620:data<=-16'd4758;
      124621:data<=-16'd5150;
      124622:data<=-16'd4243;
      124623:data<=-16'd5779;
      124624:data<=-16'd12646;
      124625:data<=-16'd14651;
      124626:data<=-16'd12684;
      124627:data<=-16'd13952;
      124628:data<=-16'd13312;
      124629:data<=-16'd11556;
      124630:data<=-16'd11755;
      124631:data<=-16'd9706;
      124632:data<=-16'd7689;
      124633:data<=-16'd7385;
      124634:data<=-16'd6088;
      124635:data<=-16'd5416;
      124636:data<=-16'd5359;
      124637:data<=-16'd4974;
      124638:data<=-16'd4457;
      124639:data<=-16'd2596;
      124640:data<=-16'd1181;
      124641:data<=-16'd1162;
      124642:data<=-16'd886;
      124643:data<=-16'd955;
      124644:data<=-16'd682;
      124645:data<=16'd694;
      124646:data<=16'd1530;
      124647:data<=16'd1862;
      124648:data<=16'd2742;
      124649:data<=16'd3994;
      124650:data<=16'd4264;
      124651:data<=16'd3832;
      124652:data<=16'd4893;
      124653:data<=16'd6146;
      124654:data<=16'd5512;
      124655:data<=16'd4335;
      124656:data<=16'd4164;
      124657:data<=16'd5156;
      124658:data<=16'd5958;
      124659:data<=16'd6658;
      124660:data<=16'd7597;
      124661:data<=16'd6693;
      124662:data<=16'd6811;
      124663:data<=16'd8621;
      124664:data<=16'd6795;
      124665:data<=16'd7708;
      124666:data<=16'd15838;
      124667:data<=16'd20181;
      124668:data<=16'd18903;
      124669:data<=16'd17829;
      124670:data<=16'd16543;
      124671:data<=16'd16636;
      124672:data<=16'd18131;
      124673:data<=16'd18266;
      124674:data<=16'd17782;
      124675:data<=16'd16694;
      124676:data<=16'd15858;
      124677:data<=16'd16202;
      124678:data<=16'd16228;
      124679:data<=16'd16609;
      124680:data<=16'd16631;
      124681:data<=16'd15644;
      124682:data<=16'd15970;
      124683:data<=16'd15946;
      124684:data<=16'd15009;
      124685:data<=16'd15659;
      124686:data<=16'd16045;
      124687:data<=16'd15201;
      124688:data<=16'd14411;
      124689:data<=16'd13439;
      124690:data<=16'd12772;
      124691:data<=16'd12445;
      124692:data<=16'd12622;
      124693:data<=16'd13159;
      124694:data<=16'd12357;
      124695:data<=16'd11837;
      124696:data<=16'd12851;
      124697:data<=16'd13124;
      124698:data<=16'd12803;
      124699:data<=16'd12739;
      124700:data<=16'd12777;
      124701:data<=16'd12804;
      124702:data<=16'd11932;
      124703:data<=16'd11307;
      124704:data<=16'd11350;
      124705:data<=16'd11145;
      124706:data<=16'd11935;
      124707:data<=16'd10176;
      124708:data<=16'd3230;
      124709:data<=-16'd1293;
      124710:data<=-16'd914;
      124711:data<=-16'd787;
      124712:data<=-16'd626;
      124713:data<=16'd106;
      124714:data<=16'd50;
      124715:data<=16'd675;
      124716:data<=16'd1321;
      124717:data<=16'd520;
      124718:data<=16'd376;
      124719:data<=16'd1801;
      124720:data<=16'd2845;
      124721:data<=16'd2881;
      124722:data<=16'd3027;
      124723:data<=16'd3013;
      124724:data<=16'd2611;
      124725:data<=16'd3102;
      124726:data<=16'd3469;
      124727:data<=16'd2893;
      124728:data<=16'd3292;
      124729:data<=16'd3842;
      124730:data<=16'd3301;
      124731:data<=16'd2875;
      124732:data<=16'd2576;
      124733:data<=16'd3099;
      124734:data<=16'd3965;
      124735:data<=16'd3072;
      124736:data<=16'd2911;
      124737:data<=16'd3694;
      124738:data<=16'd1597;
      124739:data<=-16'd942;
      124740:data<=-16'd934;
      124741:data<=-16'd450;
      124742:data<=-16'd516;
      124743:data<=-16'd616;
      124744:data<=-16'd604;
      124745:data<=-16'd1692;
      124746:data<=-16'd3560;
      124747:data<=-16'd3418;
      124748:data<=-16'd3219;
      124749:data<=-16'd3075;
      124750:data<=16'd2203;
      124751:data<=16'd7679;
      124752:data<=16'd6572;
      124753:data<=16'd4443;
      124754:data<=16'd4663;
      124755:data<=16'd4176;
      124756:data<=16'd3551;
      124757:data<=16'd3812;
      124758:data<=16'd3054;
      124759:data<=16'd1195;
      124760:data<=16'd632;
      124761:data<=16'd895;
      124762:data<=16'd385;
      124763:data<=16'd282;
      124764:data<=-16'd403;
      124765:data<=-16'd2099;
      124766:data<=-16'd2058;
      124767:data<=-16'd1812;
      124768:data<=-16'd2209;
      124769:data<=-16'd1400;
      124770:data<=-16'd1430;
      124771:data<=-16'd2414;
      124772:data<=-16'd3444;
      124773:data<=-16'd5143;
      124774:data<=-16'd5121;
      124775:data<=-16'd4488;
      124776:data<=-16'd4931;
      124777:data<=-16'd3899;
      124778:data<=-16'd3811;
      124779:data<=-16'd5865;
      124780:data<=-16'd6860;
      124781:data<=-16'd7279;
      124782:data<=-16'd6722;
      124783:data<=-16'd6149;
      124784:data<=-16'd7785;
      124785:data<=-16'd8287;
      124786:data<=-16'd8147;
      124787:data<=-16'd9453;
      124788:data<=-16'd9236;
      124789:data<=-16'd8566;
      124790:data<=-16'd8483;
      124791:data<=-16'd9051;
      124792:data<=-16'd14019;
      124793:data<=-16'd19555;
      124794:data<=-16'd20284;
      124795:data<=-16'd20058;
      124796:data<=-16'd20037;
      124797:data<=-16'd18600;
      124798:data<=-16'd18083;
      124799:data<=-16'd18594;
      124800:data<=-16'd18222;
      124801:data<=-16'd17418;
      124802:data<=-16'd16785;
      124803:data<=-16'd15773;
      124804:data<=-16'd15343;
      124805:data<=-16'd16305;
      124806:data<=-16'd15702;
      124807:data<=-16'd13617;
      124808:data<=-16'd14057;
      124809:data<=-16'd14772;
      124810:data<=-16'd13327;
      124811:data<=-16'd13100;
      124812:data<=-16'd14013;
      124813:data<=-16'd14337;
      124814:data<=-16'd15088;
      124815:data<=-16'd15201;
      124816:data<=-16'd13547;
      124817:data<=-16'd11829;
      124818:data<=-16'd11972;
      124819:data<=-16'd13361;
      124820:data<=-16'd13282;
      124821:data<=-16'd12293;
      124822:data<=-16'd11864;
      124823:data<=-16'd10266;
      124824:data<=-16'd9100;
      124825:data<=-16'd9915;
      124826:data<=-16'd9659;
      124827:data<=-16'd9263;
      124828:data<=-16'd9790;
      124829:data<=-16'd8948;
      124830:data<=-16'd8728;
      124831:data<=-16'd9414;
      124832:data<=-16'd9236;
      124833:data<=-16'd9192;
      124834:data<=-16'd5330;
      124835:data<=16'd1774;
      124836:data<=16'd3570;
      124837:data<=16'd2529;
      124838:data<=16'd2896;
      124839:data<=16'd1639;
      124840:data<=16'd1839;
      124841:data<=16'd3938;
      124842:data<=16'd3074;
      124843:data<=16'd2217;
      124844:data<=16'd3620;
      124845:data<=16'd4664;
      124846:data<=16'd4905;
      124847:data<=16'd4730;
      124848:data<=16'd4942;
      124849:data<=16'd4913;
      124850:data<=16'd4317;
      124851:data<=16'd5627;
      124852:data<=16'd7460;
      124853:data<=16'd7903;
      124854:data<=16'd8073;
      124855:data<=16'd7101;
      124856:data<=16'd5950;
      124857:data<=16'd6234;
      124858:data<=16'd6667;
      124859:data<=16'd7538;
      124860:data<=16'd8466;
      124861:data<=16'd8278;
      124862:data<=16'd7680;
      124863:data<=16'd7036;
      124864:data<=16'd7153;
      124865:data<=16'd7588;
      124866:data<=16'd7291;
      124867:data<=16'd7541;
      124868:data<=16'd7911;
      124869:data<=16'd7403;
      124870:data<=16'd6648;
      124871:data<=16'd7037;
      124872:data<=16'd9420;
      124873:data<=16'd12712;
      124874:data<=16'd21035;
      124875:data<=16'd31172;
      124876:data<=16'd25047;
      124877:data<=16'd8370;
      124878:data<=16'd2957;
      124879:data<=16'd4447;
      124880:data<=16'd3944;
      124881:data<=16'd3242;
      124882:data<=16'd2472;
      124883:data<=16'd1633;
      124884:data<=-16'd5341;
      124885:data<=-16'd14425;
      124886:data<=-16'd13750;
      124887:data<=-16'd16418;
      124888:data<=-16'd27680;
      124889:data<=-16'd30644;
      124890:data<=-16'd27326;
      124891:data<=-16'd26462;
      124892:data<=-16'd25992;
      124893:data<=-16'd18988;
      124894:data<=-16'd3482;
      124895:data<=16'd1087;
      124896:data<=-16'd8109;
      124897:data<=-16'd8884;
      124898:data<=-16'd6557;
      124899:data<=-16'd8990;
      124900:data<=-16'd7300;
      124901:data<=-16'd6338;
      124902:data<=-16'd6220;
      124903:data<=-16'd4338;
      124904:data<=-16'd6278;
      124905:data<=-16'd5888;
      124906:data<=-16'd3533;
      124907:data<=-16'd4783;
      124908:data<=-16'd4017;
      124909:data<=-16'd3615;
      124910:data<=-16'd5068;
      124911:data<=-16'd5145;
      124912:data<=-16'd6100;
      124913:data<=-16'd4582;
      124914:data<=-16'd3028;
      124915:data<=-16'd4864;
      124916:data<=-16'd3497;
      124917:data<=-16'd2593;
      124918:data<=-16'd2889;
      124919:data<=-16'd1409;
      124920:data<=-16'd3406;
      124921:data<=16'd1906;
      124922:data<=16'd15288;
      124923:data<=16'd17054;
      124924:data<=16'd14267;
      124925:data<=16'd16578;
      124926:data<=16'd15597;
      124927:data<=16'd13744;
      124928:data<=16'd13088;
      124929:data<=16'd11903;
      124930:data<=16'd11768;
      124931:data<=16'd10116;
      124932:data<=16'd9241;
      124933:data<=16'd9761;
      124934:data<=16'd8871;
      124935:data<=16'd9908;
      124936:data<=16'd9808;
      124937:data<=16'd8172;
      124938:data<=16'd9125;
      124939:data<=16'd7653;
      124940:data<=16'd8768;
      124941:data<=16'd16402;
      124942:data<=16'd18322;
      124943:data<=16'd15406;
      124944:data<=16'd13963;
      124945:data<=16'd12022;
      124946:data<=16'd12326;
      124947:data<=16'd12751;
      124948:data<=16'd10810;
      124949:data<=16'd11408;
      124950:data<=16'd11779;
      124951:data<=16'd9750;
      124952:data<=16'd9315;
      124953:data<=16'd9747;
      124954:data<=16'd9806;
      124955:data<=16'd8983;
      124956:data<=16'd7216;
      124957:data<=16'd7453;
      124958:data<=16'd7021;
      124959:data<=-16'd485;
      124960:data<=-16'd10834;
      124961:data<=-16'd13934;
      124962:data<=-16'd11843;
      124963:data<=-16'd12140;
      124964:data<=-16'd11916;
      124965:data<=-16'd9539;
      124966:data<=-16'd9414;
      124967:data<=-16'd9817;
      124968:data<=-16'd9013;
      124969:data<=-16'd8554;
      124970:data<=-16'd8197;
      124971:data<=-16'd8267;
      124972:data<=-16'd7947;
      124973:data<=-16'd7060;
      124974:data<=-16'd6880;
      124975:data<=-16'd6692;
      124976:data<=-16'd7191;
      124977:data<=-16'd7765;
      124978:data<=-16'd7840;
      124979:data<=-16'd9142;
      124980:data<=-16'd8381;
      124981:data<=-16'd6663;
      124982:data<=-16'd7843;
      124983:data<=-16'd6816;
      124984:data<=-16'd6253;
      124985:data<=-16'd11235;
      124986:data<=-16'd14217;
      124987:data<=-16'd13485;
      124988:data<=-16'd12649;
      124989:data<=-16'd11162;
      124990:data<=-16'd10141;
      124991:data<=-16'd9438;
      124992:data<=-16'd8893;
      124993:data<=-16'd8598;
      124994:data<=-16'd9022;
      124995:data<=-16'd11515;
      124996:data<=-16'd7148;
      124997:data<=16'd5066;
      124998:data<=16'd9583;
      124999:data<=16'd8062;
      125000:data<=16'd8846;
      125001:data<=16'd7917;
      125002:data<=16'd7483;
      125003:data<=16'd8654;
      125004:data<=16'd7794;
      125005:data<=16'd7595;
      125006:data<=16'd7526;
      125007:data<=16'd6431;
      125008:data<=16'd6193;
      125009:data<=16'd6128;
      125010:data<=16'd6144;
      125011:data<=16'd4878;
      125012:data<=16'd3882;
      125013:data<=16'd5830;
      125014:data<=16'd5791;
      125015:data<=16'd4567;
      125016:data<=16'd5429;
      125017:data<=16'd4510;
      125018:data<=16'd3900;
      125019:data<=16'd4308;
      125020:data<=16'd2725;
      125021:data<=16'd3377;
      125022:data<=16'd4811;
      125023:data<=16'd3532;
      125024:data<=16'd3570;
      125025:data<=16'd4085;
      125026:data<=16'd3360;
      125027:data<=16'd2156;
      125028:data<=-16'd41;
      125029:data<=16'd2431;
      125030:data<=16'd9291;
      125031:data<=16'd10305;
      125032:data<=16'd8610;
      125033:data<=16'd9448;
      125034:data<=16'd2995;
      125035:data<=-16'd8407;
      125036:data<=-16'd10284;
      125037:data<=-16'd7366;
      125038:data<=-16'd8316;
      125039:data<=-16'd8393;
      125040:data<=-16'd7377;
      125041:data<=-16'd7136;
      125042:data<=-16'd6020;
      125043:data<=-16'd6625;
      125044:data<=-16'd8187;
      125045:data<=-16'd8052;
      125046:data<=-16'd7588;
      125047:data<=-16'd6634;
      125048:data<=-16'd6108;
      125049:data<=-16'd6138;
      125050:data<=-16'd5990;
      125051:data<=-16'd7338;
      125052:data<=-16'd6692;
      125053:data<=-16'd3861;
      125054:data<=-16'd3885;
      125055:data<=-16'd3877;
      125056:data<=-16'd3322;
      125057:data<=-16'd4059;
      125058:data<=-16'd3083;
      125059:data<=-16'd2519;
      125060:data<=-16'd3356;
      125061:data<=-16'd3676;
      125062:data<=-16'd4287;
      125063:data<=-16'd3368;
      125064:data<=-16'd2566;
      125065:data<=-16'd2977;
      125066:data<=-16'd1888;
      125067:data<=-16'd2482;
      125068:data<=-16'd2808;
      125069:data<=-16'd1343;
      125070:data<=-16'd2710;
      125071:data<=16'd2070;
      125072:data<=16'd14392;
      125073:data<=16'd17996;
      125074:data<=16'd12813;
      125075:data<=16'd8965;
      125076:data<=16'd8226;
      125077:data<=16'd8398;
      125078:data<=16'd7098;
      125079:data<=16'd5965;
      125080:data<=16'd5520;
      125081:data<=16'd4907;
      125082:data<=16'd5592;
      125083:data<=16'd5404;
      125084:data<=16'd5427;
      125085:data<=16'd6934;
      125086:data<=16'd5562;
      125087:data<=16'd4821;
      125088:data<=16'd6457;
      125089:data<=16'd5441;
      125090:data<=16'd4335;
      125091:data<=16'd4651;
      125092:data<=16'd4626;
      125093:data<=16'd4496;
      125094:data<=16'd3247;
      125095:data<=16'd3004;
      125096:data<=16'd3659;
      125097:data<=16'd2719;
      125098:data<=16'd2852;
      125099:data<=16'd3935;
      125100:data<=16'd4452;
      125101:data<=16'd4414;
      125102:data<=16'd3301;
      125103:data<=16'd3480;
      125104:data<=16'd3964;
      125105:data<=16'd3301;
      125106:data<=16'd3233;
      125107:data<=16'd3027;
      125108:data<=16'd3486;
      125109:data<=-16'd1027;
      125110:data<=-16'd13113;
      125111:data<=-16'd17535;
      125112:data<=-16'd14530;
      125113:data<=-16'd15706;
      125114:data<=-16'd15617;
      125115:data<=-16'd14201;
      125116:data<=-16'd15232;
      125117:data<=-16'd14081;
      125118:data<=-16'd10386;
      125119:data<=-16'd4508;
      125120:data<=-16'd881;
      125121:data<=-16'd2528;
      125122:data<=-16'd2306;
      125123:data<=-16'd1309;
      125124:data<=-16'd1864;
      125125:data<=-16'd1478;
      125126:data<=-16'd2214;
      125127:data<=-16'd1753;
      125128:data<=-16'd2044;
      125129:data<=-16'd4579;
      125130:data<=-16'd2038;
      125131:data<=-16'd325;
      125132:data<=-16'd1469;
      125133:data<=16'd767;
      125134:data<=-16'd836;
      125135:data<=-16'd2573;
      125136:data<=16'd1004;
      125137:data<=16'd763;
      125138:data<=-16'd397;
      125139:data<=-16'd317;
      125140:data<=-16'd1456;
      125141:data<=16'd381;
      125142:data<=16'd737;
      125143:data<=16'd726;
      125144:data<=16'd2569;
      125145:data<=-16'd782;
      125146:data<=16'd2541;
      125147:data<=16'd16446;
      125148:data<=16'd21362;
      125149:data<=16'd18763;
      125150:data<=16'd19126;
      125151:data<=16'd19287;
      125152:data<=16'd18525;
      125153:data<=16'd17796;
      125154:data<=16'd16666;
      125155:data<=16'd15734;
      125156:data<=16'd15526;
      125157:data<=16'd15675;
      125158:data<=16'd14486;
      125159:data<=16'd13837;
      125160:data<=16'd14040;
      125161:data<=16'd13940;
      125162:data<=16'd15929;
      125163:data<=16'd14425;
      125164:data<=16'd7668;
      125165:data<=16'd5465;
      125166:data<=16'd5905;
      125167:data<=16'd4636;
      125168:data<=16'd5412;
      125169:data<=16'd5932;
      125170:data<=16'd4805;
      125171:data<=16'd4517;
      125172:data<=16'd4463;
      125173:data<=16'd4437;
      125174:data<=16'd4188;
      125175:data<=16'd3671;
      125176:data<=16'd3694;
      125177:data<=16'd4679;
      125178:data<=16'd5876;
      125179:data<=16'd5808;
      125180:data<=16'd6247;
      125181:data<=16'd6073;
      125182:data<=16'd5016;
      125183:data<=16'd7081;
      125184:data<=16'd2161;
      125185:data<=-16'd11397;
      125186:data<=-16'd14446;
      125187:data<=-16'd10951;
      125188:data<=-16'd12225;
      125189:data<=-16'd11339;
      125190:data<=-16'd10185;
      125191:data<=-16'd10223;
      125192:data<=-16'd8448;
      125193:data<=-16'd9197;
      125194:data<=-16'd8325;
      125195:data<=-16'd5727;
      125196:data<=-16'd7294;
      125197:data<=-16'd7263;
      125198:data<=-16'd5873;
      125199:data<=-16'd6655;
      125200:data<=-16'd6341;
      125201:data<=-16'd5591;
      125202:data<=-16'd4361;
      125203:data<=-16'd4126;
      125204:data<=-16'd5231;
      125205:data<=-16'd3862;
      125206:data<=-16'd4399;
      125207:data<=-16'd4141;
      125208:data<=16'd2299;
      125209:data<=16'd5143;
      125210:data<=16'd5059;
      125211:data<=16'd7295;
      125212:data<=16'd6636;
      125213:data<=16'd6302;
      125214:data<=16'd7262;
      125215:data<=16'd6449;
      125216:data<=16'd6931;
      125217:data<=16'd5961;
      125218:data<=16'd5209;
      125219:data<=16'd6460;
      125220:data<=16'd3686;
      125221:data<=16'd6660;
      125222:data<=16'd18656;
      125223:data<=16'd22764;
      125224:data<=16'd20635;
      125225:data<=16'd21300;
      125226:data<=16'd20727;
      125227:data<=16'd20087;
      125228:data<=16'd20974;
      125229:data<=16'd19694;
      125230:data<=16'd17825;
      125231:data<=16'd17796;
      125232:data<=16'd18116;
      125233:data<=16'd17531;
      125234:data<=16'd17197;
      125235:data<=16'd17317;
      125236:data<=16'd16339;
      125237:data<=16'd15276;
      125238:data<=16'd14172;
      125239:data<=16'd12257;
      125240:data<=16'd12405;
      125241:data<=16'd13376;
      125242:data<=16'd11755;
      125243:data<=16'd10568;
      125244:data<=16'd11503;
      125245:data<=16'd12070;
      125246:data<=16'd11759;
      125247:data<=16'd11570;
      125248:data<=16'd11618;
      125249:data<=16'd10395;
      125250:data<=16'd8909;
      125251:data<=16'd9482;
      125252:data<=16'd6928;
      125253:data<=-16'd438;
      125254:data<=-16'd2511;
      125255:data<=16'd579;
      125256:data<=-16'd663;
      125257:data<=-16'd1615;
      125258:data<=16'd996;
      125259:data<=-16'd4538;
      125260:data<=-16'd16769;
      125261:data<=-16'd20240;
      125262:data<=-16'd16231;
      125263:data<=-16'd15567;
      125264:data<=-16'd16703;
      125265:data<=-16'd15547;
      125266:data<=-16'd14651;
      125267:data<=-16'd14408;
      125268:data<=-16'd13238;
      125269:data<=-16'd12975;
      125270:data<=-16'd13837;
      125271:data<=-16'd13396;
      125272:data<=-16'd12636;
      125273:data<=-16'd12883;
      125274:data<=-16'd12266;
      125275:data<=-16'd11320;
      125276:data<=-16'd11655;
      125277:data<=-16'd11188;
      125278:data<=-16'd9626;
      125279:data<=-16'd8939;
      125280:data<=-16'd8217;
      125281:data<=-16'd7400;
      125282:data<=-16'd7116;
      125283:data<=-16'd6161;
      125284:data<=-16'd6070;
      125285:data<=-16'd7266;
      125286:data<=-16'd7037;
      125287:data<=-16'd6253;
      125288:data<=-16'd5586;
      125289:data<=-16'd4825;
      125290:data<=-16'd5356;
      125291:data<=-16'd5335;
      125292:data<=-16'd4719;
      125293:data<=-16'd4313;
      125294:data<=-16'd2870;
      125295:data<=-16'd4068;
      125296:data<=-16'd1295;
      125297:data<=16'd14186;
      125298:data<=16'd24623;
      125299:data<=16'd21778;
      125300:data<=16'd21309;
      125301:data<=16'd21952;
      125302:data<=16'd19315;
      125303:data<=16'd19027;
      125304:data<=16'd18240;
      125305:data<=16'd17666;
      125306:data<=16'd18058;
      125307:data<=16'd15402;
      125308:data<=16'd15258;
      125309:data<=16'd16260;
      125310:data<=16'd13711;
      125311:data<=16'd14663;
      125312:data<=16'd16763;
      125313:data<=16'd14698;
      125314:data<=16'd13261;
      125315:data<=16'd12803;
      125316:data<=16'd12202;
      125317:data<=16'd11455;
      125318:data<=16'd10061;
      125319:data<=16'd9868;
      125320:data<=16'd8765;
      125321:data<=16'd7914;
      125322:data<=16'd9871;
      125323:data<=16'd8978;
      125324:data<=16'd7154;
      125325:data<=16'd7824;
      125326:data<=16'd6428;
      125327:data<=16'd5712;
      125328:data<=16'd6147;
      125329:data<=16'd5156;
      125330:data<=16'd6783;
      125331:data<=16'd6579;
      125332:data<=16'd4223;
      125333:data<=16'd6719;
      125334:data<=16'd2408;
      125335:data<=-16'd11432;
      125336:data<=-16'd15690;
      125337:data<=-16'd11961;
      125338:data<=-16'd13112;
      125339:data<=-16'd14016;
      125340:data<=-16'd11637;
      125341:data<=-16'd13235;
      125342:data<=-16'd18319;
      125343:data<=-16'd20669;
      125344:data<=-16'd19832;
      125345:data<=-16'd18336;
      125346:data<=-16'd17338;
      125347:data<=-16'd17065;
      125348:data<=-16'd16208;
      125349:data<=-16'd15575;
      125350:data<=-16'd16738;
      125351:data<=-16'd16269;
      125352:data<=-16'd13902;
      125353:data<=-16'd13655;
      125354:data<=-16'd13785;
      125355:data<=-16'd12742;
      125356:data<=-16'd12584;
      125357:data<=-16'd12498;
      125358:data<=-16'd11973;
      125359:data<=-16'd11614;
      125360:data<=-16'd10969;
      125361:data<=-16'd10578;
      125362:data<=-16'd10002;
      125363:data<=-16'd8705;
      125364:data<=-16'd7949;
      125365:data<=-16'd7591;
      125366:data<=-16'd7633;
      125367:data<=-16'd8516;
      125368:data<=-16'd8290;
      125369:data<=-16'd7906;
      125370:data<=-16'd9559;
      125371:data<=-16'd6196;
      125372:data<=16'd5773;
      125373:data<=16'd12980;
      125374:data<=16'd10160;
      125375:data<=16'd8928;
      125376:data<=16'd10328;
      125377:data<=16'd9204;
      125378:data<=16'd8880;
      125379:data<=16'd9385;
      125380:data<=16'd9376;
      125381:data<=16'd9473;
      125382:data<=16'd8448;
      125383:data<=16'd9057;
      125384:data<=16'd9406;
      125385:data<=16'd6866;
      125386:data<=16'd9931;
      125387:data<=16'd15547;
      125388:data<=16'd14531;
      125389:data<=16'd13209;
      125390:data<=16'd12971;
      125391:data<=16'd11041;
      125392:data<=16'd11215;
      125393:data<=16'd10800;
      125394:data<=16'd9759;
      125395:data<=16'd11232;
      125396:data<=16'd11341;
      125397:data<=16'd10790;
      125398:data<=16'd10466;
      125399:data<=16'd8661;
      125400:data<=16'd8020;
      125401:data<=16'd7392;
      125402:data<=16'd6526;
      125403:data<=16'd6498;
      125404:data<=16'd5130;
      125405:data<=16'd5247;
      125406:data<=16'd4996;
      125407:data<=16'd3566;
      125408:data<=16'd6736;
      125409:data<=16'd2804;
      125410:data<=-16'd10918;
      125411:data<=-16'd14684;
      125412:data<=-16'd12219;
      125413:data<=-16'd13873;
      125414:data<=-16'd13230;
      125415:data<=-16'd12455;
      125416:data<=-16'd12827;
      125417:data<=-16'd11559;
      125418:data<=-16'd12681;
      125419:data<=-16'd13083;
      125420:data<=-16'd11075;
      125421:data<=-16'd11324;
      125422:data<=-16'd12002;
      125423:data<=-16'd12070;
      125424:data<=-16'd12088;
      125425:data<=-16'd11414;
      125426:data<=-16'd11191;
      125427:data<=-16'd11119;
      125428:data<=-16'd11755;
      125429:data<=-16'd12237;
      125430:data<=-16'd12963;
      125431:data<=-16'd17834;
      125432:data<=-16'd20428;
      125433:data<=-16'd17660;
      125434:data<=-16'd17810;
      125435:data<=-16'd18339;
      125436:data<=-16'd16766;
      125437:data<=-16'd16904;
      125438:data<=-16'd15734;
      125439:data<=-16'd14499;
      125440:data<=-16'd14355;
      125441:data<=-16'd12924;
      125442:data<=-16'd14070;
      125443:data<=-16'd14266;
      125444:data<=-16'd11775;
      125445:data<=-16'd14008;
      125446:data<=-16'd12599;
      125447:data<=-16'd1909;
      125448:data<=16'd4643;
      125449:data<=16'd4640;
      125450:data<=16'd4692;
      125451:data<=16'd4202;
      125452:data<=16'd3589;
      125453:data<=16'd3720;
      125454:data<=16'd3237;
      125455:data<=16'd2936;
      125456:data<=16'd3137;
      125457:data<=16'd2702;
      125458:data<=16'd2397;
      125459:data<=16'd2933;
      125460:data<=16'd3166;
      125461:data<=16'd3049;
      125462:data<=16'd2560;
      125463:data<=16'd1368;
      125464:data<=16'd581;
      125465:data<=-16'd223;
      125466:data<=-16'd385;
      125467:data<=16'd978;
      125468:data<=16'd690;
      125469:data<=-16'd124;
      125470:data<=16'd67;
      125471:data<=-16'd984;
      125472:data<=-16'd91;
      125473:data<=16'd779;
      125474:data<=-16'd1507;
      125475:data<=16'd1207;
      125476:data<=16'd6781;
      125477:data<=16'd7424;
      125478:data<=16'd6384;
      125479:data<=16'd5063;
      125480:data<=16'd5156;
      125481:data<=16'd5855;
      125482:data<=16'd3665;
      125483:data<=16'd4441;
      125484:data<=16'd1474;
      125485:data<=-16'd11458;
      125486:data<=-16'd15653;
      125487:data<=-16'd11257;
      125488:data<=-16'd12551;
      125489:data<=-16'd12925;
      125490:data<=-16'd11590;
      125491:data<=-16'd12508;
      125492:data<=-16'd11082;
      125493:data<=-16'd10232;
      125494:data<=-16'd11044;
      125495:data<=-16'd10875;
      125496:data<=-16'd11317;
      125497:data<=-16'd10910;
      125498:data<=-16'd10393;
      125499:data<=-16'd10678;
      125500:data<=-16'd9653;
      125501:data<=-16'd9397;
      125502:data<=-16'd9461;
      125503:data<=-16'd8467;
      125504:data<=-16'd8237;
      125505:data<=-16'd8073;
      125506:data<=-16'd7990;
      125507:data<=-16'd7189;
      125508:data<=-16'd5530;
      125509:data<=-16'd5636;
      125510:data<=-16'd5118;
      125511:data<=-16'd4749;
      125512:data<=-16'd6913;
      125513:data<=-16'd6862;
      125514:data<=-16'd6015;
      125515:data<=-16'd6264;
      125516:data<=-16'd4916;
      125517:data<=-16'd5348;
      125518:data<=-16'd5424;
      125519:data<=-16'd4379;
      125520:data<=-16'd9298;
      125521:data<=-16'd10354;
      125522:data<=16'd203;
      125523:data<=16'd7647;
      125524:data<=16'd7295;
      125525:data<=16'd6992;
      125526:data<=16'd6956;
      125527:data<=16'd6555;
      125528:data<=16'd5952;
      125529:data<=16'd4325;
      125530:data<=16'd3830;
      125531:data<=16'd4030;
      125532:data<=16'd3259;
      125533:data<=16'd3976;
      125534:data<=16'd5460;
      125535:data<=16'd4761;
      125536:data<=16'd4106;
      125537:data<=16'd4607;
      125538:data<=16'd4438;
      125539:data<=16'd4056;
      125540:data<=16'd3680;
      125541:data<=16'd3618;
      125542:data<=16'd4108;
      125543:data<=16'd3924;
      125544:data<=16'd4018;
      125545:data<=16'd3535;
      125546:data<=16'd1413;
      125547:data<=16'd986;
      125548:data<=16'd1152;
      125549:data<=16'd740;
      125550:data<=16'd1902;
      125551:data<=16'd1917;
      125552:data<=16'd1322;
      125553:data<=16'd1309;
      125554:data<=16'd141;
      125555:data<=16'd1921;
      125556:data<=16'd2752;
      125557:data<=-16'd244;
      125558:data<=16'd1862;
      125559:data<=-16'd1083;
      125560:data<=-16'd14713;
      125561:data<=-16'd18396;
      125562:data<=-16'd15493;
      125563:data<=-16'd18553;
      125564:data<=-16'd15776;
      125565:data<=-16'd8539;
      125566:data<=-16'd6954;
      125567:data<=-16'd6234;
      125568:data<=-16'd5893;
      125569:data<=-16'd6915;
      125570:data<=-16'd5832;
      125571:data<=-16'd5065;
      125572:data<=-16'd5796;
      125573:data<=-16'd5695;
      125574:data<=-16'd4772;
      125575:data<=-16'd4358;
      125576:data<=-16'd5012;
      125577:data<=-16'd4604;
      125578:data<=-16'd3322;
      125579:data<=-16'd3980;
      125580:data<=-16'd4954;
      125581:data<=-16'd4637;
      125582:data<=-16'd3897;
      125583:data<=-16'd3040;
      125584:data<=-16'd3096;
      125585:data<=-16'd3115;
      125586:data<=-16'd2146;
      125587:data<=-16'd1812;
      125588:data<=-16'd1403;
      125589:data<=-16'd1154;
      125590:data<=-16'd1701;
      125591:data<=-16'd980;
      125592:data<=-16'd1265;
      125593:data<=-16'd2055;
      125594:data<=16'd170;
      125595:data<=-16'd626;
      125596:data<=-16'd1343;
      125597:data<=16'd8505;
      125598:data<=16'd17264;
      125599:data<=16'd16054;
      125600:data<=16'd15543;
      125601:data<=16'd15969;
      125602:data<=16'd14060;
      125603:data<=16'd13991;
      125604:data<=16'd13685;
      125605:data<=16'd12692;
      125606:data<=16'd12985;
      125607:data<=16'd13230;
      125608:data<=16'd13661;
      125609:data<=16'd10295;
      125610:data<=16'd4143;
      125611:data<=16'd3657;
      125612:data<=16'd4778;
      125613:data<=16'd3465;
      125614:data<=16'd3651;
      125615:data<=16'd3001;
      125616:data<=16'd2026;
      125617:data<=16'd2814;
      125618:data<=16'd2453;
      125619:data<=16'd2314;
      125620:data<=16'd2246;
      125621:data<=16'd1609;
      125622:data<=16'd2684;
      125623:data<=16'd2385;
      125624:data<=16'd1251;
      125625:data<=16'd1886;
      125626:data<=16'd1941;
      125627:data<=16'd2816;
      125628:data<=16'd2473;
      125629:data<=-16'd153;
      125630:data<=16'd1068;
      125631:data<=16'd1148;
      125632:data<=-16'd1328;
      125633:data<=16'd978;
      125634:data<=-16'd2388;
      125635:data<=-16'd14460;
      125636:data<=-16'd18463;
      125637:data<=-16'd15393;
      125638:data<=-16'd15030;
      125639:data<=-16'd14671;
      125640:data<=-16'd13640;
      125641:data<=-16'd13415;
      125642:data<=-16'd12170;
      125643:data<=-16'd11022;
      125644:data<=-16'd10997;
      125645:data<=-16'd11010;
      125646:data<=-16'd11418;
      125647:data<=-16'd11508;
      125648:data<=-16'd10455;
      125649:data<=-16'd10235;
      125650:data<=-16'd10103;
      125651:data<=-16'd8793;
      125652:data<=-16'd8655;
      125653:data<=-16'd6539;
      125654:data<=-16'd429;
      125655:data<=16'd1992;
      125656:data<=16'd977;
      125657:data<=16'd2359;
      125658:data<=16'd2758;
      125659:data<=16'd1547;
      125660:data<=16'd2029;
      125661:data<=16'd2322;
      125662:data<=16'd1762;
      125663:data<=16'd1063;
      125664:data<=16'd288;
      125665:data<=16'd886;
      125666:data<=16'd1759;
      125667:data<=16'd1134;
      125668:data<=16'd704;
      125669:data<=16'd1441;
      125670:data<=16'd1530;
      125671:data<=16'd3412;
      125672:data<=16'd11949;
      125673:data<=16'd20148;
      125674:data<=16'd20031;
      125675:data<=16'd18683;
      125676:data<=16'd19434;
      125677:data<=16'd18310;
      125678:data<=16'd17867;
      125679:data<=16'd17822;
      125680:data<=16'd16354;
      125681:data<=16'd16269;
      125682:data<=16'd16327;
      125683:data<=16'd15667;
      125684:data<=16'd15549;
      125685:data<=16'd14841;
      125686:data<=16'd14054;
      125687:data<=16'd13464;
      125688:data<=16'd13456;
      125689:data<=16'd14075;
      125690:data<=16'd12853;
      125691:data<=16'd11862;
      125692:data<=16'd11963;
      125693:data<=16'd10677;
      125694:data<=16'd10293;
      125695:data<=16'd10073;
      125696:data<=16'd10228;
      125697:data<=16'd12656;
      125698:data<=16'd9667;
      125699:data<=16'd2854;
      125700:data<=16'd1615;
      125701:data<=16'd2096;
      125702:data<=16'd2388;
      125703:data<=16'd3169;
      125704:data<=16'd1902;
      125705:data<=16'd2373;
      125706:data<=16'd2114;
      125707:data<=16'd244;
      125708:data<=16'd3113;
      125709:data<=-16'd517;
      125710:data<=-16'd13682;
      125711:data<=-16'd17496;
      125712:data<=-16'd13411;
      125713:data<=-16'd12555;
      125714:data<=-16'd11696;
      125715:data<=-16'd10695;
      125716:data<=-16'd10608;
      125717:data<=-16'd9235;
      125718:data<=-16'd8595;
      125719:data<=-16'd8990;
      125720:data<=-16'd9044;
      125721:data<=-16'd8977;
      125722:data<=-16'd8502;
      125723:data<=-16'd8126;
      125724:data<=-16'd8017;
      125725:data<=-16'd7744;
      125726:data<=-16'd7289;
      125727:data<=-16'd6461;
      125728:data<=-16'd5573;
      125729:data<=-16'd4303;
      125730:data<=-16'd3239;
      125731:data<=-16'd3312;
      125732:data<=-16'd2422;
      125733:data<=-16'd984;
      125734:data<=-16'd1239;
      125735:data<=-16'd1281;
      125736:data<=-16'd685;
      125737:data<=-16'd937;
      125738:data<=-16'd1169;
      125739:data<=-16'd1043;
      125740:data<=-16'd785;
      125741:data<=-16'd459;
      125742:data<=16'd770;
      125743:data<=16'd5109;
      125744:data<=16'd9301;
      125745:data<=16'd8429;
      125746:data<=16'd9171;
      125747:data<=16'd18668;
      125748:data<=16'd27473;
      125749:data<=16'd27023;
      125750:data<=16'd24876;
      125751:data<=16'd25170;
      125752:data<=16'd23896;
      125753:data<=16'd22953;
      125754:data<=16'd22633;
      125755:data<=16'd20384;
      125756:data<=16'd19276;
      125757:data<=16'd19023;
      125758:data<=16'd17779;
      125759:data<=16'd17922;
      125760:data<=16'd17455;
      125761:data<=16'd15535;
      125762:data<=16'd15844;
      125763:data<=16'd16783;
      125764:data<=16'd16099;
      125765:data<=16'd15453;
      125766:data<=16'd15245;
      125767:data<=16'd14442;
      125768:data<=16'd13167;
      125769:data<=16'd12900;
      125770:data<=16'd12847;
      125771:data<=16'd11541;
      125772:data<=16'd10598;
      125773:data<=16'd10040;
      125774:data<=16'd9643;
      125775:data<=16'd10014;
      125776:data<=16'd9368;
      125777:data<=16'd8599;
      125778:data<=16'd7987;
      125779:data<=16'd7109;
      125780:data<=16'd9007;
      125781:data<=16'd8931;
      125782:data<=16'd6355;
      125783:data<=16'd8625;
      125784:data<=16'd4172;
      125785:data<=-16'd9365;
      125786:data<=-16'd12219;
      125787:data<=-16'd11655;
      125788:data<=-16'd19364;
      125789:data<=-16'd21123;
      125790:data<=-16'd17731;
      125791:data<=-16'd18184;
      125792:data<=-16'd17223;
      125793:data<=-16'd15985;
      125794:data<=-16'd16339;
      125795:data<=-16'd15168;
      125796:data<=-16'd14387;
      125797:data<=-16'd13267;
      125798:data<=-16'd11811;
      125799:data<=-16'd12223;
      125800:data<=-16'd11456;
      125801:data<=-16'd10122;
      125802:data<=-16'd10305;
      125803:data<=-16'd9655;
      125804:data<=-16'd9053;
      125805:data<=-16'd9151;
      125806:data<=-16'd8313;
      125807:data<=-16'd7506;
      125808:data<=-16'd7479;
      125809:data<=-16'd7817;
      125810:data<=-16'd7749;
      125811:data<=-16'd7424;
      125812:data<=-16'd7457;
      125813:data<=-16'd5938;
      125814:data<=-16'd4288;
      125815:data<=-16'd4889;
      125816:data<=-16'd4519;
      125817:data<=-16'd3853;
      125818:data<=-16'd4244;
      125819:data<=-16'd2954;
      125820:data<=-16'd3460;
      125821:data<=-16'd3764;
      125822:data<=16'd4830;
      125823:data<=16'd14272;
      125824:data<=16'd14839;
      125825:data<=16'd13444;
      125826:data<=16'd13838;
      125827:data<=16'd12965;
      125828:data<=16'd12270;
      125829:data<=16'd12734;
      125830:data<=16'd12351;
      125831:data<=16'd11721;
      125832:data<=16'd14348;
      125833:data<=16'd18860;
      125834:data<=16'd19335;
      125835:data<=16'd17014;
      125836:data<=16'd16305;
      125837:data<=16'd15844;
      125838:data<=16'd15067;
      125839:data<=16'd14330;
      125840:data<=16'd12821;
      125841:data<=16'd12116;
      125842:data<=16'd11869;
      125843:data<=16'd11139;
      125844:data<=16'd10850;
      125845:data<=16'd9571;
      125846:data<=16'd8924;
      125847:data<=16'd10537;
      125848:data<=16'd10137;
      125849:data<=16'd8758;
      125850:data<=16'd8768;
      125851:data<=16'd7491;
      125852:data<=16'd7083;
      125853:data<=16'd7494;
      125854:data<=16'd5893;
      125855:data<=16'd5738;
      125856:data<=16'd5244;
      125857:data<=16'd3741;
      125858:data<=16'd5896;
      125859:data<=16'd1812;
      125860:data<=-16'd11065;
      125861:data<=-16'd15641;
      125862:data<=-16'd12895;
      125863:data<=-16'd12947;
      125864:data<=-16'd11870;
      125865:data<=-16'd10608;
      125866:data<=-16'd11317;
      125867:data<=-16'd10402;
      125868:data<=-16'd10363;
      125869:data<=-16'd10815;
      125870:data<=-16'd9441;
      125871:data<=-16'd9539;
      125872:data<=-16'd9941;
      125873:data<=-16'd9922;
      125874:data<=-16'd10473;
      125875:data<=-16'd9027;
      125876:data<=-16'd10349;
      125877:data<=-16'd16292;
      125878:data<=-16'd17875;
      125879:data<=-16'd15309;
      125880:data<=-16'd13706;
      125881:data<=-16'd12504;
      125882:data<=-16'd12358;
      125883:data<=-16'd12228;
      125884:data<=-16'd11203;
      125885:data<=-16'd10936;
      125886:data<=-16'd10198;
      125887:data<=-16'd9820;
      125888:data<=-16'd10346;
      125889:data<=-16'd9611;
      125890:data<=-16'd9222;
      125891:data<=-16'd8763;
      125892:data<=-16'd7805;
      125893:data<=-16'd8448;
      125894:data<=-16'd8037;
      125895:data<=-16'd8179;
      125896:data<=-16'd8349;
      125897:data<=16'd711;
      125898:data<=16'd11365;
      125899:data<=16'd11797;
      125900:data<=16'd10275;
      125901:data<=16'd10977;
      125902:data<=16'd10002;
      125903:data<=16'd9206;
      125904:data<=16'd8805;
      125905:data<=16'd8546;
      125906:data<=16'd8282;
      125907:data<=16'd6874;
      125908:data<=16'd6740;
      125909:data<=16'd7216;
      125910:data<=16'd6351;
      125911:data<=16'd5474;
      125912:data<=16'd4904;
      125913:data<=16'd6120;
      125914:data<=16'd7330;
      125915:data<=16'd6009;
      125916:data<=16'd6053;
      125917:data<=16'd6093;
      125918:data<=16'd4657;
      125919:data<=16'd5034;
      125920:data<=16'd4375;
      125921:data<=16'd5645;
      125922:data<=16'd11250;
      125923:data<=16'd11652;
      125924:data<=16'd9483;
      125925:data<=16'd10151;
      125926:data<=16'd8458;
      125927:data<=16'd7671;
      125928:data<=16'd8275;
      125929:data<=16'd6733;
      125930:data<=16'd7864;
      125931:data<=16'd7915;
      125932:data<=16'd6070;
      125933:data<=16'd8869;
      125934:data<=16'd4986;
      125935:data<=-16'd8022;
      125936:data<=-16'd12663;
      125937:data<=-16'd10693;
      125938:data<=-16'd11652;
      125939:data<=-16'd11119;
      125940:data<=-16'd9650;
      125941:data<=-16'd10863;
      125942:data<=-16'd11110;
      125943:data<=-16'd10295;
      125944:data<=-16'd10248;
      125945:data<=-16'd9136;
      125946:data<=-16'd8611;
      125947:data<=-16'd9727;
      125948:data<=-16'd9001;
      125949:data<=-16'd7709;
      125950:data<=-16'd8241;
      125951:data<=-16'd8487;
      125952:data<=-16'd8279;
      125953:data<=-16'd7932;
      125954:data<=-16'd7192;
      125955:data<=-16'd7197;
      125956:data<=-16'd7100;
      125957:data<=-16'd6745;
      125958:data<=-16'd6552;
      125959:data<=-16'd5877;
      125960:data<=-16'd5727;
      125961:data<=-16'd5127;
      125962:data<=-16'd4652;
      125963:data<=-16'd6310;
      125964:data<=-16'd6701;
      125965:data<=-16'd8081;
      125966:data<=-16'd13538;
      125967:data<=-16'd16178;
      125968:data<=-16'd15127;
      125969:data<=-16'd13900;
      125970:data<=-16'd13626;
      125971:data<=-16'd14624;
      125972:data<=-16'd7970;
      125973:data<=16'd4082;
      125974:data<=16'd6072;
      125975:data<=16'd3697;
      125976:data<=16'd5115;
      125977:data<=16'd4523;
      125978:data<=16'd3885;
      125979:data<=16'd4144;
      125980:data<=16'd2701;
      125981:data<=16'd2100;
      125982:data<=16'd1237;
      125983:data<=16'd611;
      125984:data<=16'd1134;
      125985:data<=16'd45;
      125986:data<=-16'd193;
      125987:data<=16'd681;
      125988:data<=16'd716;
      125989:data<=16'd1104;
      125990:data<=16'd318;
      125991:data<=16'd123;
      125992:data<=16'd1309;
      125993:data<=16'd296;
      125994:data<=-16'd229;
      125995:data<=16'd26;
      125996:data<=-16'd869;
      125997:data<=-16'd1146;
      125998:data<=-16'd2819;
      125999:data<=-16'd3704;
      126000:data<=-16'd2164;
      126001:data<=-16'd2784;
      126002:data<=-16'd2566;
      126003:data<=-16'd2079;
      126004:data<=-16'd3686;
      126005:data<=-16'd1762;
      126006:data<=-16'd1274;
      126007:data<=-16'd2852;
      126008:data<=-16'd170;
      126009:data<=-16'd5024;
      126010:data<=-16'd14698;
      126011:data<=-16'd12035;
      126012:data<=-16'd7955;
      126013:data<=-16'd11351;
      126014:data<=-16'd12037;
      126015:data<=-16'd10722;
      126016:data<=-16'd10681;
      126017:data<=-16'd9867;
      126018:data<=-16'd9730;
      126019:data<=-16'd9474;
      126020:data<=-16'd8240;
      126021:data<=-16'd8132;
      126022:data<=-16'd8960;
      126023:data<=-16'd9376;
      126024:data<=-16'd8658;
      126025:data<=-16'd7436;
      126026:data<=-16'd7112;
      126027:data<=-16'd7159;
      126028:data<=-16'd6487;
      126029:data<=-16'd5638;
      126030:data<=-16'd5908;
      126031:data<=-16'd6862;
      126032:data<=-16'd6710;
      126033:data<=-16'd5794;
      126034:data<=-16'd5389;
      126035:data<=-16'd5028;
      126036:data<=-16'd4397;
      126037:data<=-16'd4331;
      126038:data<=-16'd4420;
      126039:data<=-16'd3859;
      126040:data<=-16'd4003;
      126041:data<=-16'd4607;
      126042:data<=-16'd4570;
      126043:data<=-16'd5145;
      126044:data<=-16'd4144;
      126045:data<=-16'd2584;
      126046:data<=-16'd4646;
      126047:data<=-16'd446;
      126048:data<=16'd12000;
      126049:data<=16'd15371;
      126050:data<=16'd11712;
      126051:data<=16'd12225;
      126052:data<=16'd11676;
      126053:data<=16'd10774;
      126054:data<=16'd10598;
      126055:data<=16'd5074;
      126056:data<=16'd738;
      126057:data<=16'd1266;
      126058:data<=16'd854;
      126059:data<=16'd1017;
      126060:data<=16'd1572;
      126061:data<=16'd925;
      126062:data<=16'd1650;
      126063:data<=16'd1550;
      126064:data<=16'd14;
      126065:data<=-16'd335;
      126066:data<=-16'd600;
      126067:data<=-16'd617;
      126068:data<=-16'd174;
      126069:data<=-16'd767;
      126070:data<=-16'd1626;
      126071:data<=-16'd1530;
      126072:data<=-16'd669;
      126073:data<=-16'd872;
      126074:data<=-16'd2158;
      126075:data<=-16'd2137;
      126076:data<=-16'd1343;
      126077:data<=-16'd540;
      126078:data<=-16'd27;
      126079:data<=-16'd364;
      126080:data<=-16'd211;
      126081:data<=-16'd1767;
      126082:data<=-16'd3372;
      126083:data<=-16'd258;
      126084:data<=-16'd3139;
      126085:data<=-16'd15452;
      126086:data<=-16'd20562;
      126087:data<=-16'd17908;
      126088:data<=-16'd17459;
      126089:data<=-16'd17003;
      126090:data<=-16'd15908;
      126091:data<=-16'd15585;
      126092:data<=-16'd14565;
      126093:data<=-16'd13885;
      126094:data<=-16'd13509;
      126095:data<=-16'd12599;
      126096:data<=-16'd11094;
      126097:data<=-16'd11116;
      126098:data<=-16'd13820;
      126099:data<=-16'd11226;
      126100:data<=-16'd3377;
      126101:data<=-16'd1521;
      126102:data<=-16'd2608;
      126103:data<=-16'd1201;
      126104:data<=-16'd1574;
      126105:data<=-16'd1513;
      126106:data<=16'd118;
      126107:data<=16'd77;
      126108:data<=16'd378;
      126109:data<=16'd535;
      126110:data<=16'd85;
      126111:data<=16'd1401;
      126112:data<=16'd1859;
      126113:data<=16'd440;
      126114:data<=-16'd1017;
      126115:data<=-16'd2059;
      126116:data<=-16'd895;
      126117:data<=16'd38;
      126118:data<=-16'd1340;
      126119:data<=-16'd299;
      126120:data<=16'd287;
      126121:data<=-16'd2352;
      126122:data<=16'd3541;
      126123:data<=16'd16879;
      126124:data<=16'd20478;
      126125:data<=16'd17006;
      126126:data<=16'd17384;
      126127:data<=16'd16857;
      126128:data<=16'd14847;
      126129:data<=16'd15282;
      126130:data<=16'd13875;
      126131:data<=16'd11953;
      126132:data<=16'd12211;
      126133:data<=16'd10969;
      126134:data<=16'd10088;
      126135:data<=16'd10655;
      126136:data<=16'd10070;
      126137:data<=16'd10058;
      126138:data<=16'd9779;
      126139:data<=16'd8860;
      126140:data<=16'd9379;
      126141:data<=16'd8525;
      126142:data<=16'd7661;
      126143:data<=16'd8126;
      126144:data<=16'd3479;
      126145:data<=-16'd2796;
      126146:data<=-16'd2987;
      126147:data<=-16'd2473;
      126148:data<=-16'd4408;
      126149:data<=-16'd4247;
      126150:data<=-16'd3181;
      126151:data<=-16'd3380;
      126152:data<=-16'd2874;
      126153:data<=-16'd2752;
      126154:data<=-16'd3357;
      126155:data<=-16'd1932;
      126156:data<=-16'd1450;
      126157:data<=-16'd2303;
      126158:data<=16'd79;
      126159:data<=-16'd2640;
      126160:data<=-16'd14659;
      126161:data<=-16'd20506;
      126162:data<=-16'd17892;
      126163:data<=-16'd17935;
      126164:data<=-16'd18541;
      126165:data<=-16'd17503;
      126166:data<=-16'd17596;
      126167:data<=-16'd16539;
      126168:data<=-16'd15355;
      126169:data<=-16'd15405;
      126170:data<=-16'd13988;
      126171:data<=-16'd12583;
      126172:data<=-16'd12496;
      126173:data<=-16'd12016;
      126174:data<=-16'd11118;
      126175:data<=-16'd10185;
      126176:data<=-16'd9711;
      126177:data<=-16'd9160;
      126178:data<=-16'd7556;
      126179:data<=-16'd6540;
      126180:data<=-16'd6799;
      126181:data<=-16'd7535;
      126182:data<=-16'd7714;
      126183:data<=-16'd6399;
      126184:data<=-16'd6050;
      126185:data<=-16'd6278;
      126186:data<=-16'd4720;
      126187:data<=-16'd4787;
      126188:data<=-16'd3457;
      126189:data<=16'd3081;
      126190:data<=16'd5638;
      126191:data<=16'd3856;
      126192:data<=16'd4501;
      126193:data<=16'd4112;
      126194:data<=16'd4660;
      126195:data<=16'd6240;
      126196:data<=16'd3492;
      126197:data<=16'd7908;
      126198:data<=16'd20447;
      126199:data<=16'd22973;
      126200:data<=16'd19543;
      126201:data<=16'd20319;
      126202:data<=16'd19726;
      126203:data<=16'd18199;
      126204:data<=16'd18011;
      126205:data<=16'd17136;
      126206:data<=16'd17282;
      126207:data<=16'd17124;
      126208:data<=16'd15402;
      126209:data<=16'd14765;
      126210:data<=16'd14991;
      126211:data<=16'd14980;
      126212:data<=16'd14383;
      126213:data<=16'd13588;
      126214:data<=16'd13207;
      126215:data<=16'd12383;
      126216:data<=16'd12116;
      126217:data<=16'd12184;
      126218:data<=16'd11012;
      126219:data<=16'd10551;
      126220:data<=16'd10370;
      126221:data<=16'd9323;
      126222:data<=16'd9166;
      126223:data<=16'd9039;
      126224:data<=16'd8934;
      126225:data<=16'd9421;
      126226:data<=16'd9080;
      126227:data<=16'd9109;
      126228:data<=16'd9124;
      126229:data<=16'd8385;
      126230:data<=16'd8968;
      126231:data<=16'd9726;
      126232:data<=16'd10581;
      126233:data<=16'd9570;
      126234:data<=-16'd637;
      126235:data<=-16'd14223;
      126236:data<=-16'd18501;
      126237:data<=-16'd16832;
      126238:data<=-16'd16572;
      126239:data<=-16'd16051;
      126240:data<=-16'd14636;
      126241:data<=-16'd14286;
      126242:data<=-16'd14037;
      126243:data<=-16'd13333;
      126244:data<=-16'd12698;
      126245:data<=-16'd11374;
      126246:data<=-16'd10261;
      126247:data<=-16'd9518;
      126248:data<=-16'd7918;
      126249:data<=-16'd7509;
      126250:data<=-16'd7515;
      126251:data<=-16'd5877;
      126252:data<=-16'd5460;
      126253:data<=-16'd5582;
      126254:data<=-16'd5037;
      126255:data<=-16'd5438;
      126256:data<=-16'd4637;
      126257:data<=-16'd3744;
      126258:data<=-16'd4088;
      126259:data<=-16'd3034;
      126260:data<=-16'd2679;
      126261:data<=-16'd2666;
      126262:data<=-16'd1867;
      126263:data<=-16'd2648;
      126264:data<=-16'd1428;
      126265:data<=16'd698;
      126266:data<=16'd133;
      126267:data<=16'd168;
      126268:data<=-16'd757;
      126269:data<=-16'd531;
      126270:data<=16'd1562;
      126271:data<=-16'd1039;
      126272:data<=16'd3566;
      126273:data<=16'd17613;
      126274:data<=16'd20524;
      126275:data<=16'd16803;
      126276:data<=16'd17068;
      126277:data<=16'd17253;
      126278:data<=16'd21500;
      126279:data<=16'd25426;
      126280:data<=16'd22982;
      126281:data<=16'd23017;
      126282:data<=16'd23975;
      126283:data<=16'd22051;
      126284:data<=16'd21632;
      126285:data<=16'd21155;
      126286:data<=16'd20169;
      126287:data<=16'd19508;
      126288:data<=16'd18509;
      126289:data<=16'd18274;
      126290:data<=16'd17033;
      126291:data<=16'd16004;
      126292:data<=16'd16107;
      126293:data<=16'd14483;
      126294:data<=16'd13841;
      126295:data<=16'd13324;
      126296:data<=16'd11091;
      126297:data<=16'd11899;
      126298:data<=16'd13191;
      126299:data<=16'd12630;
      126300:data<=16'd12988;
      126301:data<=16'd12082;
      126302:data<=16'd11180;
      126303:data<=16'd11218;
      126304:data<=16'd9861;
      126305:data<=16'd9915;
      126306:data<=16'd9403;
      126307:data<=16'd7729;
      126308:data<=16'd9647;
      126309:data<=16'd6432;
      126310:data<=-16'd5935;
      126311:data<=-16'd12891;
      126312:data<=-16'd11546;
      126313:data<=-16'd11160;
      126314:data<=-16'd10906;
      126315:data<=-16'd8388;
      126316:data<=-16'd7656;
      126317:data<=-16'd8141;
      126318:data<=-16'd6922;
      126319:data<=-16'd6755;
      126320:data<=-16'd7153;
      126321:data<=-16'd5717;
      126322:data<=-16'd7911;
      126323:data<=-16'd14035;
      126324:data<=-16'd15863;
      126325:data<=-16'd13806;
      126326:data<=-16'd13100;
      126327:data<=-16'd13003;
      126328:data<=-16'd12759;
      126329:data<=-16'd13483;
      126330:data<=-16'd13292;
      126331:data<=-16'd10925;
      126332:data<=-16'd8909;
      126333:data<=-16'd8190;
      126334:data<=-16'd8035;
      126335:data<=-16'd8050;
      126336:data<=-16'd6860;
      126337:data<=-16'd6370;
      126338:data<=-16'd7699;
      126339:data<=-16'd7338;
      126340:data<=-16'd6699;
      126341:data<=-16'd6636;
      126342:data<=-16'd5542;
      126343:data<=-16'd6710;
      126344:data<=-16'd6708;
      126345:data<=-16'd4860;
      126346:data<=-16'd7756;
      126347:data<=-16'd3134;
      126348:data<=16'd12607;
      126349:data<=16'd17849;
      126350:data<=16'd14219;
      126351:data<=16'd14747;
      126352:data<=16'd13869;
      126353:data<=16'd12326;
      126354:data<=16'd12841;
      126355:data<=16'd11356;
      126356:data<=16'd11126;
      126357:data<=16'd11734;
      126358:data<=16'd10173;
      126359:data<=16'd9652;
      126360:data<=16'd9323;
      126361:data<=16'd8463;
      126362:data<=16'd8251;
      126363:data<=16'd7286;
      126364:data<=16'd7368;
      126365:data<=16'd8469;
      126366:data<=16'd9276;
      126367:data<=16'd12598;
      126368:data<=16'd16125;
      126369:data<=16'd15876;
      126370:data<=16'd14046;
      126371:data<=16'd13022;
      126372:data<=16'd12962;
      126373:data<=16'd12534;
      126374:data<=16'd11847;
      126375:data<=16'd12047;
      126376:data<=16'd11288;
      126377:data<=16'd10434;
      126378:data<=16'd10528;
      126379:data<=16'd9148;
      126380:data<=16'd8598;
      126381:data<=16'd9118;
      126382:data<=16'd8771;
      126383:data<=16'd10442;
      126384:data<=16'd7436;
      126385:data<=-16'd4507;
      126386:data<=-16'd11215;
      126387:data<=-16'd9700;
      126388:data<=-16'd9597;
      126389:data<=-16'd9699;
      126390:data<=-16'd8801;
      126391:data<=-16'd8758;
      126392:data<=-16'd8152;
      126393:data<=-16'd8499;
      126394:data<=-16'd9059;
      126395:data<=-16'd7667;
      126396:data<=-16'd7131;
      126397:data<=-16'd7410;
      126398:data<=-16'd6557;
      126399:data<=-16'd5497;
      126400:data<=-16'd4790;
      126401:data<=-16'd4858;
      126402:data<=-16'd5190;
      126403:data<=-16'd5103;
      126404:data<=-16'd5174;
      126405:data<=-16'd4760;
      126406:data<=-16'd4241;
      126407:data<=-16'd4156;
      126408:data<=-16'd3533;
      126409:data<=-16'd3136;
      126410:data<=-16'd2930;
      126411:data<=-16'd4670;
      126412:data<=-16'd10763;
      126413:data<=-16'd14117;
      126414:data<=-16'd11608;
      126415:data<=-16'd10360;
      126416:data<=-16'd9784;
      126417:data<=-16'd8790;
      126418:data<=-16'd9794;
      126419:data<=-16'd7649;
      126420:data<=-16'd5702;
      126421:data<=-16'd8934;
      126422:data<=-16'd3407;
      126423:data<=16'd10558;
      126424:data<=16'd14119;
      126425:data<=16'd11122;
      126426:data<=16'd11721;
      126427:data<=16'd10766;
      126428:data<=16'd9454;
      126429:data<=16'd9941;
      126430:data<=16'd8199;
      126431:data<=16'd8012;
      126432:data<=16'd9882;
      126433:data<=16'd8771;
      126434:data<=16'd7749;
      126435:data<=16'd7841;
      126436:data<=16'd6781;
      126437:data<=16'd6766;
      126438:data<=16'd6968;
      126439:data<=16'd6302;
      126440:data<=16'd6284;
      126441:data<=16'd5906;
      126442:data<=16'd5764;
      126443:data<=16'd5702;
      126444:data<=16'd3864;
      126445:data<=16'd3087;
      126446:data<=16'd3714;
      126447:data<=16'd3118;
      126448:data<=16'd3339;
      126449:data<=16'd4648;
      126450:data<=16'd4740;
      126451:data<=16'd4413;
      126452:data<=16'd4367;
      126453:data<=16'd3795;
      126454:data<=16'd2523;
      126455:data<=16'd2130;
      126456:data<=16'd4278;
      126457:data<=16'd8158;
      126458:data<=16'd11185;
      126459:data<=16'd7902;
      126460:data<=-16'd3121;
      126461:data<=-16'd11311;
      126462:data<=-16'd10994;
      126463:data<=-16'd9787;
      126464:data<=-16'd10066;
      126465:data<=-16'd8564;
      126466:data<=-16'd7153;
      126467:data<=-16'd7189;
      126468:data<=-16'd7236;
      126469:data<=-16'd7107;
      126470:data<=-16'd6980;
      126471:data<=-16'd6522;
      126472:data<=-16'd5846;
      126473:data<=-16'd6085;
      126474:data<=-16'd6851;
      126475:data<=-16'd6299;
      126476:data<=-16'd5712;
      126477:data<=-16'd6238;
      126478:data<=-16'd6273;
      126479:data<=-16'd5999;
      126480:data<=-16'd5570;
      126481:data<=-16'd4692;
      126482:data<=-16'd4740;
      126483:data<=-16'd5021;
      126484:data<=-16'd4737;
      126485:data<=-16'd4528;
      126486:data<=-16'd3993;
      126487:data<=-16'd4498;
      126488:data<=-16'd5426;
      126489:data<=-16'd4634;
      126490:data<=-16'd4696;
      126491:data<=-16'd4905;
      126492:data<=-16'd4196;
      126493:data<=-16'd5664;
      126494:data<=-16'd5219;
      126495:data<=-16'd3709;
      126496:data<=-16'd6346;
      126497:data<=-16'd1519;
      126498:data<=16'd11618;
      126499:data<=16'd14851;
      126500:data<=16'd9611;
      126501:data<=16'd6040;
      126502:data<=16'd3410;
      126503:data<=16'd2763;
      126504:data<=16'd2877;
      126505:data<=16'd1779;
      126506:data<=16'd1999;
      126507:data<=16'd1786;
      126508:data<=16'd704;
      126509:data<=16'd643;
      126510:data<=16'd617;
      126511:data<=16'd1165;
      126512:data<=16'd1042;
      126513:data<=16'd12;
      126514:data<=16'd267;
      126515:data<=-16'd1040;
      126516:data<=-16'd2807;
      126517:data<=-16'd1889;
      126518:data<=-16'd2223;
      126519:data<=-16'd3306;
      126520:data<=-16'd2946;
      126521:data<=-16'd3413;
      126522:data<=-16'd3560;
      126523:data<=-16'd3412;
      126524:data<=-16'd3874;
      126525:data<=-16'd3015;
      126526:data<=-16'd2563;
      126527:data<=-16'd3143;
      126528:data<=-16'd3063;
      126529:data<=-16'd3348;
      126530:data<=-16'd3134;
      126531:data<=-16'd3184;
      126532:data<=-16'd5153;
      126533:data<=-16'd5254;
      126534:data<=-16'd6778;
      126535:data<=-16'd16283;
      126536:data<=-16'd24256;
      126537:data<=-16'd22818;
      126538:data<=-16'd20996;
      126539:data<=-16'd21864;
      126540:data<=-16'd20415;
      126541:data<=-16'd19121;
      126542:data<=-16'd18788;
      126543:data<=-16'd17646;
      126544:data<=-16'd17734;
      126545:data<=-16'd15534;
      126546:data<=-16'd9661;
      126547:data<=-16'd7322;
      126548:data<=-16'd8654;
      126549:data<=-16'd9392;
      126550:data<=-16'd9427;
      126551:data<=-16'd9030;
      126552:data<=-16'd9135;
      126553:data<=-16'd8969;
      126554:data<=-16'd7929;
      126555:data<=-16'd8009;
      126556:data<=-16'd7867;
      126557:data<=-16'd7022;
      126558:data<=-16'd6795;
      126559:data<=-16'd6297;
      126560:data<=-16'd6252;
      126561:data<=-16'd5956;
      126562:data<=-16'd5347;
      126563:data<=-16'd6024;
      126564:data<=-16'd5453;
      126565:data<=-16'd5588;
      126566:data<=-16'd7420;
      126567:data<=-16'd6569;
      126568:data<=-16'd6743;
      126569:data<=-16'd6840;
      126570:data<=-16'd4581;
      126571:data<=-16'd6663;
      126572:data<=-16'd2534;
      126573:data<=16'd11762;
      126574:data<=16'd15437;
      126575:data<=16'd11347;
      126576:data<=16'd12405;
      126577:data<=16'd12266;
      126578:data<=16'd11408;
      126579:data<=16'd11694;
      126580:data<=16'd10082;
      126581:data<=16'd9659;
      126582:data<=16'd8595;
      126583:data<=16'd6296;
      126584:data<=16'd6194;
      126585:data<=16'd6044;
      126586:data<=16'd6153;
      126587:data<=16'd6413;
      126588:data<=16'd5483;
      126589:data<=16'd4787;
      126590:data<=16'd1439;
      126591:data<=-16'd2106;
      126592:data<=-16'd1703;
      126593:data<=-16'd2411;
      126594:data<=-16'd3015;
      126595:data<=-16'd1566;
      126596:data<=-16'd1768;
      126597:data<=-16'd1158;
      126598:data<=-16'd1213;
      126599:data<=-16'd3750;
      126600:data<=-16'd3190;
      126601:data<=-16'd2308;
      126602:data<=-16'd3785;
      126603:data<=-16'd3633;
      126604:data<=-16'd3280;
      126605:data<=-16'd2921;
      126606:data<=-16'd2159;
      126607:data<=-16'd2955;
      126608:data<=-16'd2297;
      126609:data<=-16'd3657;
      126610:data<=-16'd13041;
      126611:data<=-16'd21008;
      126612:data<=-16'd20668;
      126613:data<=-16'd19012;
      126614:data<=-16'd18697;
      126615:data<=-16'd18146;
      126616:data<=-16'd18750;
      126617:data<=-16'd18951;
      126618:data<=-16'd17801;
      126619:data<=-16'd17564;
      126620:data<=-16'd16753;
      126621:data<=-16'd14763;
      126622:data<=-16'd14369;
      126623:data<=-16'd14518;
      126624:data<=-16'd13656;
      126625:data<=-16'd12565;
      126626:data<=-16'd11574;
      126627:data<=-16'd11335;
      126628:data<=-16'd11097;
      126629:data<=-16'd10325;
      126630:data<=-16'd9841;
      126631:data<=-16'd8980;
      126632:data<=-16'd9406;
      126633:data<=-16'd11069;
      126634:data<=-16'd8698;
      126635:data<=-16'd3519;
      126636:data<=-16'd1154;
      126637:data<=-16'd1456;
      126638:data<=-16'd1512;
      126639:data<=-16'd713;
      126640:data<=-16'd1016;
      126641:data<=-16'd1196;
      126642:data<=-16'd237;
      126643:data<=-16'd1271;
      126644:data<=-16'd1025;
      126645:data<=16'd168;
      126646:data<=-16'd2438;
      126647:data<=16'd2975;
      126648:data<=16'd16688;
      126649:data<=16'd19023;
      126650:data<=16'd14489;
      126651:data<=16'd14895;
      126652:data<=16'd14616;
      126653:data<=16'd14169;
      126654:data<=16'd14683;
      126655:data<=16'd12956;
      126656:data<=16'd12689;
      126657:data<=16'd13306;
      126658:data<=16'd12693;
      126659:data<=16'd12610;
      126660:data<=16'd11621;
      126661:data<=16'd11041;
      126662:data<=16'd11605;
      126663:data<=16'd10968;
      126664:data<=16'd10901;
      126665:data<=16'd10314;
      126666:data<=16'd8282;
      126667:data<=16'd8026;
      126668:data<=16'd7353;
      126669:data<=16'd5753;
      126670:data<=16'd6147;
      126671:data<=16'd6490;
      126672:data<=16'd6302;
      126673:data<=16'd5988;
      126674:data<=16'd5115;
      126675:data<=16'd5858;
      126676:data<=16'd6106;
      126677:data<=16'd5039;
      126678:data<=16'd5507;
      126679:data<=16'd3142;
      126680:data<=-16'd1362;
      126681:data<=-16'd1530;
      126682:data<=-16'd1500;
      126683:data<=-16'd2754;
      126684:data<=-16'd4352;
      126685:data<=-16'd12933;
      126686:data<=-16'd21663;
      126687:data<=-16'd20606;
      126688:data<=-16'd18691;
      126689:data<=-16'd19256;
      126690:data<=-16'd17423;
      126691:data<=-16'd16433;
      126692:data<=-16'd16210;
      126693:data<=-16'd15173;
      126694:data<=-16'd15174;
      126695:data<=-16'd14038;
      126696:data<=-16'd12363;
      126697:data<=-16'd12219;
      126698:data<=-16'd12239;
      126699:data<=-16'd13069;
      126700:data<=-16'd13376;
      126701:data<=-16'd12408;
      126702:data<=-16'd12621;
      126703:data<=-16'd12173;
      126704:data<=-16'd10837;
      126705:data<=-16'd10270;
      126706:data<=-16'd9259;
      126707:data<=-16'd9342;
      126708:data<=-16'd9805;
      126709:data<=-16'd8510;
      126710:data<=-16'd7918;
      126711:data<=-16'd7517;
      126712:data<=-16'd6649;
      126713:data<=-16'd6252;
      126714:data<=-16'd5106;
      126715:data<=-16'd5485;
      126716:data<=-16'd6575;
      126717:data<=-16'd5512;
      126718:data<=-16'd5788;
      126719:data<=-16'd5570;
      126720:data<=-16'd4297;
      126721:data<=-16'd6475;
      126722:data<=-16'd2372;
      126723:data<=16'd11941;
      126724:data<=16'd20592;
      126725:data<=16'd20061;
      126726:data<=16'd19246;
      126727:data<=16'd19144;
      126728:data<=16'd18838;
      126729:data<=16'd18545;
      126730:data<=16'd17884;
      126731:data<=16'd17750;
      126732:data<=16'd17020;
      126733:data<=16'd14706;
      126734:data<=16'd13162;
      126735:data<=16'd13206;
      126736:data<=16'd13403;
      126737:data<=16'd13303;
      126738:data<=16'd12756;
      126739:data<=16'd12002;
      126740:data<=16'd11691;
      126741:data<=16'd11276;
      126742:data<=16'd10634;
      126743:data<=16'd10336;
      126744:data<=16'd10238;
      126745:data<=16'd10410;
      126746:data<=16'd10243;
      126747:data<=16'd9665;
      126748:data<=16'd9732;
      126749:data<=16'd9627;
      126750:data<=16'd9427;
      126751:data<=16'd9323;
      126752:data<=16'd8073;
      126753:data<=16'd7905;
      126754:data<=16'd8751;
      126755:data<=16'd8100;
      126756:data<=16'd7803;
      126757:data<=16'd7377;
      126758:data<=16'd7327;
      126759:data<=16'd7342;
      126760:data<=-16'd939;
      126761:data<=-16'd11667;
      126762:data<=-16'd12096;
      126763:data<=-16'd9765;
      126764:data<=-16'd10216;
      126765:data<=-16'd9130;
      126766:data<=-16'd7650;
      126767:data<=-16'd6044;
      126768:data<=-16'd7398;
      126769:data<=-16'd12495;
      126770:data<=-16'd12975;
      126771:data<=-16'd10818;
      126772:data<=-16'd11163;
      126773:data<=-16'd10775;
      126774:data<=-16'd10319;
      126775:data<=-16'd9903;
      126776:data<=-16'd8840;
      126777:data<=-16'd9019;
      126778:data<=-16'd8223;
      126779:data<=-16'd7142;
      126780:data<=-16'd7319;
      126781:data<=-16'd6586;
      126782:data<=-16'd6002;
      126783:data<=-16'd4701;
      126784:data<=-16'd2931;
      126785:data<=-16'd3633;
      126786:data<=-16'd3510;
      126787:data<=-16'd2739;
      126788:data<=-16'd3130;
      126789:data<=-16'd2176;
      126790:data<=-16'd2478;
      126791:data<=-16'd2641;
      126792:data<=-16'd484;
      126793:data<=-16'd1386;
      126794:data<=-16'd1908;
      126795:data<=-16'd1040;
      126796:data<=-16'd3657;
      126797:data<=16'd951;
      126798:data<=16'd13994;
      126799:data<=16'd19120;
      126800:data<=16'd17547;
      126801:data<=16'd18048;
      126802:data<=16'd18116;
      126803:data<=16'd16982;
      126804:data<=16'd16371;
      126805:data<=16'd15935;
      126806:data<=16'd15935;
      126807:data<=16'd15826;
      126808:data<=16'd15159;
      126809:data<=16'd14895;
      126810:data<=16'd14722;
      126811:data<=16'd13535;
      126812:data<=16'd13449;
      126813:data<=16'd16424;
      126814:data<=16'd18683;
      126815:data<=16'd18430;
      126816:data<=16'd18871;
      126817:data<=16'd19073;
      126818:data<=16'd17585;
      126819:data<=16'd17021;
      126820:data<=16'd16997;
      126821:data<=16'd16298;
      126822:data<=16'd16075;
      126823:data<=16'd15168;
      126824:data<=16'd13840;
      126825:data<=16'd14431;
      126826:data<=16'd14380;
      126827:data<=16'd12499;
      126828:data<=16'd12119;
      126829:data<=16'd12005;
      126830:data<=16'd11004;
      126831:data<=16'd11019;
      126832:data<=16'd10642;
      126833:data<=16'd11520;
      126834:data<=16'd12778;
      126835:data<=16'd5081;
      126836:data<=-16'd6222;
      126837:data<=-16'd8006;
      126838:data<=-16'd6038;
      126839:data<=-16'd6822;
      126840:data<=-16'd6369;
      126841:data<=-16'd5418;
      126842:data<=-16'd5623;
      126843:data<=-16'd5861;
      126844:data<=-16'd5812;
      126845:data<=-16'd4871;
      126846:data<=-16'd4660;
      126847:data<=-16'd5480;
      126848:data<=-16'd5040;
      126849:data<=-16'd3736;
      126850:data<=-16'd2279;
      126851:data<=-16'd1941;
      126852:data<=-16'd2875;
      126853:data<=-16'd2388;
      126854:data<=-16'd2147;
      126855:data<=-16'd2525;
      126856:data<=-16'd1321;
      126857:data<=-16'd3134;
      126858:data<=-16'd7846;
      126859:data<=-16'd9329;
      126860:data<=-16'd8924;
      126861:data<=-16'd8499;
      126862:data<=-16'd7774;
      126863:data<=-16'd7752;
      126864:data<=-16'd7444;
      126865:data<=-16'd7195;
      126866:data<=-16'd6360;
      126867:data<=-16'd4291;
      126868:data<=-16'd4205;
      126869:data<=-16'd3751;
      126870:data<=-16'd3112;
      126871:data<=-16'd6096;
      126872:data<=-16'd1900;
      126873:data<=16'd11215;
      126874:data<=16'd16066;
      126875:data<=16'd13482;
      126876:data<=16'd13496;
      126877:data<=16'd12950;
      126878:data<=16'd11740;
      126879:data<=16'd12017;
      126880:data<=16'd11195;
      126881:data<=16'd10320;
      126882:data<=16'd10715;
      126883:data<=16'd11157;
      126884:data<=16'd11141;
      126885:data<=16'd10728;
      126886:data<=16'd10487;
      126887:data<=16'd9793;
      126888:data<=16'd8901;
      126889:data<=16'd8918;
      126890:data<=16'd8508;
      126891:data<=16'd8108;
      126892:data<=16'd8217;
      126893:data<=16'd7459;
      126894:data<=16'd7350;
      126895:data<=16'd7423;
      126896:data<=16'd6657;
      126897:data<=16'd7286;
      126898:data<=16'd7353;
      126899:data<=16'd6631;
      126900:data<=16'd7694;
      126901:data<=16'd7629;
      126902:data<=16'd8878;
      126903:data<=16'd13743;
      126904:data<=16'd14041;
      126905:data<=16'd11406;
      126906:data<=16'd12179;
      126907:data<=16'd11427;
      126908:data<=16'd10426;
      126909:data<=16'd10897;
      126910:data<=16'd3620;
      126911:data<=-16'd7109;
      126912:data<=-16'd9459;
      126913:data<=-16'd8343;
      126914:data<=-16'd9329;
      126915:data<=-16'd9031;
      126916:data<=-16'd7474;
      126917:data<=-16'd6358;
      126918:data<=-16'd5985;
      126919:data<=-16'd6279;
      126920:data<=-16'd5826;
      126921:data<=-16'd5294;
      126922:data<=-16'd5351;
      126923:data<=-16'd4743;
      126924:data<=-16'd4440;
      126925:data<=-16'd4722;
      126926:data<=-16'd4510;
      126927:data<=-16'd4367;
      126928:data<=-16'd4194;
      126929:data<=-16'd4158;
      126930:data<=-16'd4034;
      126931:data<=-16'd3116;
      126932:data<=-16'd3256;
      126933:data<=-16'd3462;
      126934:data<=-16'd2265;
      126935:data<=-16'd2235;
      126936:data<=-16'd2176;
      126937:data<=-16'd1554;
      126938:data<=-16'd2326;
      126939:data<=-16'd2067;
      126940:data<=-16'd1962;
      126941:data<=-16'd2781;
      126942:data<=-16'd1416;
      126943:data<=-16'd1583;
      126944:data<=-16'd2184;
      126945:data<=-16'd905;
      126946:data<=-16'd4766;
      126947:data<=-16'd5656;
      126948:data<=16'd4479;
      126949:data<=16'd10351;
      126950:data<=16'd9407;
      126951:data<=16'd10768;
      126952:data<=16'd10113;
      126953:data<=16'd8768;
      126954:data<=16'd10408;
      126955:data<=16'd9583;
      126956:data<=16'd7817;
      126957:data<=16'd8002;
      126958:data<=16'd7473;
      126959:data<=16'd6639;
      126960:data<=16'd6056;
      126961:data<=16'd5827;
      126962:data<=16'd5796;
      126963:data<=16'd4636;
      126964:data<=16'd4335;
      126965:data<=16'd4752;
      126966:data<=16'd4105;
      126967:data<=16'd4725;
      126968:data<=16'd5303;
      126969:data<=16'd4511;
      126970:data<=16'd5300;
      126971:data<=16'd5674;
      126972:data<=16'd4423;
      126973:data<=16'd3950;
      126974:data<=16'd3472;
      126975:data<=16'd3351;
      126976:data<=16'd2949;
      126977:data<=16'd1568;
      126978:data<=16'd2547;
      126979:data<=16'd2655;
      126980:data<=16'd482;
      126981:data<=16'd1403;
      126982:data<=16'd1325;
      126983:data<=16'd914;
      126984:data<=16'd4458;
      126985:data<=-16'd922;
      126986:data<=-16'd13975;
      126987:data<=-16'd16674;
      126988:data<=-16'd13647;
      126989:data<=-16'd14257;
      126990:data<=-16'd14260;
      126991:data<=-16'd11908;
      126992:data<=-16'd7935;
      126993:data<=-16'd5846;
      126994:data<=-16'd6915;
      126995:data<=-16'd6102;
      126996:data<=-16'd5471;
      126997:data<=-16'd6416;
      126998:data<=-16'd5507;
      126999:data<=-16'd5333;
      127000:data<=-16'd4883;
      127001:data<=-16'd2808;
      127002:data<=-16'd3262;
      127003:data<=-16'd3703;
      127004:data<=-16'd2723;
      127005:data<=-16'd3137;
      127006:data<=-16'd3392;
      127007:data<=-16'd3759;
      127008:data<=-16'd4276;
      127009:data<=-16'd3920;
      127010:data<=-16'd4434;
      127011:data<=-16'd4391;
      127012:data<=-16'd3773;
      127013:data<=-16'd3976;
      127014:data<=-16'd3294;
      127015:data<=-16'd3747;
      127016:data<=-16'd4573;
      127017:data<=-16'd2972;
      127018:data<=-16'd2849;
      127019:data<=-16'd3106;
      127020:data<=-16'd2825;
      127021:data<=-16'd5438;
      127022:data<=-16'd1927;
      127023:data<=16'd9982;
      127024:data<=16'd14810;
      127025:data<=16'd12107;
      127026:data<=16'd11884;
      127027:data<=16'd11709;
      127028:data<=16'd10292;
      127029:data<=16'd10383;
      127030:data<=16'd9784;
      127031:data<=16'd9089;
      127032:data<=16'd9010;
      127033:data<=16'd6918;
      127034:data<=16'd5093;
      127035:data<=16'd3671;
      127036:data<=-16'd302;
      127037:data<=-16'd2954;
      127038:data<=-16'd3275;
      127039:data<=-16'd4065;
      127040:data<=-16'd3612;
      127041:data<=-16'd3162;
      127042:data<=-16'd3909;
      127043:data<=-16'd3812;
      127044:data<=-16'd4044;
      127045:data<=-16'd3630;
      127046:data<=-16'd2228;
      127047:data<=-16'd2508;
      127048:data<=-16'd2872;
      127049:data<=-16'd3530;
      127050:data<=-16'd4887;
      127051:data<=-16'd5048;
      127052:data<=-16'd6073;
      127053:data<=-16'd6476;
      127054:data<=-16'd5802;
      127055:data<=-16'd6990;
      127056:data<=-16'd6344;
      127057:data<=-16'd6035;
      127058:data<=-16'd7183;
      127059:data<=-16'd4306;
      127060:data<=-16'd8442;
      127061:data<=-16'd20927;
      127062:data<=-16'd23595;
      127063:data<=-16'd20885;
      127064:data<=-16'd21767;
      127065:data<=-16'd20383;
      127066:data<=-16'd19397;
      127067:data<=-16'd20651;
      127068:data<=-16'd20891;
      127069:data<=-16'd20991;
      127070:data<=-16'd19376;
      127071:data<=-16'd17546;
      127072:data<=-16'd17705;
      127073:data<=-16'd17167;
      127074:data<=-16'd16484;
      127075:data<=-16'd15913;
      127076:data<=-16'd15171;
      127077:data<=-16'd14929;
      127078:data<=-16'd13861;
      127079:data<=-16'd13364;
      127080:data<=-16'd11453;
      127081:data<=-16'd6344;
      127082:data<=-16'd4777;
      127083:data<=-16'd5990;
      127084:data<=-16'd5947;
      127085:data<=-16'd6837;
      127086:data<=-16'd6595;
      127087:data<=-16'd6108;
      127088:data<=-16'd7150;
      127089:data<=-16'd5805;
      127090:data<=-16'd5062;
      127091:data<=-16'd5783;
      127092:data<=-16'd4501;
      127093:data<=-16'd4461;
      127094:data<=-16'd3961;
      127095:data<=-16'd2848;
      127096:data<=-16'd5529;
      127097:data<=-16'd2438;
      127098:data<=16'd9295;
      127099:data<=16'd15057;
      127100:data<=16'd12871;
      127101:data<=16'd11113;
      127102:data<=16'd10593;
      127103:data<=16'd10202;
      127104:data<=16'd10055;
      127105:data<=16'd9497;
      127106:data<=16'd8793;
      127107:data<=16'd8573;
      127108:data<=16'd8478;
      127109:data<=16'd8226;
      127110:data<=16'd8075;
      127111:data<=16'd7600;
      127112:data<=16'd6981;
      127113:data<=16'd6721;
      127114:data<=16'd6232;
      127115:data<=16'd5915;
      127116:data<=16'd5404;
      127117:data<=16'd3852;
      127118:data<=16'd3175;
      127119:data<=16'd3330;
      127120:data<=16'd2801;
      127121:data<=16'd2773;
      127122:data<=16'd3178;
      127123:data<=16'd3081;
      127124:data<=16'd2090;
      127125:data<=-16'd984;
      127126:data<=-16'd4549;
      127127:data<=-16'd5333;
      127128:data<=-16'd3874;
      127129:data<=-16'd3683;
      127130:data<=-16'd4775;
      127131:data<=-16'd4196;
      127132:data<=-16'd3741;
      127133:data<=-16'd3692;
      127134:data<=-16'd2302;
      127135:data<=-16'd7385;
      127136:data<=-16'd18201;
      127137:data<=-16'd20742;
      127138:data<=-16'd17767;
      127139:data<=-16'd18089;
      127140:data<=-16'd17798;
      127141:data<=-16'd16665;
      127142:data<=-16'd16618;
      127143:data<=-16'd15946;
      127144:data<=-16'd15659;
      127145:data<=-16'd14762;
      127146:data<=-16'd13317;
      127147:data<=-16'd13317;
      127148:data<=-16'd12474;
      127149:data<=-16'd11433;
      127150:data<=-16'd11862;
      127151:data<=-16'd11699;
      127152:data<=-16'd11388;
      127153:data<=-16'd11320;
      127154:data<=-16'd11019;
      127155:data<=-16'd10800;
      127156:data<=-16'd9717;
      127157:data<=-16'd9165;
      127158:data<=-16'd9715;
      127159:data<=-16'd9424;
      127160:data<=-16'd8840;
      127161:data<=-16'd7955;
      127162:data<=-16'd7210;
      127163:data<=-16'd7139;
      127164:data<=-16'd6237;
      127165:data<=-16'd6255;
      127166:data<=-16'd6314;
      127167:data<=-16'd5278;
      127168:data<=-16'd6898;
      127169:data<=-16'd5459;
      127170:data<=16'd268;
      127171:data<=16'd290;
      127172:data<=16'd2478;
      127173:data<=16'd12704;
      127174:data<=16'd16920;
      127175:data<=16'd15209;
      127176:data<=16'd15543;
      127177:data<=16'd15003;
      127178:data<=16'd14166;
      127179:data<=16'd14405;
      127180:data<=16'd14242;
      127181:data<=16'd14295;
      127182:data<=16'd13397;
      127183:data<=16'd11929;
      127184:data<=16'd10960;
      127185:data<=16'd9717;
      127186:data<=16'd9391;
      127187:data<=16'd8962;
      127188:data<=16'd7832;
      127189:data<=16'd8147;
      127190:data<=16'd8332;
      127191:data<=16'd7940;
      127192:data<=16'd8102;
      127193:data<=16'd7503;
      127194:data<=16'd7090;
      127195:data<=16'd7448;
      127196:data<=16'd7550;
      127197:data<=16'd7576;
      127198:data<=16'd6924;
      127199:data<=16'd6592;
      127200:data<=16'd6631;
      127201:data<=16'd4673;
      127202:data<=16'd3374;
      127203:data<=16'd4400;
      127204:data<=16'd4099;
      127205:data<=16'd3122;
      127206:data<=16'd3530;
      127207:data<=16'd2954;
      127208:data<=16'd2391;
      127209:data<=16'd4173;
      127210:data<=16'd1093;
      127211:data<=-16'd9288;
      127212:data<=-16'd13279;
      127213:data<=-16'd9592;
      127214:data<=-16'd12017;
      127215:data<=-16'd16967;
      127216:data<=-16'd16327;
      127217:data<=-16'd16166;
      127218:data<=-16'd17444;
      127219:data<=-16'd16468;
      127220:data<=-16'd15333;
      127221:data<=-16'd14598;
      127222:data<=-16'd13641;
      127223:data<=-16'd12932;
      127224:data<=-16'd12128;
      127225:data<=-16'd11373;
      127226:data<=-16'd10743;
      127227:data<=-16'd10310;
      127228:data<=-16'd9922;
      127229:data<=-16'd9239;
      127230:data<=-16'd8809;
      127231:data<=-16'd8558;
      127232:data<=-16'd8445;
      127233:data<=-16'd8235;
      127234:data<=-16'd8009;
      127235:data<=-16'd9160;
      127236:data<=-16'd9606;
      127237:data<=-16'd8069;
      127238:data<=-16'd7444;
      127239:data<=-16'd6989;
      127240:data<=-16'd6278;
      127241:data<=-16'd6304;
      127242:data<=-16'd5166;
      127243:data<=-16'd4397;
      127244:data<=-16'd4282;
      127245:data<=-16'd3369;
      127246:data<=-16'd4200;
      127247:data<=-16'd1653;
      127248:data<=16'd7630;
      127249:data<=16'd12925;
      127250:data<=16'd11508;
      127251:data<=16'd10040;
      127252:data<=16'd9489;
      127253:data<=16'd9562;
      127254:data<=16'd9658;
      127255:data<=16'd9353;
      127256:data<=16'd9420;
      127257:data<=16'd8646;
      127258:data<=16'd9368;
      127259:data<=16'd13145;
      127260:data<=16'd15024;
      127261:data<=16'd14431;
      127262:data<=16'd14123;
      127263:data<=16'd13444;
      127264:data<=16'd12665;
      127265:data<=16'd12331;
      127266:data<=16'd11900;
      127267:data<=16'd11283;
      127268:data<=16'd10031;
      127269:data<=16'd8990;
      127270:data<=16'd9048;
      127271:data<=16'd9270;
      127272:data<=16'd9670;
      127273:data<=16'd9832;
      127274:data<=16'd8887;
      127275:data<=16'd8580;
      127276:data<=16'd9022;
      127277:data<=16'd8713;
      127278:data<=16'd8705;
      127279:data<=16'd8153;
      127280:data<=16'd6954;
      127281:data<=16'd7800;
      127282:data<=16'd7371;
      127283:data<=16'd5893;
      127284:data<=16'd8046;
      127285:data<=16'd4443;
      127286:data<=-16'd6925;
      127287:data<=-16'd10008;
      127288:data<=-16'd6619;
      127289:data<=-16'd7327;
      127290:data<=-16'd7473;
      127291:data<=-16'd6244;
      127292:data<=-16'd6590;
      127293:data<=-16'd6270;
      127294:data<=-16'd6109;
      127295:data<=-16'd5573;
      127296:data<=-16'd4150;
      127297:data<=-16'd4270;
      127298:data<=-16'd4152;
      127299:data<=-16'd3609;
      127300:data<=-16'd3604;
      127301:data<=-16'd1532;
      127302:data<=16'd382;
      127303:data<=-16'd1707;
      127304:data<=-16'd5477;
      127305:data<=-16'd6892;
      127306:data<=-16'd5912;
      127307:data<=-16'd5661;
      127308:data<=-16'd5705;
      127309:data<=-16'd4804;
      127310:data<=-16'd4672;
      127311:data<=-16'd4055;
      127312:data<=-16'd3297;
      127313:data<=-16'd4193;
      127314:data<=-16'd3644;
      127315:data<=-16'd2657;
      127316:data<=-16'd3163;
      127317:data<=-16'd1930;
      127318:data<=-16'd279;
      127319:data<=16'd705;
      127320:data<=16'd1747;
      127321:data<=16'd355;
      127322:data<=16'd2112;
      127323:data<=16'd11051;
      127324:data<=16'd16713;
      127325:data<=16'd15541;
      127326:data<=16'd14463;
      127327:data<=16'd14354;
      127328:data<=16'd14222;
      127329:data<=16'd14331;
      127330:data<=16'd13679;
      127331:data<=16'd13499;
      127332:data<=16'd13403;
      127333:data<=16'd11997;
      127334:data<=16'd12252;
      127335:data<=16'd13805;
      127336:data<=16'd13300;
      127337:data<=16'd12625;
      127338:data<=16'd12683;
      127339:data<=16'd12044;
      127340:data<=16'd11594;
      127341:data<=16'd10939;
      127342:data<=16'd10207;
      127343:data<=16'd10331;
      127344:data<=16'd10188;
      127345:data<=16'd9912;
      127346:data<=16'd8971;
      127347:data<=16'd8834;
      127348:data<=16'd12845;
      127349:data<=16'd15503;
      127350:data<=16'd14352;
      127351:data<=16'd15150;
      127352:data<=16'd15670;
      127353:data<=16'd14527;
      127354:data<=16'd14272;
      127355:data<=16'd12725;
      127356:data<=16'd12032;
      127357:data<=16'd12352;
      127358:data<=16'd11529;
      127359:data<=16'd12762;
      127360:data<=16'd8604;
      127361:data<=-16'd2848;
      127362:data<=-16'd6055;
      127363:data<=-16'd3109;
      127364:data<=-16'd3765;
      127365:data<=-16'd3720;
      127366:data<=-16'd3538;
      127367:data<=-16'd3936;
      127368:data<=-16'd2000;
      127369:data<=-16'd1486;
      127370:data<=-16'd1748;
      127371:data<=-16'd719;
      127372:data<=-16'd946;
      127373:data<=-16'd1121;
      127374:data<=-16'd864;
      127375:data<=-16'd996;
      127376:data<=-16'd696;
      127377:data<=-16'd1043;
      127378:data<=-16'd826;
      127379:data<=16'd44;
      127380:data<=-16'd584;
      127381:data<=-16'd529;
      127382:data<=-16'd176;
      127383:data<=-16'd1259;
      127384:data<=-16'd738;
      127385:data<=16'd869;
      127386:data<=16'd970;
      127387:data<=16'd911;
      127388:data<=16'd1169;
      127389:data<=16'd748;
      127390:data<=16'd729;
      127391:data<=16'd2030;
      127392:data<=16'd920;
      127393:data<=-16'd3888;
      127394:data<=-16'd5567;
      127395:data<=-16'd4232;
      127396:data<=-16'd5714;
      127397:data<=-16'd3617;
      127398:data<=16'd5827;
      127399:data<=16'd11718;
      127400:data<=16'd10696;
      127401:data<=16'd10103;
      127402:data<=16'd11013;
      127403:data<=16'd10869;
      127404:data<=16'd10439;
      127405:data<=16'd10252;
      127406:data<=16'd9829;
      127407:data<=16'd9209;
      127408:data<=16'd8642;
      127409:data<=16'd8587;
      127410:data<=16'd8373;
      127411:data<=16'd7426;
      127412:data<=16'd6974;
      127413:data<=16'd6717;
      127414:data<=16'd5979;
      127415:data<=16'd5705;
      127416:data<=16'd5383;
      127417:data<=16'd5301;
      127418:data<=16'd6256;
      127419:data<=16'd6727;
      127420:data<=16'd6928;
      127421:data<=16'd6877;
      127422:data<=16'd5855;
      127423:data<=16'd5771;
      127424:data<=16'd5641;
      127425:data<=16'd4651;
      127426:data<=16'd4816;
      127427:data<=16'd4449;
      127428:data<=16'd3993;
      127429:data<=16'd4340;
      127430:data<=16'd3099;
      127431:data<=16'd2960;
      127432:data<=16'd2968;
      127433:data<=16'd1463;
      127434:data<=16'd3785;
      127435:data<=16'd1268;
      127436:data<=-16'd10040;
      127437:data<=-16'd11033;
      127438:data<=-16'd3570;
      127439:data<=-16'd3585;
      127440:data<=-16'd4775;
      127441:data<=-16'd3714;
      127442:data<=-16'd5010;
      127443:data<=-16'd5236;
      127444:data<=-16'd5115;
      127445:data<=-16'd5545;
      127446:data<=-16'd4214;
      127447:data<=-16'd4026;
      127448:data<=-16'd4567;
      127449:data<=-16'd4087;
      127450:data<=-16'd4266;
      127451:data<=-16'd3560;
      127452:data<=-16'd2355;
      127453:data<=-16'd2560;
      127454:data<=-16'd2282;
      127455:data<=-16'd1844;
      127456:data<=-16'd2390;
      127457:data<=-16'd2817;
      127458:data<=-16'd2666;
      127459:data<=-16'd1868;
      127460:data<=-16'd1853;
      127461:data<=-16'd3045;
      127462:data<=-16'd3025;
      127463:data<=-16'd2322;
      127464:data<=-16'd2450;
      127465:data<=-16'd2397;
      127466:data<=-16'd2112;
      127467:data<=-16'd1883;
      127468:data<=-16'd1253;
      127469:data<=-16'd331;
      127470:data<=-16'd191;
      127471:data<=-16'd1557;
      127472:data<=16'd74;
      127473:data<=16'd8241;
      127474:data<=16'd14827;
      127475:data<=16'd13673;
      127476:data<=16'd11541;
      127477:data<=16'd11966;
      127478:data<=16'd11406;
      127479:data<=16'd10960;
      127480:data<=16'd11485;
      127481:data<=16'd9277;
      127482:data<=16'd5002;
      127483:data<=16'd2890;
      127484:data<=16'd3256;
      127485:data<=16'd3824;
      127486:data<=16'd3805;
      127487:data<=16'd3688;
      127488:data<=16'd3237;
      127489:data<=16'd2569;
      127490:data<=16'd2720;
      127491:data<=16'd2761;
      127492:data<=16'd1905;
      127493:data<=16'd1448;
      127494:data<=16'd1209;
      127495:data<=16'd807;
      127496:data<=16'd628;
      127497:data<=16'd284;
      127498:data<=16'd467;
      127499:data<=16'd734;
      127500:data<=16'd276;
      127501:data<=16'd954;
      127502:data<=16'd1571;
      127503:data<=16'd409;
      127504:data<=-16'd161;
      127505:data<=16'd171;
      127506:data<=16'd329;
      127507:data<=-16'd356;
      127508:data<=-16'd899;
      127509:data<=16'd752;
      127510:data<=-16'd3008;
      127511:data<=-16'd14210;
      127512:data<=-16'd17634;
      127513:data<=-16'd13890;
      127514:data<=-16'd14789;
      127515:data<=-16'd14901;
      127516:data<=-16'd12848;
      127517:data<=-16'd13772;
      127518:data<=-16'd13104;
      127519:data<=-16'd11414;
      127520:data<=-16'd11309;
      127521:data<=-16'd10464;
      127522:data<=-16'd10605;
      127523:data<=-16'd10616;
      127524:data<=-16'd9985;
      127525:data<=-16'd11057;
      127526:data<=-16'd8349;
      127527:data<=-16'd2881;
      127528:data<=-16'd2411;
      127529:data<=-16'd3366;
      127530:data<=-16'd2625;
      127531:data<=-16'd2784;
      127532:data<=-16'd2971;
      127533:data<=-16'd2996;
      127534:data<=-16'd2958;
      127535:data<=-16'd2023;
      127536:data<=-16'd1119;
      127537:data<=-16'd649;
      127538:data<=-16'd958;
      127539:data<=-16'd1416;
      127540:data<=-16'd1024;
      127541:data<=-16'd981;
      127542:data<=-16'd1019;
      127543:data<=-16'd949;
      127544:data<=-16'd1213;
      127545:data<=-16'd1028;
      127546:data<=-16'd1842;
      127547:data<=-16'd482;
      127548:data<=16'd7626;
      127549:data<=16'd14128;
      127550:data<=16'd13182;
      127551:data<=16'd11449;
      127552:data<=16'd11248;
      127553:data<=16'd10787;
      127554:data<=16'd10605;
      127555:data<=16'd10420;
      127556:data<=16'd10340;
      127557:data<=16'd9832;
      127558:data<=16'd8486;
      127559:data<=16'd8006;
      127560:data<=16'd7885;
      127561:data<=16'd7112;
      127562:data<=16'd6396;
      127563:data<=16'd5618;
      127564:data<=16'd5066;
      127565:data<=16'd4810;
      127566:data<=16'd4328;
      127567:data<=16'd3703;
      127568:data<=16'd2731;
      127569:data<=16'd2278;
      127570:data<=16'd1064;
      127571:data<=-16'd3407;
      127572:data<=-16'd6347;
      127573:data<=-16'd5200;
      127574:data<=-16'd5198;
      127575:data<=-16'd5668;
      127576:data<=-16'd4814;
      127577:data<=-16'd5554;
      127578:data<=-16'd5887;
      127579:data<=-16'd5057;
      127580:data<=-16'd5438;
      127581:data<=-16'd5362;
      127582:data<=-16'd5962;
      127583:data<=-16'd6504;
      127584:data<=-16'd4440;
      127585:data<=-16'd9007;
      127586:data<=-16'd20553;
      127587:data<=-16'd23971;
      127588:data<=-16'd20961;
      127589:data<=-16'd20841;
      127590:data<=-16'd20436;
      127591:data<=-16'd19610;
      127592:data<=-16'd20054;
      127593:data<=-16'd19165;
      127594:data<=-16'd18324;
      127595:data<=-16'd17963;
      127596:data<=-16'd17036;
      127597:data<=-16'd16615;
      127598:data<=-16'd15854;
      127599:data<=-16'd15382;
      127600:data<=-16'd15488;
      127601:data<=-16'd14616;
      127602:data<=-16'd14753;
      127603:data<=-16'd15129;
      127604:data<=-16'd14051;
      127605:data<=-16'd14026;
      127606:data<=-16'd13479;
      127607:data<=-16'd12260;
      127608:data<=-16'd13006;
      127609:data<=-16'd12430;
      127610:data<=-16'd11206;
      127611:data<=-16'd11671;
      127612:data<=-16'd10279;
      127613:data<=-16'd9527;
      127614:data<=-16'd10804;
      127615:data<=-16'd8128;
      127616:data<=-16'd3456;
      127617:data<=-16'd1760;
      127618:data<=-16'd2431;
      127619:data<=-16'd3930;
      127620:data<=-16'd4252;
      127621:data<=-16'd4334;
      127622:data<=-16'd3277;
      127623:data<=16'd3903;
      127624:data<=16'd11229;
      127625:data<=16'd11391;
      127626:data<=16'd10158;
      127627:data<=16'd10464;
      127628:data<=16'd9994;
      127629:data<=16'd9608;
      127630:data<=16'd9183;
      127631:data<=16'd9156;
      127632:data<=16'd9320;
      127633:data<=16'd8166;
      127634:data<=16'd7817;
      127635:data<=16'd7415;
      127636:data<=16'd5570;
      127637:data<=16'd5668;
      127638:data<=16'd5893;
      127639:data<=16'd4543;
      127640:data<=16'd4716;
      127641:data<=16'd4758;
      127642:data<=16'd4056;
      127643:data<=16'd4073;
      127644:data<=16'd3597;
      127645:data<=16'd3926;
      127646:data<=16'd4109;
      127647:data<=16'd2977;
      127648:data<=16'd3365;
      127649:data<=16'd2949;
      127650:data<=16'd1774;
      127651:data<=16'd2666;
      127652:data<=16'd1665;
      127653:data<=16'd303;
      127654:data<=16'd943;
      127655:data<=16'd267;
      127656:data<=16'd658;
      127657:data<=16'd628;
      127658:data<=-16'd406;
      127659:data<=16'd1836;
      127660:data<=-16'd4156;
      127661:data<=-16'd18877;
      127662:data<=-16'd22554;
      127663:data<=-16'd18989;
      127664:data<=-16'd19105;
      127665:data<=-16'd18142;
      127666:data<=-16'd17432;
      127667:data<=-16'd17461;
      127668:data<=-16'd16072;
      127669:data<=-16'd17130;
      127670:data<=-16'd17606;
      127671:data<=-16'd15802;
      127672:data<=-16'd15773;
      127673:data<=-16'd15338;
      127674:data<=-16'd14255;
      127675:data<=-16'd13949;
      127676:data<=-16'd12668;
      127677:data<=-16'd11708;
      127678:data<=-16'd11215;
      127679:data<=-16'd10763;
      127680:data<=-16'd10847;
      127681:data<=-16'd9345;
      127682:data<=-16'd8251;
      127683:data<=-16'd8804;
      127684:data<=-16'd7655;
      127685:data<=-16'd7768;
      127686:data<=-16'd10126;
      127687:data<=-16'd9486;
      127688:data<=-16'd7841;
      127689:data<=-16'd7926;
      127690:data<=-16'd7301;
      127691:data<=-16'd6537;
      127692:data<=-16'd6026;
      127693:data<=-16'd5213;
      127694:data<=-16'd5319;
      127695:data<=-16'd4824;
      127696:data<=-16'd4356;
      127697:data<=-16'd4167;
      127698:data<=16'd2848;
      127699:data<=16'd12422;
      127700:data<=16'd12894;
      127701:data<=16'd10784;
      127702:data<=16'd11371;
      127703:data<=16'd9135;
      127704:data<=16'd9691;
      127705:data<=16'd14875;
      127706:data<=16'd16057;
      127707:data<=16'd14947;
      127708:data<=16'd14959;
      127709:data<=16'd14522;
      127710:data<=16'd14132;
      127711:data<=16'd13232;
      127712:data<=16'd12583;
      127713:data<=16'd12480;
      127714:data<=16'd11652;
      127715:data<=16'd11923;
      127716:data<=16'd11964;
      127717:data<=16'd10954;
      127718:data<=16'd10862;
      127719:data<=16'd9643;
      127720:data<=16'd8693;
      127721:data<=16'd8969;
      127722:data<=16'd7961;
      127723:data<=16'd8420;
      127724:data<=16'd8539;
      127725:data<=16'd6828;
      127726:data<=16'd7891;
      127727:data<=16'd7765;
      127728:data<=16'd6006;
      127729:data<=16'd6843;
      127730:data<=16'd6643;
      127731:data<=16'd6956;
      127732:data<=16'd7212;
      127733:data<=16'd5359;
      127734:data<=16'd7476;
      127735:data<=16'd4115;
      127736:data<=-16'd8848;
      127737:data<=-16'd12613;
      127738:data<=-16'd9286;
      127739:data<=-16'd10032;
      127740:data<=-16'd9552;
      127741:data<=-16'd8892;
      127742:data<=-16'd9168;
      127743:data<=-16'd7935;
      127744:data<=-16'd8258;
      127745:data<=-16'd7794;
      127746:data<=-16'd6805;
      127747:data<=-16'd7216;
      127748:data<=-16'd5424;
      127749:data<=-16'd6843;
      127750:data<=-16'd12022;
      127751:data<=-16'd12003;
      127752:data<=-16'd10880;
      127753:data<=-16'd12094;
      127754:data<=-16'd11250;
      127755:data<=-16'd10105;
      127756:data<=-16'd9374;
      127757:data<=-16'd8533;
      127758:data<=-16'd8677;
      127759:data<=-16'd7873;
      127760:data<=-16'd7483;
      127761:data<=-16'd8066;
      127762:data<=-16'd6619;
      127763:data<=-16'd6040;
      127764:data<=-16'd6889;
      127765:data<=-16'd5491;
      127766:data<=-16'd4228;
      127767:data<=-16'd4181;
      127768:data<=-16'd4077;
      127769:data<=-16'd5054;
      127770:data<=-16'd4919;
      127771:data<=-16'd4259;
      127772:data<=-16'd4191;
      127773:data<=16'd2435;
      127774:data<=16'd11812;
      127775:data<=16'd12581;
      127776:data<=16'd10684;
      127777:data<=16'd11652;
      127778:data<=16'd10909;
      127779:data<=16'd10654;
      127780:data<=16'd11445;
      127781:data<=16'd10452;
      127782:data<=16'd10137;
      127783:data<=16'd10231;
      127784:data<=16'd10164;
      127785:data<=16'd10273;
      127786:data<=16'd8328;
      127787:data<=16'd7197;
      127788:data<=16'd7809;
      127789:data<=16'd6986;
      127790:data<=16'd7413;
      127791:data<=16'd8240;
      127792:data<=16'd6611;
      127793:data<=16'd7241;
      127794:data<=16'd10994;
      127795:data<=16'd13329;
      127796:data<=16'd13024;
      127797:data<=16'd12063;
      127798:data<=16'd11966;
      127799:data<=16'd11248;
      127800:data<=16'd10677;
      127801:data<=16'd11141;
      127802:data<=16'd9530;
      127803:data<=16'd8023;
      127804:data<=16'd8367;
      127805:data<=16'd7620;
      127806:data<=16'd7806;
      127807:data<=16'd8012;
      127808:data<=16'd7307;
      127809:data<=16'd9166;
      127810:data<=16'd5251;
      127811:data<=-16'd6097;
      127812:data<=-16'd9582;
      127813:data<=-16'd6605;
      127814:data<=-16'd6913;
      127815:data<=-16'd7021;
      127816:data<=-16'd6743;
      127817:data<=-16'd7538;
      127818:data<=-16'd6222;
      127819:data<=-16'd5189;
      127820:data<=-16'd5645;
      127821:data<=-16'd5127;
      127822:data<=-16'd4673;
      127823:data<=-16'd4266;
      127824:data<=-16'd3548;
      127825:data<=-16'd3636;
      127826:data<=-16'd3445;
      127827:data<=-16'd3055;
      127828:data<=-16'd2995;
      127829:data<=-16'd2372;
      127830:data<=-16'd2174;
      127831:data<=-16'd2082;
      127832:data<=-16'd1428;
      127833:data<=-16'd1333;
      127834:data<=-16'd698;
      127835:data<=-16'd315;
      127836:data<=-16'd185;
      127837:data<=16'd2358;
      127838:data<=16'd1340;
      127839:data<=-16'd4270;
      127840:data<=-16'd4775;
      127841:data<=-16'd3268;
      127842:data<=-16'd4356;
      127843:data<=-16'd3459;
      127844:data<=-16'd2981;
      127845:data<=-16'd2955;
      127846:data<=-16'd1935;
      127847:data<=-16'd2752;
      127848:data<=16'd2734;
      127849:data<=16'd13229;
      127850:data<=16'd14310;
      127851:data<=16'd11687;
      127852:data<=16'd13200;
      127853:data<=16'd13644;
      127854:data<=16'd13806;
      127855:data<=16'd14111;
      127856:data<=16'd13306;
      127857:data<=16'd13427;
      127858:data<=16'd12865;
      127859:data<=16'd12279;
      127860:data<=16'd12595;
      127861:data<=16'd11755;
      127862:data<=16'd11462;
      127863:data<=16'd11283;
      127864:data<=16'd10410;
      127865:data<=16'd10710;
      127866:data<=16'd10433;
      127867:data<=16'd9667;
      127868:data<=16'd9465;
      127869:data<=16'd9189;
      127870:data<=16'd10249;
      127871:data<=16'd10608;
      127872:data<=16'd9585;
      127873:data<=16'd9674;
      127874:data<=16'd8851;
      127875:data<=16'd8229;
      127876:data<=16'd8934;
      127877:data<=16'd7858;
      127878:data<=16'd7177;
      127879:data<=16'd7165;
      127880:data<=16'd6531;
      127881:data<=16'd7210;
      127882:data<=16'd6807;
      127883:data<=16'd8617;
      127884:data<=16'd14320;
      127885:data<=16'd10710;
      127886:data<=-16'd241;
      127887:data<=-16'd3095;
      127888:data<=-16'd1221;
      127889:data<=-16'd1676;
      127890:data<=-16'd1895;
      127891:data<=-16'd2043;
      127892:data<=-16'd2391;
      127893:data<=-16'd1889;
      127894:data<=-16'd1703;
      127895:data<=-16'd1670;
      127896:data<=-16'd1679;
      127897:data<=-16'd2218;
      127898:data<=-16'd2087;
      127899:data<=-16'd1541;
      127900:data<=-16'd1522;
      127901:data<=-16'd1058;
      127902:data<=-16'd520;
      127903:data<=-16'd297;
      127904:data<=16'd573;
      127905:data<=16'd772;
      127906:data<=16'd381;
      127907:data<=16'd811;
      127908:data<=16'd429;
      127909:data<=16'd24;
      127910:data<=16'd503;
      127911:data<=16'd9;
      127912:data<=16'd173;
      127913:data<=16'd729;
      127914:data<=16'd446;
      127915:data<=16'd1339;
      127916:data<=16'd1049;
      127917:data<=-16'd29;
      127918:data<=16'd481;
      127919:data<=-16'd59;
      127920:data<=16'd1709;
      127921:data<=16'd3312;
      127922:data<=16'd102;
      127923:data<=16'd5721;
      127924:data<=16'd17068;
      127925:data<=16'd17182;
      127926:data<=16'd15158;
      127927:data<=16'd14418;
      127928:data<=16'd8158;
      127929:data<=16'd6302;
      127930:data<=16'd8184;
      127931:data<=16'd6572;
      127932:data<=16'd6437;
      127933:data<=16'd6617;
      127934:data<=16'd5940;
      127935:data<=16'd6502;
      127936:data<=16'd6179;
      127937:data<=16'd7040;
      127938:data<=16'd7661;
      127939:data<=16'd5981;
      127940:data<=16'd6341;
      127941:data<=16'd6250;
      127942:data<=16'd4730;
      127943:data<=16'd5137;
      127944:data<=16'd4833;
      127945:data<=16'd4096;
      127946:data<=16'd3650;
      127947:data<=16'd2914;
      127948:data<=16'd3923;
      127949:data<=16'd3554;
      127950:data<=16'd2311;
      127951:data<=16'd3018;
      127952:data<=16'd2121;
      127953:data<=16'd2670;
      127954:data<=16'd4725;
      127955:data<=16'd3227;
      127956:data<=16'd3459;
      127957:data<=16'd4034;
      127958:data<=16'd2432;
      127959:data<=16'd4708;
      127960:data<=16'd1662;
      127961:data<=-16'd9978;
      127962:data<=-16'd14377;
      127963:data<=-16'd12439;
      127964:data<=-16'd12706;
      127965:data<=-16'd12730;
      127966:data<=-16'd12307;
      127967:data<=-16'd12093;
      127968:data<=-16'd11644;
      127969:data<=-16'd10957;
      127970:data<=-16'd9562;
      127971:data<=-16'd9353;
      127972:data<=-16'd7218;
      127973:data<=-16'd1774;
      127974:data<=-16'd717;
      127975:data<=-16'd2177;
      127976:data<=-16'd820;
      127977:data<=-16'd989;
      127978:data<=-16'd2076;
      127979:data<=-16'd1873;
      127980:data<=-16'd2896;
      127981:data<=-16'd2834;
      127982:data<=-16'd1357;
      127983:data<=-16'd1521;
      127984:data<=-16'd1735;
      127985:data<=-16'd1770;
      127986:data<=-16'd1623;
      127987:data<=16'd226;
      127988:data<=16'd557;
      127989:data<=-16'd581;
      127990:data<=16'd256;
      127991:data<=16'd162;
      127992:data<=-16'd1031;
      127993:data<=-16'd960;
      127994:data<=-16'd1817;
      127995:data<=-16'd1387;
      127996:data<=-16'd607;
      127997:data<=-16'd3271;
      127998:data<=16'd983;
      127999:data<=16'd12251;
      128000:data<=16'd14571;
      128001:data<=16'd11823;
      128002:data<=16'd12542;
      128003:data<=16'd12111;
      128004:data<=16'd12161;
      128005:data<=16'd13009;
      128006:data<=16'd11632;
      128007:data<=16'd11126;
      128008:data<=16'd10302;
      128009:data<=16'd9276;
      128010:data<=16'd10040;
      128011:data<=16'd8927;
      128012:data<=16'd7811;
      128013:data<=16'd7655;
      128014:data<=16'd6108;
      128015:data<=16'd6702;
      128016:data<=16'd5888;
      128017:data<=16'd540;
      128018:data<=-16'd1932;
      128019:data<=-16'd1137;
      128020:data<=-16'd370;
      128021:data<=16'd194;
      128022:data<=-16'd440;
      128023:data<=-16'd705;
      128024:data<=-16'd893;
      128025:data<=-16'd1007;
      128026:data<=-16'd88;
      128027:data<=-16'd1380;
      128028:data<=-16'd2217;
      128029:data<=-16'd1202;
      128030:data<=-16'd2240;
      128031:data<=-16'd1698;
      128032:data<=-16'd1444;
      128033:data<=-16'd3253;
      128034:data<=-16'd817;
      128035:data<=-16'd3518;
      128036:data<=-16'd14402;
      128037:data<=-16'd17233;
      128038:data<=-16'd14384;
      128039:data<=-16'd14775;
      128040:data<=-16'd14639;
      128041:data<=-16'd14552;
      128042:data<=-16'd14697;
      128043:data<=-16'd13750;
      128044:data<=-16'd13916;
      128045:data<=-16'd13494;
      128046:data<=-16'd12790;
      128047:data<=-16'd13274;
      128048:data<=-16'd12434;
      128049:data<=-16'd11251;
      128050:data<=-16'd11188;
      128051:data<=-16'd11247;
      128052:data<=-16'd11116;
      128053:data<=-16'd10008;
      128054:data<=-16'd8915;
      128055:data<=-16'd8757;
      128056:data<=-16'd8373;
      128057:data<=-16'd7944;
      128058:data<=-16'd7298;
      128059:data<=-16'd7156;
      128060:data<=-16'd8120;
      128061:data<=-16'd5671;
      128062:data<=-16'd146;
      128063:data<=16'd1122;
      128064:data<=-16'd513;
      128065:data<=-16'd114;
      128066:data<=-16'd503;
      128067:data<=-16'd1459;
      128068:data<=-16'd876;
      128069:data<=-16'd1512;
      128070:data<=-16'd649;
      128071:data<=16'd1075;
      128072:data<=-16'd1224;
      128073:data<=16'd3140;
      128074:data<=16'd14713;
      128075:data<=16'd16110;
      128076:data<=16'd12404;
      128077:data<=16'd13424;
      128078:data<=16'd12455;
      128079:data<=16'd11512;
      128080:data<=16'd12489;
      128081:data<=16'd11151;
      128082:data<=16'd10522;
      128083:data<=16'd10040;
      128084:data<=16'd8796;
      128085:data<=16'd8895;
      128086:data<=16'd7776;
      128087:data<=16'd6971;
      128088:data<=16'd7034;
      128089:data<=16'd5562;
      128090:data<=16'd5647;
      128091:data<=16'd6029;
      128092:data<=16'd5090;
      128093:data<=16'd5174;
      128094:data<=16'd4240;
      128095:data<=16'd3290;
      128096:data<=16'd3483;
      128097:data<=16'd2767;
      128098:data<=16'd2875;
      128099:data<=16'd2344;
      128100:data<=16'd1001;
      128101:data<=16'd1715;
      128102:data<=16'd998;
      128103:data<=-16'd443;
      128104:data<=-16'd276;
      128105:data<=-16'd2041;
      128106:data<=-16'd5059;
      128107:data<=-16'd8194;
      128108:data<=-16'd9256;
      128109:data<=-16'd6446;
      128110:data<=-16'd9427;
      128111:data<=-16'd19226;
      128112:data<=-16'd23347;
      128113:data<=-16'd21716;
      128114:data<=-16'd20829;
      128115:data<=-16'd20624;
      128116:data<=-16'd20422;
      128117:data<=-16'd20169;
      128118:data<=-16'd19875;
      128119:data<=-16'd19650;
      128120:data<=-16'd19331;
      128121:data<=-16'd19164;
      128122:data<=-16'd18870;
      128123:data<=-16'd18131;
      128124:data<=-16'd17235;
      128125:data<=-16'd16847;
      128126:data<=-16'd16446;
      128127:data<=-16'd15250;
      128128:data<=-16'd14797;
      128129:data<=-16'd14663;
      128130:data<=-16'd13747;
      128131:data<=-16'd13353;
      128132:data<=-16'd12436;
      128133:data<=-16'd11605;
      128134:data<=-16'd12151;
      128135:data<=-16'd11555;
      128136:data<=-16'd11156;
      128137:data<=-16'd11891;
      128138:data<=-16'd11724;
      128139:data<=-16'd11638;
      128140:data<=-16'd10701;
      128141:data<=-16'd9690;
      128142:data<=-16'd10301;
      128143:data<=-16'd10016;
      128144:data<=-16'd10053;
      128145:data<=-16'd9327;
      128146:data<=-16'd7877;
      128147:data<=-16'd9903;
      128148:data<=-16'd5556;
      128149:data<=16'd5943;
      128150:data<=16'd9988;
      128151:data<=16'd11782;
      128152:data<=16'd14918;
      128153:data<=16'd12305;
      128154:data<=16'd10655;
      128155:data<=16'd10928;
      128156:data<=16'd9327;
      128157:data<=16'd9887;
      128158:data<=16'd9950;
      128159:data<=16'd9097;
      128160:data<=16'd9356;
      128161:data<=16'd8251;
      128162:data<=16'd8436;
      128163:data<=16'd8746;
      128164:data<=16'd7098;
      128165:data<=16'd7166;
      128166:data<=16'd6951;
      128167:data<=16'd6231;
      128168:data<=16'd6540;
      128169:data<=16'd5711;
      128170:data<=16'd5165;
      128171:data<=16'd3641;
      128172:data<=16'd1589;
      128173:data<=16'd2497;
      128174:data<=16'd2206;
      128175:data<=16'd1588;
      128176:data<=16'd2661;
      128177:data<=16'd1454;
      128178:data<=16'd1756;
      128179:data<=16'd3218;
      128180:data<=16'd1847;
      128181:data<=16'd2191;
      128182:data<=16'd2268;
      128183:data<=16'd1183;
      128184:data<=16'd3284;
      128185:data<=16'd682;
      128186:data<=-16'd9295;
      128187:data<=-16'd15380;
      128188:data<=-16'd14935;
      128189:data<=-16'd14046;
      128190:data<=-16'd14170;
      128191:data<=-16'd13412;
      128192:data<=-16'd12869;
      128193:data<=-16'd12646;
      128194:data<=-16'd11674;
      128195:data<=-16'd13612;
      128196:data<=-16'd17111;
      128197:data<=-16'd17030;
      128198:data<=-16'd16107;
      128199:data<=-16'd15684;
      128200:data<=-16'd14800;
      128201:data<=-16'd14572;
      128202:data<=-16'd13350;
      128203:data<=-16'd12578;
      128204:data<=-16'd13794;
      128205:data<=-16'd13954;
      128206:data<=-16'd13424;
      128207:data<=-16'd12665;
      128208:data<=-16'd11298;
      128209:data<=-16'd10575;
      128210:data<=-16'd9905;
      128211:data<=-16'd9538;
      128212:data<=-16'd8828;
      128213:data<=-16'd7503;
      128214:data<=-16'd7550;
      128215:data<=-16'd6981;
      128216:data<=-16'd6222;
      128217:data<=-16'd6733;
      128218:data<=-16'd6049;
      128219:data<=-16'd6026;
      128220:data<=-16'd5685;
      128221:data<=-16'd5187;
      128222:data<=-16'd8348;
      128223:data<=-16'd3976;
      128224:data<=16'd8464;
      128225:data<=16'd11079;
      128226:data<=16'd8451;
      128227:data<=16'd9940;
      128228:data<=16'd9524;
      128229:data<=16'd8715;
      128230:data<=16'd9564;
      128231:data<=16'd9477;
      128232:data<=16'd9389;
      128233:data<=16'd8809;
      128234:data<=16'd8602;
      128235:data<=16'd8837;
      128236:data<=16'd8214;
      128237:data<=16'd7871;
      128238:data<=16'd5955;
      128239:data<=16'd5603;
      128240:data<=16'd10451;
      128241:data<=16'd12645;
      128242:data<=16'd11135;
      128243:data<=16'd11233;
      128244:data<=16'd11056;
      128245:data<=16'd10586;
      128246:data<=16'd10539;
      128247:data<=16'd9993;
      128248:data<=16'd9817;
      128249:data<=16'd9213;
      128250:data<=16'd8986;
      128251:data<=16'd9148;
      128252:data<=16'd8050;
      128253:data<=16'd7991;
      128254:data<=16'd7623;
      128255:data<=16'd5794;
      128256:data<=16'd6182;
      128257:data<=16'd6009;
      128258:data<=16'd4814;
      128259:data<=16'd6590;
      128260:data<=16'd4394;
      128261:data<=-16'd5104;
      128262:data<=-16'd11079;
      128263:data<=-16'd10094;
      128264:data<=-16'd9206;
      128265:data<=-16'd9371;
      128266:data<=-16'd8314;
      128267:data<=-16'd8200;
      128268:data<=-16'd8504;
      128269:data<=-16'd7347;
      128270:data<=-16'd7283;
      128271:data<=-16'd8317;
      128272:data<=-16'd8607;
      128273:data<=-16'd8393;
      128274:data<=-16'd7291;
      128275:data<=-16'd6974;
      128276:data<=-16'd7441;
      128277:data<=-16'd6078;
      128278:data<=-16'd5389;
      128279:data<=-16'd5767;
      128280:data<=-16'd4831;
      128281:data<=-16'd4786;
      128282:data<=-16'd4457;
      128283:data<=-16'd2763;
      128284:data<=-16'd4555;
      128285:data<=-16'd8578;
      128286:data<=-16'd9503;
      128287:data<=-16'd8922;
      128288:data<=-16'd9935;
      128289:data<=-16'd10252;
      128290:data<=-16'd8778;
      128291:data<=-16'd8951;
      128292:data<=-16'd9401;
      128293:data<=-16'd8208;
      128294:data<=-16'd8319;
      128295:data<=-16'd6904;
      128296:data<=-16'd4845;
      128297:data<=-16'd6986;
      128298:data<=-16'd2667;
      128299:data<=16'd9412;
      128300:data<=16'd12501;
      128301:data<=16'd9477;
      128302:data<=16'd10514;
      128303:data<=16'd10477;
      128304:data<=16'd8731;
      128305:data<=16'd8561;
      128306:data<=16'd8090;
      128307:data<=16'd7630;
      128308:data<=16'd7780;
      128309:data<=16'd8129;
      128310:data<=16'd8440;
      128311:data<=16'd8031;
      128312:data<=16'd8041;
      128313:data<=16'd8000;
      128314:data<=16'd6901;
      128315:data<=16'd6619;
      128316:data<=16'd6733;
      128317:data<=16'd6231;
      128318:data<=16'd6114;
      128319:data<=16'd6023;
      128320:data<=16'd5679;
      128321:data<=16'd4846;
      128322:data<=16'd3641;
      128323:data<=16'd3486;
      128324:data<=16'd3633;
      128325:data<=16'd3741;
      128326:data<=16'd4179;
      128327:data<=16'd3421;
      128328:data<=16'd4244;
      128329:data<=16'd8602;
      128330:data<=16'd11154;
      128331:data<=16'd10851;
      128332:data<=16'd10269;
      128333:data<=16'd9288;
      128334:data<=16'd9768;
      128335:data<=16'd8492;
      128336:data<=16'd85;
      128337:data<=-16'd7585;
      128338:data<=-16'd8237;
      128339:data<=-16'd7776;
      128340:data<=-16'd7785;
      128341:data<=-16'd6909;
      128342:data<=-16'd7136;
      128343:data<=-16'd7215;
      128344:data<=-16'd6554;
      128345:data<=-16'd6405;
      128346:data<=-16'd5833;
      128347:data<=-16'd5653;
      128348:data<=-16'd5832;
      128349:data<=-16'd4978;
      128350:data<=-16'd4939;
      128351:data<=-16'd5090;
      128352:data<=-16'd3721;
      128353:data<=-16'd3171;
      128354:data<=-16'd3491;
      128355:data<=-16'd3178;
      128356:data<=-16'd2708;
      128357:data<=-16'd1976;
      128358:data<=-16'd1591;
      128359:data<=-16'd1621;
      128360:data<=-16'd1237;
      128361:data<=-16'd1168;
      128362:data<=-16'd998;
      128363:data<=-16'd743;
      128364:data<=-16'd977;
      128365:data<=-16'd258;
      128366:data<=16'd182;
      128367:data<=-16'd261;
      128368:data<=16'd144;
      128369:data<=-16'd32;
      128370:data<=16'd886;
      128371:data<=16'd3206;
      128372:data<=16'd2372;
      128373:data<=16'd4267;
      128374:data<=16'd11520;
      128375:data<=16'd13236;
      128376:data<=16'd10989;
      128377:data<=16'd11832;
      128378:data<=16'd11544;
      128379:data<=16'd10352;
      128380:data<=16'd10696;
      128381:data<=16'd10229;
      128382:data<=16'd10013;
      128383:data<=16'd10249;
      128384:data<=16'd9958;
      128385:data<=16'd10002;
      128386:data<=16'd9464;
      128387:data<=16'd9682;
      128388:data<=16'd11300;
      128389:data<=16'd11163;
      128390:data<=16'd10205;
      128391:data<=16'd9962;
      128392:data<=16'd9556;
      128393:data<=16'd9524;
      128394:data<=16'd9235;
      128395:data<=16'd8664;
      128396:data<=16'd8461;
      128397:data<=16'd7483;
      128398:data<=16'd7148;
      128399:data<=16'd7796;
      128400:data<=16'd7197;
      128401:data<=16'd6660;
      128402:data<=16'd6599;
      128403:data<=16'd6161;
      128404:data<=16'd7034;
      128405:data<=16'd8472;
      128406:data<=16'd8831;
      128407:data<=16'd8217;
      128408:data<=16'd7221;
      128409:data<=16'd7877;
      128410:data<=16'd6387;
      128411:data<=-16'd2121;
      128412:data<=-16'd9051;
      128413:data<=-16'd8645;
      128414:data<=-16'd8085;
      128415:data<=-16'd8367;
      128416:data<=-16'd7533;
      128417:data<=-16'd7507;
      128418:data<=-16'd4696;
      128419:data<=-16'd183;
      128420:data<=16'd35;
      128421:data<=-16'd2;
      128422:data<=16'd1818;
      128423:data<=16'd1971;
      128424:data<=16'd2208;
      128425:data<=16'd2309;
      128426:data<=16'd1372;
      128427:data<=16'd1961;
      128428:data<=16'd2646;
      128429:data<=16'd2522;
      128430:data<=16'd2417;
      128431:data<=16'd1723;
      128432:data<=16'd2079;
      128433:data<=16'd2746;
      128434:data<=16'd2287;
      128435:data<=16'd2420;
      128436:data<=16'd2232;
      128437:data<=16'd2419;
      128438:data<=16'd4105;
      128439:data<=16'd4505;
      128440:data<=16'd4300;
      128441:data<=16'd4053;
      128442:data<=16'd3407;
      128443:data<=16'd3751;
      128444:data<=16'd3058;
      128445:data<=16'd3215;
      128446:data<=16'd4473;
      128447:data<=16'd2262;
      128448:data<=16'd6056;
      128449:data<=16'd17374;
      128450:data<=16'd19607;
      128451:data<=16'd16452;
      128452:data<=16'd17590;
      128453:data<=16'd16483;
      128454:data<=16'd15033;
      128455:data<=16'd16920;
      128456:data<=16'd16903;
      128457:data<=16'd16145;
      128458:data<=16'd16160;
      128459:data<=16'd14728;
      128460:data<=16'd13794;
      128461:data<=16'd13940;
      128462:data<=16'd11788;
      128463:data<=16'd7080;
      128464:data<=16'd4378;
      128465:data<=16'd4857;
      128466:data<=16'd4678;
      128467:data<=16'd3783;
      128468:data<=16'd3501;
      128469:data<=16'd2751;
      128470:data<=16'd2532;
      128471:data<=16'd3427;
      128472:data<=16'd4090;
      128473:data<=16'd4055;
      128474:data<=16'd3510;
      128475:data<=16'd3271;
      128476:data<=16'd3362;
      128477:data<=16'd3254;
      128478:data<=16'd3107;
      128479:data<=16'd2682;
      128480:data<=16'd2440;
      128481:data<=16'd2446;
      128482:data<=16'd1689;
      128483:data<=16'd1111;
      128484:data<=16'd1971;
      128485:data<=16'd1262;
      128486:data<=-16'd5524;
      128487:data<=-16'd12942;
      128488:data<=-16'd12205;
      128489:data<=-16'd9310;
      128490:data<=-16'd9914;
      128491:data<=-16'd9256;
      128492:data<=-16'd9101;
      128493:data<=-16'd10320;
      128494:data<=-16'd9318;
      128495:data<=-16'd8912;
      128496:data<=-16'd8848;
      128497:data<=-16'd8235;
      128498:data<=-16'd9059;
      128499:data<=-16'd8446;
      128500:data<=-16'd7824;
      128501:data<=-16'd8552;
      128502:data<=-16'd7562;
      128503:data<=-16'd7445;
      128504:data<=-16'd6910;
      128505:data<=-16'd4837;
      128506:data<=-16'd5462;
      128507:data<=-16'd3955;
      128508:data<=16'd252;
      128509:data<=16'd878;
      128510:data<=16'd497;
      128511:data<=16'd2;
      128512:data<=-16'd889;
      128513:data<=-16'd335;
      128514:data<=-16'd361;
      128515:data<=16'd167;
      128516:data<=16'd256;
      128517:data<=-16'd1404;
      128518:data<=-16'd779;
      128519:data<=-16'd1045;
      128520:data<=-16'd1839;
      128521:data<=16'd155;
      128522:data<=-16'd467;
      128523:data<=16'd3231;
      128524:data<=16'd14443;
      128525:data<=16'd17329;
      128526:data<=16'd14087;
      128527:data<=16'd14736;
      128528:data<=16'd14202;
      128529:data<=16'd12560;
      128530:data<=16'd12090;
      128531:data<=16'd11083;
      128532:data<=16'd11292;
      128533:data<=16'd11688;
      128534:data<=16'd10924;
      128535:data<=16'd10126;
      128536:data<=16'd9069;
      128537:data<=16'd8822;
      128538:data<=16'd9567;
      128539:data<=16'd10025;
      128540:data<=16'd9611;
      128541:data<=16'd8181;
      128542:data<=16'd7598;
      128543:data<=16'd7744;
      128544:data<=16'd6833;
      128545:data<=16'd5940;
      128546:data<=16'd5591;
      128547:data<=16'd5542;
      128548:data<=16'd5388;
      128549:data<=16'd4554;
      128550:data<=16'd4313;
      128551:data<=16'd3516;
      128552:data<=16'd717;
      128553:data<=-16'd1190;
      128554:data<=-16'd1104;
      128555:data<=-16'd293;
      128556:data<=16'd637;
      128557:data<=16'd373;
      128558:data<=-16'd896;
      128559:data<=-16'd951;
      128560:data<=-16'd1671;
      128561:data<=-16'd8305;
      128562:data<=-16'd16337;
      128563:data<=-16'd16800;
      128564:data<=-16'd14747;
      128565:data<=-16'd15555;
      128566:data<=-16'd14888;
      128567:data<=-16'd13958;
      128568:data<=-16'd14173;
      128569:data<=-16'd13646;
      128570:data<=-16'd13998;
      128571:data<=-16'd13221;
      128572:data<=-16'd11204;
      128573:data<=-16'd10978;
      128574:data<=-16'd10006;
      128575:data<=-16'd9479;
      128576:data<=-16'd10539;
      128577:data<=-16'd9646;
      128578:data<=-16'd9075;
      128579:data<=-16'd9276;
      128580:data<=-16'd8457;
      128581:data<=-16'd8863;
      128582:data<=-16'd8883;
      128583:data<=-16'd8150;
      128584:data<=-16'd8210;
      128585:data<=-16'd7233;
      128586:data<=-16'd6896;
      128587:data<=-16'd7233;
      128588:data<=-16'd6141;
      128589:data<=-16'd5303;
      128590:data<=-16'd4269;
      128591:data<=-16'd4032;
      128592:data<=-16'd5021;
      128593:data<=-16'd4252;
      128594:data<=-16'd4817;
      128595:data<=-16'd5541;
      128596:data<=-16'd2749;
      128597:data<=-16'd1400;
      128598:data<=16'd3042;
      128599:data<=16'd13556;
      128600:data<=16'd17042;
      128601:data<=16'd14363;
      128602:data<=16'd14612;
      128603:data<=16'd13903;
      128604:data<=16'd12669;
      128605:data<=16'd13850;
      128606:data<=16'd13850;
      128607:data<=16'd13209;
      128608:data<=16'd12901;
      128609:data<=16'd11893;
      128610:data<=16'd11803;
      128611:data<=16'd11499;
      128612:data<=16'd9787;
      128613:data<=16'd9194;
      128614:data<=16'd9726;
      128615:data<=16'd9445;
      128616:data<=16'd8442;
      128617:data<=16'd8050;
      128618:data<=16'd8161;
      128619:data<=16'd6962;
      128620:data<=16'd5607;
      128621:data<=16'd5729;
      128622:data<=16'd5210;
      128623:data<=16'd4537;
      128624:data<=16'd4934;
      128625:data<=16'd4188;
      128626:data<=16'd3618;
      128627:data<=16'd4356;
      128628:data<=16'd3852;
      128629:data<=16'd3054;
      128630:data<=16'd2661;
      128631:data<=16'd2099;
      128632:data<=16'd2305;
      128633:data<=16'd1694;
      128634:data<=16'd1474;
      128635:data<=16'd1334;
      128636:data<=-16'd5589;
      128637:data<=-16'd14075;
      128638:data<=-16'd15185;
      128639:data<=-16'd14838;
      128640:data<=-16'd16269;
      128641:data<=-16'd17373;
      128642:data<=-16'd19237;
      128643:data<=-16'd19133;
      128644:data<=-16'd17482;
      128645:data<=-16'd17490;
      128646:data<=-16'd16883;
      128647:data<=-16'd16177;
      128648:data<=-16'd16020;
      128649:data<=-16'd14872;
      128650:data<=-16'd14872;
      128651:data<=-16'd15051;
      128652:data<=-16'd13990;
      128653:data<=-16'd13582;
      128654:data<=-16'd12881;
      128655:data<=-16'd12918;
      128656:data<=-16'd14418;
      128657:data<=-16'd14157;
      128658:data<=-16'd13368;
      128659:data<=-16'd13261;
      128660:data<=-16'd12505;
      128661:data<=-16'd12452;
      128662:data<=-16'd12468;
      128663:data<=-16'd11637;
      128664:data<=-16'd11004;
      128665:data<=-16'd10355;
      128666:data<=-16'd10363;
      128667:data<=-16'd10076;
      128668:data<=-16'd9045;
      128669:data<=-16'd9638;
      128670:data<=-16'd9047;
      128671:data<=-16'd8064;
      128672:data<=-16'd10845;
      128673:data<=-16'd7721;
      128674:data<=16'd3430;
      128675:data<=16'd7259;
      128676:data<=16'd4792;
      128677:data<=16'd5794;
      128678:data<=16'd5927;
      128679:data<=16'd4643;
      128680:data<=16'd5288;
      128681:data<=16'd4798;
      128682:data<=16'd4684;
      128683:data<=16'd5466;
      128684:data<=16'd4123;
      128685:data<=16'd4915;
      128686:data<=16'd8176;
      128687:data<=16'd8525;
      128688:data<=16'd7218;
      128689:data<=16'd5923;
      128690:data<=16'd4908;
      128691:data<=16'd5333;
      128692:data<=16'd5253;
      128693:data<=16'd4619;
      128694:data<=16'd4431;
      128695:data<=16'd3943;
      128696:data<=16'd4338;
      128697:data<=16'd4215;
      128698:data<=16'd2729;
      128699:data<=16'd2699;
      128700:data<=16'd2839;
      128701:data<=16'd2587;
      128702:data<=16'd2968;
      128703:data<=16'd2634;
      128704:data<=16'd2917;
      128705:data<=16'd2291;
      128706:data<=-16'd176;
      128707:data<=-16'd88;
      128708:data<=-16'd274;
      128709:data<=-16'd887;
      128710:data<=16'd523;
      128711:data<=-16'd5576;
      128712:data<=-16'd15194;
      128713:data<=-16'd15154;
      128714:data<=-16'd13285;
      128715:data<=-16'd14316;
      128716:data<=-16'd13239;
      128717:data<=-16'd13341;
      128718:data<=-16'd13380;
      128719:data<=-16'd11723;
      128720:data<=-16'd12020;
      128721:data<=-16'd12051;
      128722:data<=-16'd12140;
      128723:data<=-16'd13080;
      128724:data<=-16'd11900;
      128725:data<=-16'd11432;
      128726:data<=-16'd11549;
      128727:data<=-16'd10100;
      128728:data<=-16'd9809;
      128729:data<=-16'd9409;
      128730:data<=-16'd10160;
      128731:data<=-16'd13841;
      128732:data<=-16'd14093;
      128733:data<=-16'd11768;
      128734:data<=-16'd11555;
      128735:data<=-16'd11210;
      128736:data<=-16'd10681;
      128737:data<=-16'd10037;
      128738:data<=-16'd9204;
      128739:data<=-16'd10140;
      128740:data<=-16'd10592;
      128741:data<=-16'd10138;
      128742:data<=-16'd9573;
      128743:data<=-16'd7882;
      128744:data<=-16'd7956;
      128745:data<=-16'd7987;
      128746:data<=-16'd6764;
      128747:data<=-16'd8519;
      128748:data<=-16'd4655;
      128749:data<=16'd6933;
      128750:data<=16'd10290;
      128751:data<=16'd7392;
      128752:data<=16'd8561;
      128753:data<=16'd9194;
      128754:data<=16'd8813;
      128755:data<=16'd8809;
      128756:data<=16'd6281;
      128757:data<=16'd5313;
      128758:data<=16'd6522;
      128759:data<=16'd5915;
      128760:data<=16'd5288;
      128761:data<=16'd4921;
      128762:data<=16'd4432;
      128763:data<=16'd5106;
      128764:data<=16'd5100;
      128765:data<=16'd4764;
      128766:data<=16'd5125;
      128767:data<=16'd5069;
      128768:data<=16'd5554;
      128769:data<=16'd5028;
      128770:data<=16'd3383;
      128771:data<=16'd4517;
      128772:data<=16'd4511;
      128773:data<=16'd1535;
      128774:data<=16'd2403;
      128775:data<=16'd5336;
      128776:data<=16'd5977;
      128777:data<=16'd6331;
      128778:data<=16'd5887;
      128779:data<=16'd5234;
      128780:data<=16'd5426;
      128781:data<=16'd4980;
      128782:data<=16'd5395;
      128783:data<=16'd5228;
      128784:data<=16'd4384;
      128785:data<=16'd5288;
      128786:data<=16'd18;
      128787:data<=-16'd9837;
      128788:data<=-16'd11596;
      128789:data<=-16'd10951;
      128790:data<=-16'd12907;
      128791:data<=-16'd11345;
      128792:data<=-16'd10290;
      128793:data<=-16'd10781;
      128794:data<=-16'd9459;
      128795:data<=-16'd9679;
      128796:data<=-16'd9527;
      128797:data<=-16'd8308;
      128798:data<=-16'd8658;
      128799:data<=-16'd7770;
      128800:data<=-16'd7266;
      128801:data<=-16'd7973;
      128802:data<=-16'd7207;
      128803:data<=-16'd7107;
      128804:data<=-16'd6346;
      128805:data<=-16'd5536;
      128806:data<=-16'd7617;
      128807:data<=-16'd7521;
      128808:data<=-16'd6085;
      128809:data<=-16'd6399;
      128810:data<=-16'd5369;
      128811:data<=-16'd5322;
      128812:data<=-16'd5532;
      128813:data<=-16'd3795;
      128814:data<=-16'd3946;
      128815:data<=-16'd3651;
      128816:data<=-16'd2919;
      128817:data<=-16'd3500;
      128818:data<=-16'd1683;
      128819:data<=-16'd2884;
      128820:data<=-16'd6661;
      128821:data<=-16'd5847;
      128822:data<=-16'd6796;
      128823:data<=-16'd4886;
      128824:data<=16'd5909;
      128825:data<=16'd9800;
      128826:data<=16'd7298;
      128827:data<=16'd9333;
      128828:data<=16'd9206;
      128829:data<=16'd7632;
      128830:data<=16'd9135;
      128831:data<=16'd8655;
      128832:data<=16'd7837;
      128833:data<=16'd8420;
      128834:data<=16'd8011;
      128835:data<=16'd8087;
      128836:data<=16'd7771;
      128837:data<=16'd6863;
      128838:data<=16'd7128;
      128839:data<=16'd6446;
      128840:data<=16'd5112;
      128841:data<=16'd4817;
      128842:data<=16'd4589;
      128843:data<=16'd4807;
      128844:data<=16'd5062;
      128845:data<=16'd4713;
      128846:data<=16'd4711;
      128847:data<=16'd4294;
      128848:data<=16'd4014;
      128849:data<=16'd4584;
      128850:data<=16'd4062;
      128851:data<=16'd3506;
      128852:data<=16'd3535;
      128853:data<=16'd2783;
      128854:data<=16'd3245;
      128855:data<=16'd3359;
      128856:data<=16'd1438;
      128857:data<=16'd1598;
      128858:data<=16'd1726;
      128859:data<=16'd1007;
      128860:data<=16'd2742;
      128861:data<=-16'd2011;
      128862:data<=-16'd12801;
      128863:data<=-16'd14237;
      128864:data<=-16'd9966;
      128865:data<=-16'd8907;
      128866:data<=-16'd7512;
      128867:data<=-16'd7063;
      128868:data<=-16'd7783;
      128869:data<=-16'd6815;
      128870:data<=-16'd6598;
      128871:data<=-16'd6328;
      128872:data<=-16'd6184;
      128873:data<=-16'd7608;
      128874:data<=-16'd7203;
      128875:data<=-16'd6455;
      128876:data<=-16'd6772;
      128877:data<=-16'd6049;
      128878:data<=-16'd6153;
      128879:data<=-16'd6029;
      128880:data<=-16'd5077;
      128881:data<=-16'd5357;
      128882:data<=-16'd4112;
      128883:data<=-16'd2719;
      128884:data<=-16'd3442;
      128885:data<=-16'd3039;
      128886:data<=-16'd2617;
      128887:data<=-16'd2632;
      128888:data<=-16'd1771;
      128889:data<=-16'd1706;
      128890:data<=-16'd1134;
      128891:data<=-16'd925;
      128892:data<=-16'd1827;
      128893:data<=-16'd817;
      128894:data<=-16'd646;
      128895:data<=-16'd792;
      128896:data<=16'd429;
      128897:data<=-16'd1357;
      128898:data<=16'd1832;
      128899:data<=16'd13071;
      128900:data<=16'd16756;
      128901:data<=16'd14254;
      128902:data<=16'd15446;
      128903:data<=16'd15173;
      128904:data<=16'd13638;
      128905:data<=16'd14217;
      128906:data<=16'd14489;
      128907:data<=16'd15807;
      128908:data<=16'd15393;
      128909:data<=16'd10921;
      128910:data<=16'd9266;
      128911:data<=16'd10194;
      128912:data<=16'd9429;
      128913:data<=16'd9172;
      128914:data<=16'd8987;
      128915:data<=16'd8116;
      128916:data<=16'd8308;
      128917:data<=16'd8341;
      128918:data<=16'd8217;
      128919:data<=16'd8090;
      128920:data<=16'd6877;
      128921:data<=16'd6693;
      128922:data<=16'd7632;
      128923:data<=16'd8207;
      128924:data<=16'd8805;
      128925:data<=16'd8026;
      128926:data<=16'd7156;
      128927:data<=16'd7680;
      128928:data<=16'd6927;
      128929:data<=16'd6508;
      128930:data<=16'd6949;
      128931:data<=16'd6147;
      128932:data<=16'd6724;
      128933:data<=16'd6616;
      128934:data<=16'd5603;
      128935:data<=16'd7507;
      128936:data<=16'd2860;
      128937:data<=-16'd8539;
      128938:data<=-16'd11168;
      128939:data<=-16'd8278;
      128940:data<=-16'd8046;
      128941:data<=-16'd6896;
      128942:data<=-16'd6449;
      128943:data<=-16'd6895;
      128944:data<=-16'd5896;
      128945:data<=-16'd6088;
      128946:data<=-16'd6070;
      128947:data<=-16'd5498;
      128948:data<=-16'd6122;
      128949:data<=-16'd5385;
      128950:data<=-16'd4479;
      128951:data<=-16'd4933;
      128952:data<=-16'd4358;
      128953:data<=-16'd2343;
      128954:data<=16'd237;
      128955:data<=16'd873;
      128956:data<=16'd438;
      128957:data<=16'd2405;
      128958:data<=16'd3133;
      128959:data<=16'd2196;
      128960:data<=16'd3175;
      128961:data<=16'd3028;
      128962:data<=16'd2129;
      128963:data<=16'd2581;
      128964:data<=16'd2375;
      128965:data<=16'd2813;
      128966:data<=16'd2931;
      128967:data<=16'd1817;
      128968:data<=16'd2488;
      128969:data<=16'd2507;
      128970:data<=16'd1988;
      128971:data<=16'd2593;
      128972:data<=16'd1313;
      128973:data<=16'd5432;
      128974:data<=16'd16909;
      128975:data<=16'd20862;
      128976:data<=16'd17935;
      128977:data<=16'd18258;
      128978:data<=16'd18274;
      128979:data<=16'd16950;
      128980:data<=16'd16850;
      128981:data<=16'd15805;
      128982:data<=16'd15329;
      128983:data<=16'd15673;
      128984:data<=16'd14616;
      128985:data<=16'd14143;
      128986:data<=16'd13843;
      128987:data<=16'd12433;
      128988:data<=16'd11929;
      128989:data<=16'd12138;
      128990:data<=16'd12578;
      128991:data<=16'd12983;
      128992:data<=16'd12283;
      128993:data<=16'd11937;
      128994:data<=16'd11447;
      128995:data<=16'd10246;
      128996:data<=16'd10630;
      128997:data<=16'd9529;
      128998:data<=16'd5883;
      128999:data<=16'd4672;
      129000:data<=16'd4343;
      129001:data<=16'd3112;
      129002:data<=16'd3057;
      129003:data<=16'd2796;
      129004:data<=16'd2649;
      129005:data<=16'd2393;
      129006:data<=16'd1604;
      129007:data<=16'd3626;
      129008:data<=16'd4390;
      129009:data<=16'd2898;
      129010:data<=16'd4608;
      129011:data<=16'd370;
      129012:data<=-16'd10675;
      129013:data<=-16'd12860;
      129014:data<=-16'd10463;
      129015:data<=-16'd12105;
      129016:data<=-16'd11785;
      129017:data<=-16'd10874;
      129018:data<=-16'd11577;
      129019:data<=-16'd10733;
      129020:data<=-16'd10561;
      129021:data<=-16'd10913;
      129022:data<=-16'd10009;
      129023:data<=-16'd8893;
      129024:data<=-16'd7291;
      129025:data<=-16'd6684;
      129026:data<=-16'd7034;
      129027:data<=-16'd6322;
      129028:data<=-16'd5955;
      129029:data<=-16'd5973;
      129030:data<=-16'd5814;
      129031:data<=-16'd5921;
      129032:data<=-16'd5312;
      129033:data<=-16'd4946;
      129034:data<=-16'd4986;
      129035:data<=-16'd4472;
      129036:data<=-16'd4388;
      129037:data<=-16'd4184;
      129038:data<=-16'd4109;
      129039:data<=-16'd3667;
      129040:data<=-16'd1619;
      129041:data<=-16'd1659;
      129042:data<=-16'd1348;
      129043:data<=16'd2746;
      129044:data<=16'd3419;
      129045:data<=16'd2290;
      129046:data<=16'd3503;
      129047:data<=16'd1541;
      129048:data<=16'd3647;
      129049:data<=16'd14249;
      129050:data<=16'd18776;
      129051:data<=16'd16419;
      129052:data<=16'd16271;
      129053:data<=16'd15858;
      129054:data<=16'd14751;
      129055:data<=16'd14941;
      129056:data<=16'd14851;
      129057:data<=16'd15276;
      129058:data<=16'd15467;
      129059:data<=16'd14195;
      129060:data<=16'd13306;
      129061:data<=16'd12772;
      129062:data<=16'd12157;
      129063:data<=16'd11585;
      129064:data<=16'd10543;
      129065:data<=16'd10053;
      129066:data<=16'd9899;
      129067:data<=16'd9283;
      129068:data<=16'd9321;
      129069:data<=16'd9051;
      129070:data<=16'd8035;
      129071:data<=16'd7811;
      129072:data<=16'd7435;
      129073:data<=16'd7638;
      129074:data<=16'd9309;
      129075:data<=16'd9156;
      129076:data<=16'd7774;
      129077:data<=16'd7151;
      129078:data<=16'd5924;
      129079:data<=16'd5841;
      129080:data<=16'd6132;
      129081:data<=16'd4673;
      129082:data<=16'd4775;
      129083:data<=16'd4323;
      129084:data<=16'd3180;
      129085:data<=16'd5579;
      129086:data<=16'd693;
      129087:data<=-16'd13042;
      129088:data<=-16'd17517;
      129089:data<=-16'd14681;
      129090:data<=-16'd14944;
      129091:data<=-16'd13929;
      129092:data<=-16'd12625;
      129093:data<=-16'd13065;
      129094:data<=-16'd12273;
      129095:data<=-16'd12777;
      129096:data<=-16'd13361;
      129097:data<=-16'd11844;
      129098:data<=-16'd11444;
      129099:data<=-16'd11298;
      129100:data<=-16'd10689;
      129101:data<=-16'd10719;
      129102:data<=-16'd10158;
      129103:data<=-16'd9555;
      129104:data<=-16'd9304;
      129105:data<=-16'd9304;
      129106:data<=-16'd9218;
      129107:data<=-16'd7579;
      129108:data<=-16'd6398;
      129109:data<=-16'd6385;
      129110:data<=-16'd6076;
      129111:data<=-16'd6473;
      129112:data<=-16'd6088;
      129113:data<=-16'd5186;
      129114:data<=-16'd5506;
      129115:data<=-16'd4899;
      129116:data<=-16'd5332;
      129117:data<=-16'd6229;
      129118:data<=-16'd4316;
      129119:data<=-16'd4595;
      129120:data<=-16'd5377;
      129121:data<=-16'd3741;
      129122:data<=-16'd5436;
      129123:data<=-16'd2528;
      129124:data<=16'd9175;
      129125:data<=16'd14076;
      129126:data<=16'd11599;
      129127:data<=16'd11729;
      129128:data<=16'd12260;
      129129:data<=16'd11726;
      129130:data<=16'd11307;
      129131:data<=16'd11409;
      129132:data<=16'd13805;
      129133:data<=16'd15086;
      129134:data<=16'd13276;
      129135:data<=16'd12460;
      129136:data<=16'd12549;
      129137:data<=16'd11670;
      129138:data<=16'd10985;
      129139:data<=16'd10505;
      129140:data<=16'd10185;
      129141:data<=16'd10739;
      129142:data<=16'd11136;
      129143:data<=16'd10818;
      129144:data<=16'd10325;
      129145:data<=16'd9451;
      129146:data<=16'd8772;
      129147:data<=16'd8695;
      129148:data<=16'd8402;
      129149:data<=16'd7849;
      129150:data<=16'd6717;
      129151:data<=16'd5536;
      129152:data<=16'd5410;
      129153:data<=16'd4899;
      129154:data<=16'd4493;
      129155:data<=16'd4733;
      129156:data<=16'd3761;
      129157:data<=16'd3463;
      129158:data<=16'd3189;
      129159:data<=16'd2337;
      129160:data<=16'd4444;
      129161:data<=16'd752;
      129162:data<=-16'd11106;
      129163:data<=-16'd14316;
      129164:data<=-16'd11141;
      129165:data<=-16'd12874;
      129166:data<=-16'd13086;
      129167:data<=-16'd11664;
      129168:data<=-16'd12363;
      129169:data<=-16'd11773;
      129170:data<=-16'd11969;
      129171:data<=-16'd12181;
      129172:data<=-16'd10473;
      129173:data<=-16'd11094;
      129174:data<=-16'd12270;
      129175:data<=-16'd12269;
      129176:data<=-16'd13803;
      129177:data<=-16'd15279;
      129178:data<=-16'd15383;
      129179:data<=-16'd14804;
      129180:data<=-16'd14345;
      129181:data<=-16'd14407;
      129182:data<=-16'd13872;
      129183:data<=-16'd13766;
      129184:data<=-16'd13662;
      129185:data<=-16'd12248;
      129186:data<=-16'd12002;
      129187:data<=-16'd12026;
      129188:data<=-16'd10988;
      129189:data<=-16'd10463;
      129190:data<=-16'd9926;
      129191:data<=-16'd10731;
      129192:data<=-16'd11673;
      129193:data<=-16'd10214;
      129194:data<=-16'd10404;
      129195:data<=-16'd10575;
      129196:data<=-16'd8981;
      129197:data<=-16'd10698;
      129198:data<=-16'd8396;
      129199:data<=16'd2223;
      129200:data<=16'd7796;
      129201:data<=16'd6343;
      129202:data<=16'd6288;
      129203:data<=16'd6630;
      129204:data<=16'd6199;
      129205:data<=16'd6255;
      129206:data<=16'd5040;
      129207:data<=16'd3466;
      129208:data<=16'd3483;
      129209:data<=16'd3404;
      129210:data<=16'd2723;
      129211:data<=16'd2711;
      129212:data<=16'd2576;
      129213:data<=16'd2173;
      129214:data<=16'd2276;
      129215:data<=16'd1967;
      129216:data<=16'd1527;
      129217:data<=16'd1815;
      129218:data<=16'd1871;
      129219:data<=16'd1697;
      129220:data<=16'd2641;
      129221:data<=16'd4693;
      129222:data<=16'd5482;
      129223:data<=16'd4317;
      129224:data<=16'd3501;
      129225:data<=16'd2698;
      129226:data<=16'd1580;
      129227:data<=16'd1407;
      129228:data<=16'd992;
      129229:data<=16'd1019;
      129230:data<=16'd1216;
      129231:data<=16'd217;
      129232:data<=16'd1293;
      129233:data<=16'd1606;
      129234:data<=-16'd446;
      129235:data<=16'd970;
      129236:data<=-16'd2428;
      129237:data<=-16'd13565;
      129238:data<=-16'd16530;
      129239:data<=-16'd13744;
      129240:data<=-16'd15573;
      129241:data<=-16'd16443;
      129242:data<=-16'd15346;
      129243:data<=-16'd15076;
      129244:data<=-16'd14427;
      129245:data<=-16'd14731;
      129246:data<=-16'd14892;
      129247:data<=-16'd13881;
      129248:data<=-16'd13164;
      129249:data<=-16'd12393;
      129250:data<=-16'd12084;
      129251:data<=-16'd11614;
      129252:data<=-16'd10502;
      129253:data<=-16'd10270;
      129254:data<=-16'd9862;
      129255:data<=-16'd9285;
      129256:data<=-16'd9433;
      129257:data<=-16'd9949;
      129258:data<=-16'd11326;
      129259:data<=-16'd11402;
      129260:data<=-16'd10016;
      129261:data<=-16'd10009;
      129262:data<=-16'd9744;
      129263:data<=-16'd8860;
      129264:data<=-16'd8467;
      129265:data<=-16'd8455;
      129266:data<=-16'd10564;
      129267:data<=-16'd11568;
      129268:data<=-16'd9676;
      129269:data<=-16'd9959;
      129270:data<=-16'd10103;
      129271:data<=-16'd8288;
      129272:data<=-16'd9132;
      129273:data<=-16'd7586;
      129274:data<=16'd534;
      129275:data<=16'd6387;
      129276:data<=16'd6187;
      129277:data<=16'd5620;
      129278:data<=16'd6031;
      129279:data<=16'd5683;
      129280:data<=16'd5827;
      129281:data<=16'd6041;
      129282:data<=16'd5463;
      129283:data<=16'd5987;
      129284:data<=16'd6234;
      129285:data<=16'd5221;
      129286:data<=16'd5560;
      129287:data<=16'd5676;
      129288:data<=16'd4711;
      129289:data<=16'd4996;
      129290:data<=16'd4446;
      129291:data<=16'd2406;
      129292:data<=16'd1894;
      129293:data<=16'd2378;
      129294:data<=16'd2217;
      129295:data<=16'd2112;
      129296:data<=16'd2315;
      129297:data<=16'd1670;
      129298:data<=16'd1199;
      129299:data<=16'd2112;
      129300:data<=16'd2121;
      129301:data<=16'd1742;
      129302:data<=16'd2006;
      129303:data<=16'd967;
      129304:data<=16'd966;
      129305:data<=16'd1823;
      129306:data<=16'd1025;
      129307:data<=16'd1011;
      129308:data<=-16'd688;
      129309:data<=-16'd1454;
      129310:data<=16'd4212;
      129311:data<=16'd1970;
      129312:data<=-16'd10393;
      129313:data<=-16'd13693;
      129314:data<=-16'd10906;
      129315:data<=-16'd11527;
      129316:data<=-16'd10657;
      129317:data<=-16'd9762;
      129318:data<=-16'd10035;
      129319:data<=-16'd8777;
      129320:data<=-16'd8831;
      129321:data<=-16'd9259;
      129322:data<=-16'd8167;
      129323:data<=-16'd7988;
      129324:data<=-16'd8871;
      129325:data<=-16'd9577;
      129326:data<=-16'd9027;
      129327:data<=-16'd7931;
      129328:data<=-16'd7780;
      129329:data<=-16'd7256;
      129330:data<=-16'd6831;
      129331:data<=-16'd7244;
      129332:data<=-16'd6769;
      129333:data<=-16'd6219;
      129334:data<=-16'd6102;
      129335:data<=-16'd5503;
      129336:data<=-16'd5077;
      129337:data<=-16'd4607;
      129338:data<=-16'd3853;
      129339:data<=-16'd3068;
      129340:data<=-16'd2602;
      129341:data<=-16'd3489;
      129342:data<=-16'd4099;
      129343:data<=-16'd3442;
      129344:data<=-16'd3673;
      129345:data<=-16'd3732;
      129346:data<=-16'd3054;
      129347:data<=-16'd3952;
      129348:data<=-16'd2044;
      129349:data<=16'd6936;
      129350:data<=16'd14126;
      129351:data<=16'd13127;
      129352:data<=16'd12217;
      129353:data<=16'd14029;
      129354:data<=16'd11782;
      129355:data<=16'd8144;
      129356:data<=16'd7636;
      129357:data<=16'd6887;
      129358:data<=16'd5612;
      129359:data<=16'd5362;
      129360:data<=16'd5069;
      129361:data<=16'd5269;
      129362:data<=16'd5571;
      129363:data<=16'd5062;
      129364:data<=16'd4895;
      129365:data<=16'd4872;
      129366:data<=16'd4510;
      129367:data<=16'd4660;
      129368:data<=16'd5004;
      129369:data<=16'd4937;
      129370:data<=16'd5065;
      129371:data<=16'd5083;
      129372:data<=16'd4455;
      129373:data<=16'd4425;
      129374:data<=16'd3756;
      129375:data<=16'd1409;
      129376:data<=16'd1416;
      129377:data<=16'd2416;
      129378:data<=16'd1045;
      129379:data<=16'd1512;
      129380:data<=16'd2214;
      129381:data<=16'd846;
      129382:data<=16'd2272;
      129383:data<=16'd2221;
      129384:data<=16'd328;
      129385:data<=16'd3243;
      129386:data<=16'd26;
      129387:data<=-16'd11640;
      129388:data<=-16'd14675;
      129389:data<=-16'd11724;
      129390:data<=-16'd12901;
      129391:data<=-16'd13559;
      129392:data<=-16'd12918;
      129393:data<=-16'd13089;
      129394:data<=-16'd12398;
      129395:data<=-16'd11819;
      129396:data<=-16'd11668;
      129397:data<=-16'd11662;
      129398:data<=-16'd11136;
      129399:data<=-16'd8128;
      129400:data<=-16'd5162;
      129401:data<=-16'd4387;
      129402:data<=-16'd3908;
      129403:data<=-16'd3777;
      129404:data<=-16'd3853;
      129405:data<=-16'd3193;
      129406:data<=-16'd2773;
      129407:data<=-16'd3069;
      129408:data<=-16'd4059;
      129409:data<=-16'd4734;
      129410:data<=-16'd4079;
      129411:data<=-16'd3644;
      129412:data<=-16'd3240;
      129413:data<=-16'd2214;
      129414:data<=-16'd2347;
      129415:data<=-16'd2328;
      129416:data<=-16'd1169;
      129417:data<=-16'd843;
      129418:data<=-16'd328;
      129419:data<=16'd59;
      129420:data<=-16'd678;
      129421:data<=-16'd9;
      129422:data<=16'd174;
      129423:data<=16'd917;
      129424:data<=16'd9033;
      129425:data<=16'd17106;
      129426:data<=16'd16302;
      129427:data<=16'd14822;
      129428:data<=16'd15767;
      129429:data<=16'd14684;
      129430:data<=16'd14457;
      129431:data<=16'd15073;
      129432:data<=16'd14057;
      129433:data<=16'd13844;
      129434:data<=16'd14113;
      129435:data<=16'd13741;
      129436:data<=16'd13675;
      129437:data<=16'd13176;
      129438:data<=16'd12612;
      129439:data<=16'd12273;
      129440:data<=16'd11624;
      129441:data<=16'd12214;
      129442:data<=16'd13370;
      129443:data<=16'd12128;
      129444:data<=16'd9037;
      129445:data<=16'd7445;
      129446:data<=16'd7870;
      129447:data<=16'd7595;
      129448:data<=16'd7247;
      129449:data<=16'd7955;
      129450:data<=16'd7098;
      129451:data<=16'd6111;
      129452:data<=16'd6478;
      129453:data<=16'd5615;
      129454:data<=16'd5416;
      129455:data<=16'd5735;
      129456:data<=16'd4679;
      129457:data<=16'd6068;
      129458:data<=16'd7221;
      129459:data<=16'd6363;
      129460:data<=16'd8240;
      129461:data<=16'd4376;
      129462:data<=-16'd7037;
      129463:data<=-16'd10163;
      129464:data<=-16'd7436;
      129465:data<=-16'd8728;
      129466:data<=-16'd8589;
      129467:data<=-16'd7219;
      129468:data<=-16'd8058;
      129469:data<=-16'd7608;
      129470:data<=-16'd6836;
      129471:data<=-16'd6990;
      129472:data<=-16'd6684;
      129473:data<=-16'd6381;
      129474:data<=-16'd5171;
      129475:data<=-16'd3794;
      129476:data<=-16'd3518;
      129477:data<=-16'd2955;
      129478:data<=-16'd2622;
      129479:data<=-16'd2311;
      129480:data<=-16'd1522;
      129481:data<=-16'd1689;
      129482:data<=-16'd1647;
      129483:data<=-16'd1481;
      129484:data<=-16'd2049;
      129485:data<=-16'd1530;
      129486:data<=-16'd1510;
      129487:data<=-16'd1676;
      129488:data<=16'd1280;
      129489:data<=16'd3853;
      129490:data<=16'd4258;
      129491:data<=16'd5527;
      129492:data<=16'd6724;
      129493:data<=16'd7103;
      129494:data<=16'd6708;
      129495:data<=16'd5852;
      129496:data<=16'd6690;
      129497:data<=16'd6378;
      129498:data<=16'd6122;
      129499:data<=16'd13529;
      129500:data<=16'd21528;
      129501:data<=16'd21083;
      129502:data<=16'd19713;
      129503:data<=16'd20212;
      129504:data<=16'd18578;
      129505:data<=16'd17760;
      129506:data<=16'd17788;
      129507:data<=16'd17029;
      129508:data<=16'd17966;
      129509:data<=16'd18727;
      129510:data<=16'd17855;
      129511:data<=16'd17526;
      129512:data<=16'd16727;
      129513:data<=16'd15682;
      129514:data<=16'd15756;
      129515:data<=16'd15288;
      129516:data<=16'd14273;
      129517:data<=16'd13506;
      129518:data<=16'd12765;
      129519:data<=16'd12455;
      129520:data<=16'd12245;
      129521:data<=16'd12066;
      129522:data<=16'd11536;
      129523:data<=16'd10339;
      129524:data<=16'd10399;
      129525:data<=16'd11194;
      129526:data<=16'd11126;
      129527:data<=16'd10850;
      129528:data<=16'd9829;
      129529:data<=16'd9041;
      129530:data<=16'd9185;
      129531:data<=16'd8525;
      129532:data<=16'd7612;
      129533:data<=16'd4854;
      129534:data<=16'd1820;
      129535:data<=16'd3409;
      129536:data<=16'd88;
      129537:data<=-16'd11157;
      129538:data<=-16'd14343;
      129539:data<=-16'd11236;
      129540:data<=-16'd12393;
      129541:data<=-16'd11673;
      129542:data<=-16'd8839;
      129543:data<=-16'd9341;
      129544:data<=-16'd9632;
      129545:data<=-16'd9030;
      129546:data<=-16'd9113;
      129547:data<=-16'd8903;
      129548:data<=-16'd8731;
      129549:data<=-16'd8055;
      129550:data<=-16'd7282;
      129551:data<=-16'd7447;
      129552:data<=-16'd7509;
      129553:data<=-16'd7489;
      129554:data<=-16'd7056;
      129555:data<=-16'd6272;
      129556:data<=-16'd6583;
      129557:data<=-16'd6299;
      129558:data<=-16'd4595;
      129559:data<=-16'd3507;
      129560:data<=-16'd3275;
      129561:data<=-16'd3422;
      129562:data<=-16'd2860;
      129563:data<=-16'd1668;
      129564:data<=-16'd2259;
      129565:data<=-16'd3011;
      129566:data<=-16'd2291;
      129567:data<=-16'd2393;
      129568:data<=-16'd2170;
      129569:data<=-16'd1574;
      129570:data<=-16'd2520;
      129571:data<=-16'd1880;
      129572:data<=-16'd1486;
      129573:data<=-16'd2378;
      129574:data<=16'd5222;
      129575:data<=16'd15901;
      129576:data<=16'd15858;
      129577:data<=16'd14478;
      129578:data<=16'd18160;
      129579:data<=16'd17837;
      129580:data<=16'd16111;
      129581:data<=16'd16449;
      129582:data<=16'd15473;
      129583:data<=16'd15547;
      129584:data<=16'd15524;
      129585:data<=16'd13628;
      129586:data<=16'd13123;
      129587:data<=16'd12709;
      129588:data<=16'd12240;
      129589:data<=16'd12272;
      129590:data<=16'd10696;
      129591:data<=16'd10473;
      129592:data<=16'd11740;
      129593:data<=16'd11383;
      129594:data<=16'd10968;
      129595:data<=16'd10056;
      129596:data<=16'd8983;
      129597:data<=16'd9476;
      129598:data<=16'd9159;
      129599:data<=16'd8202;
      129600:data<=16'd7594;
      129601:data<=16'd6708;
      129602:data<=16'd6266;
      129603:data<=16'd5544;
      129604:data<=16'd5300;
      129605:data<=16'd5139;
      129606:data<=16'd3626;
      129607:data<=16'd4341;
      129608:data<=16'd5219;
      129609:data<=16'd4631;
      129610:data<=16'd6830;
      129611:data<=16'd3089;
      129612:data<=-16'd8420;
      129613:data<=-16'd12014;
      129614:data<=-16'd9561;
      129615:data<=-16'd10295;
      129616:data<=-16'd10273;
      129617:data<=-16'd9606;
      129618:data<=-16'd10151;
      129619:data<=-16'd9896;
      129620:data<=-16'd9973;
      129621:data<=-16'd10727;
      129622:data<=-16'd12328;
      129623:data<=-16'd14389;
      129624:data<=-16'd13853;
      129625:data<=-16'd11814;
      129626:data<=-16'd10733;
      129627:data<=-16'd10246;
      129628:data<=-16'd10349;
      129629:data<=-16'd10146;
      129630:data<=-16'd9288;
      129631:data<=-16'd9147;
      129632:data<=-16'd9256;
      129633:data<=-16'd9094;
      129634:data<=-16'd9294;
      129635:data<=-16'd9326;
      129636:data<=-16'd8987;
      129637:data<=-16'd8652;
      129638:data<=-16'd7730;
      129639:data<=-16'd7075;
      129640:data<=-16'd7467;
      129641:data<=-16'd6805;
      129642:data<=-16'd5233;
      129643:data<=-16'd4608;
      129644:data<=-16'd4560;
      129645:data<=-16'd4749;
      129646:data<=-16'd4081;
      129647:data<=-16'd3961;
      129648:data<=-16'd4922;
      129649:data<=16'd1425;
      129650:data<=16'd11617;
      129651:data<=16'd11888;
      129652:data<=16'd8856;
      129653:data<=16'd9814;
      129654:data<=16'd8611;
      129655:data<=16'd7885;
      129656:data<=16'd8651;
      129657:data<=16'd7679;
      129658:data<=16'd8751;
      129659:data<=16'd9576;
      129660:data<=16'd8337;
      129661:data<=16'd8648;
      129662:data<=16'd8164;
      129663:data<=16'd7418;
      129664:data<=16'd7421;
      129665:data<=16'd6087;
      129666:data<=16'd7090;
      129667:data<=16'd9470;
      129668:data<=16'd9257;
      129669:data<=16'd8675;
      129670:data<=16'd8009;
      129671:data<=16'd7574;
      129672:data<=16'd7780;
      129673:data<=16'd6898;
      129674:data<=16'd6422;
      129675:data<=16'd6120;
      129676:data<=16'd5705;
      129677:data<=16'd6475;
      129678:data<=16'd6140;
      129679:data<=16'd5533;
      129680:data<=16'd5156;
      129681:data<=16'd3694;
      129682:data<=16'd4208;
      129683:data<=16'd3971;
      129684:data<=16'd2488;
      129685:data<=16'd4460;
      129686:data<=16'd602;
      129687:data<=-16'd10678;
      129688:data<=-16'd14357;
      129689:data<=-16'd12031;
      129690:data<=-16'd12422;
      129691:data<=-16'd12681;
      129692:data<=-16'd12154;
      129693:data<=-16'd12255;
      129694:data<=-16'd11952;
      129695:data<=-16'd11822;
      129696:data<=-16'd11812;
      129697:data<=-16'd11311;
      129698:data<=-16'd10651;
      129699:data<=-16'd10378;
      129700:data<=-16'd10627;
      129701:data<=-16'd10470;
      129702:data<=-16'd9950;
      129703:data<=-16'd9635;
      129704:data<=-16'd9095;
      129705:data<=-16'd8933;
      129706:data<=-16'd9274;
      129707:data<=-16'd8900;
      129708:data<=-16'd8752;
      129709:data<=-16'd9605;
      129710:data<=-16'd10290;
      129711:data<=-16'd12028;
      129712:data<=-16'd14336;
      129713:data<=-16'd13609;
      129714:data<=-16'd12326;
      129715:data<=-16'd12800;
      129716:data<=-16'd12019;
      129717:data<=-16'd11388;
      129718:data<=-16'd11119;
      129719:data<=-16'd9768;
      129720:data<=-16'd10219;
      129721:data<=-16'd9620;
      129722:data<=-16'd8696;
      129723:data<=-16'd10825;
      129724:data<=-16'd4799;
      129725:data<=16'd5984;
      129726:data<=16'd5362;
      129727:data<=16'd2776;
      129728:data<=16'd4951;
      129729:data<=16'd3512;
      129730:data<=16'd2605;
      129731:data<=16'd3595;
      129732:data<=16'd2748;
      129733:data<=16'd3055;
      129734:data<=16'd2924;
      129735:data<=16'd2323;
      129736:data<=16'd2972;
      129737:data<=16'd2296;
      129738:data<=16'd2302;
      129739:data<=16'd2570;
      129740:data<=16'd1369;
      129741:data<=16'd1519;
      129742:data<=16'd567;
      129743:data<=-16'd1356;
      129744:data<=-16'd1115;
      129745:data<=-16'd1527;
      129746:data<=-16'd1497;
      129747:data<=-16'd444;
      129748:data<=-16'd1221;
      129749:data<=-16'd1583;
      129750:data<=-16'd1839;
      129751:data<=-16'd2373;
      129752:data<=-16'd1256;
      129753:data<=-16'd1654;
      129754:data<=-16'd2590;
      129755:data<=-16'd1063;
      129756:data<=16'd819;
      129757:data<=16'd2669;
      129758:data<=16'd1997;
      129759:data<=-16'd525;
      129760:data<=16'd490;
      129761:data<=-16'd2532;
      129762:data<=-16'd12991;
      129763:data<=-16'd17356;
      129764:data<=-16'd15076;
      129765:data<=-16'd15109;
      129766:data<=-16'd14880;
      129767:data<=-16'd13540;
      129768:data<=-16'd13773;
      129769:data<=-16'd12972;
      129770:data<=-16'd11822;
      129771:data<=-16'd12346;
      129772:data<=-16'd12296;
      129773:data<=-16'd11511;
      129774:data<=-16'd10966;
      129775:data<=-16'd10851;
      129776:data<=-16'd11724;
      129777:data<=-16'd11855;
      129778:data<=-16'd10912;
      129779:data<=-16'd10599;
      129780:data<=-16'd10223;
      129781:data<=-16'd9796;
      129782:data<=-16'd9577;
      129783:data<=-16'd9132;
      129784:data<=-16'd9162;
      129785:data<=-16'd8739;
      129786:data<=-16'd8088;
      129787:data<=-16'd7671;
      129788:data<=-16'd6126;
      129789:data<=-16'd6250;
      129790:data<=-16'd7162;
      129791:data<=-16'd5730;
      129792:data<=-16'd6514;
      129793:data<=-16'd7532;
      129794:data<=-16'd6065;
      129795:data<=-16'd7087;
      129796:data<=-16'd6273;
      129797:data<=-16'd4777;
      129798:data<=-16'd7351;
      129799:data<=-16'd1265;
      129800:data<=16'd9121;
      129801:data<=16'd7494;
      129802:data<=16'd4535;
      129803:data<=16'd6196;
      129804:data<=16'd4945;
      129805:data<=16'd4722;
      129806:data<=16'd5386;
      129807:data<=16'd4407;
      129808:data<=16'd4843;
      129809:data<=16'd3967;
      129810:data<=16'd2291;
      129811:data<=16'd2617;
      129812:data<=16'd2379;
      129813:data<=16'd2284;
      129814:data<=16'd2444;
      129815:data<=16'd1812;
      129816:data<=16'd2164;
      129817:data<=16'd2267;
      129818:data<=16'd1873;
      129819:data<=16'd1873;
      129820:data<=16'd1242;
      129821:data<=16'd1613;
      129822:data<=16'd2315;
      129823:data<=16'd1774;
      129824:data<=16'd1815;
      129825:data<=16'd591;
      129826:data<=-16'd1742;
      129827:data<=-16'd1656;
      129828:data<=-16'd1307;
      129829:data<=-16'd1577;
      129830:data<=-16'd1300;
      129831:data<=-16'd1753;
      129832:data<=-16'd1521;
      129833:data<=-16'd1177;
      129834:data<=-16'd1456;
      129835:data<=16'd259;
      129836:data<=-16'd2581;
      129837:data<=-16'd12806;
      129838:data<=-16'd17559;
      129839:data<=-16'd15374;
      129840:data<=-16'd15013;
      129841:data<=-16'd14504;
      129842:data<=-16'd14137;
      129843:data<=-16'd16073;
      129844:data<=-16'd14375;
      129845:data<=-16'd10336;
      129846:data<=-16'd9233;
      129847:data<=-16'd8580;
      129848:data<=-16'd7952;
      129849:data<=-16'd8366;
      129850:data<=-16'd8008;
      129851:data<=-16'd7148;
      129852:data<=-16'd6291;
      129853:data<=-16'd5947;
      129854:data<=-16'd6208;
      129855:data<=-16'd5403;
      129856:data<=-16'd4440;
      129857:data<=-16'd4112;
      129858:data<=-16'd4059;
      129859:data<=-16'd5143;
      129860:data<=-16'd5705;
      129861:data<=-16'd5360;
      129862:data<=-16'd5221;
      129863:data<=-16'd3888;
      129864:data<=-16'd2975;
      129865:data<=-16'd2508;
      129866:data<=-16'd720;
      129867:data<=-16'd899;
      129868:data<=-16'd1072;
      129869:data<=16'd699;
      129870:data<=16'd212;
      129871:data<=16'd907;
      129872:data<=16'd1695;
      129873:data<=-16'd1387;
      129874:data<=16'd3256;
      129875:data<=16'd13658;
      129876:data<=16'd14296;
      129877:data<=16'd11614;
      129878:data<=16'd12428;
      129879:data<=16'd11188;
      129880:data<=16'd10622;
      129881:data<=16'd11499;
      129882:data<=16'd10604;
      129883:data<=16'd10519;
      129884:data<=16'd10734;
      129885:data<=16'd10017;
      129886:data<=16'd9812;
      129887:data<=16'd9885;
      129888:data<=16'd10154;
      129889:data<=16'd8448;
      129890:data<=16'd5169;
      129891:data<=16'd4607;
      129892:data<=16'd4053;
      129893:data<=16'd2085;
      129894:data<=16'd2353;
      129895:data<=16'd2516;
      129896:data<=16'd1898;
      129897:data<=16'd2764;
      129898:data<=16'd2784;
      129899:data<=16'd2264;
      129900:data<=16'd2402;
      129901:data<=16'd1905;
      129902:data<=16'd2071;
      129903:data<=16'd2789;
      129904:data<=16'd2848;
      129905:data<=16'd2669;
      129906:data<=16'd1992;
      129907:data<=16'd2197;
      129908:data<=16'd2578;
      129909:data<=16'd1569;
      129910:data<=16'd1745;
      129911:data<=-16'd1071;
      129912:data<=-16'd9996;
      129913:data<=-16'd14366;
      129914:data<=-16'd12026;
      129915:data<=-16'd11637;
      129916:data<=-16'd11961;
      129917:data<=-16'd10715;
      129918:data<=-16'd10433;
      129919:data<=-16'd9688;
      129920:data<=-16'd8316;
      129921:data<=-16'd8257;
      129922:data<=-16'd8348;
      129923:data<=-16'd7494;
      129924:data<=-16'd6213;
      129925:data<=-16'd5958;
      129926:data<=-16'd6983;
      129927:data<=-16'd7174;
      129928:data<=-16'd6796;
      129929:data<=-16'd6798;
      129930:data<=-16'd5773;
      129931:data<=-16'd4925;
      129932:data<=-16'd5477;
      129933:data<=-16'd4739;
      129934:data<=-16'd2140;
      129935:data<=-16'd141;
      129936:data<=16'd252;
      129937:data<=16'd482;
      129938:data<=16'd1580;
      129939:data<=16'd1556;
      129940:data<=16'd886;
      129941:data<=16'd1780;
      129942:data<=16'd1472;
      129943:data<=16'd397;
      129944:data<=16'd1192;
      129945:data<=16'd869;
      129946:data<=16'd1230;
      129947:data<=16'd2746;
      129948:data<=16'd757;
      129949:data<=16'd4200;
      129950:data<=16'd15057;
      129951:data<=16'd17452;
      129952:data<=16'd14204;
      129953:data<=16'd15165;
      129954:data<=16'd14425;
      129955:data<=16'd13066;
      129956:data<=16'd14363;
      129957:data<=16'd13664;
      129958:data<=16'd12915;
      129959:data<=16'd13374;
      129960:data<=16'd12672;
      129961:data<=16'd12622;
      129962:data<=16'd12595;
      129963:data<=16'd11671;
      129964:data<=16'd11157;
      129965:data<=16'd10478;
      129966:data<=16'd10116;
      129967:data<=16'd10255;
      129968:data<=16'd10085;
      129969:data<=16'd9644;
      129970:data<=16'd8921;
      129971:data<=16'd9127;
      129972:data<=16'd9406;
      129973:data<=16'd8687;
      129974:data<=16'd8869;
      129975:data<=16'd8625;
      129976:data<=16'd8658;
      129977:data<=16'd10748;
      129978:data<=16'd9335;
      129979:data<=16'd5238;
      129980:data<=16'd4279;
      129981:data<=16'd4197;
      129982:data<=16'd4040;
      129983:data<=16'd3789;
      129984:data<=16'd2661;
      129985:data<=16'd3621;
      129986:data<=16'd1821;
      129987:data<=-16'd6363;
      129988:data<=-16'd11033;
      129989:data<=-16'd9800;
      129990:data<=-16'd9276;
      129991:data<=-16'd9288;
      129992:data<=-16'd8351;
      129993:data<=-16'd7098;
      129994:data<=-16'd5615;
      129995:data<=-16'd4775;
      129996:data<=-16'd4758;
      129997:data<=-16'd4942;
      129998:data<=-16'd4657;
      129999:data<=-16'd3929;
      130000:data<=-16'd3912;
      130001:data<=-16'd4047;
      130002:data<=-16'd3559;
      130003:data<=-16'd3360;
      130004:data<=-16'd3066;
      130005:data<=-16'd2285;
      130006:data<=-16'd1891;
      130007:data<=-16'd1783;
      130008:data<=-16'd1742;
      130009:data<=-16'd1246;
      130010:data<=16'd340;
      130011:data<=16'd1192;
      130012:data<=16'd887;
      130013:data<=16'd1418;
      130014:data<=16'd1569;
      130015:data<=16'd917;
      130016:data<=16'd1430;
      130017:data<=16'd1666;
      130018:data<=16'd1712;
      130019:data<=16'd2666;
      130020:data<=16'd2416;
      130021:data<=16'd2572;
      130022:data<=16'd2779;
      130023:data<=16'd2030;
      130024:data<=16'd8960;
      130025:data<=16'd20027;
      130026:data<=16'd21643;
      130027:data<=16'd20151;
      130028:data<=16'd21714;
      130029:data<=16'd20225;
      130030:data<=16'd18812;
      130031:data<=16'd19294;
      130032:data<=16'd17775;
      130033:data<=16'd16976;
      130034:data<=16'd17106;
      130035:data<=16'd16166;
      130036:data<=16'd15465;
      130037:data<=16'd14800;
      130038:data<=16'd14504;
      130039:data<=16'd14178;
      130040:data<=16'd12909;
      130041:data<=16'd12232;
      130042:data<=16'd11941;
      130043:data<=16'd12195;
      130044:data<=16'd12868;
      130045:data<=16'd12052;
      130046:data<=16'd11819;
      130047:data<=16'd12339;
      130048:data<=16'd11403;
      130049:data<=16'd10975;
      130050:data<=16'd10654;
      130051:data<=16'd9847;
      130052:data<=16'd10158;
      130053:data<=16'd9483;
      130054:data<=16'd8059;
      130055:data<=16'd7444;
      130056:data<=16'd6596;
      130057:data<=16'd6721;
      130058:data<=16'd6570;
      130059:data<=16'd5899;
      130060:data<=16'd7830;
      130061:data<=16'd6061;
      130062:data<=-16'd2458;
      130063:data<=-16'd7388;
      130064:data<=-16'd7009;
      130065:data<=-16'd7153;
      130066:data<=-16'd6924;
      130067:data<=-16'd7077;
      130068:data<=-16'd9638;
      130069:data<=-16'd11166;
      130070:data<=-16'd10495;
      130071:data<=-16'd10102;
      130072:data<=-16'd9962;
      130073:data<=-16'd9321;
      130074:data<=-16'd8947;
      130075:data<=-16'd8912;
      130076:data<=-16'd7811;
      130077:data<=-16'd5667;
      130078:data<=-16'd4958;
      130079:data<=-16'd5670;
      130080:data<=-16'd5436;
      130081:data<=-16'd5071;
      130082:data<=-16'd5277;
      130083:data<=-16'd4877;
      130084:data<=-16'd4981;
      130085:data<=-16'd5612;
      130086:data<=-16'd5354;
      130087:data<=-16'd4892;
      130088:data<=-16'd4478;
      130089:data<=-16'd4607;
      130090:data<=-16'd5171;
      130091:data<=-16'd4478;
      130092:data<=-16'd3598;
      130093:data<=-16'd2411;
      130094:data<=-16'd505;
      130095:data<=-16'd532;
      130096:data<=-16'd150;
      130097:data<=16'd511;
      130098:data<=-16'd1733;
      130099:data<=16'd1736;
      130100:data<=16'd11338;
      130101:data<=16'd13585;
      130102:data<=16'd11110;
      130103:data<=16'd11462;
      130104:data<=16'd10619;
      130105:data<=16'd9491;
      130106:data<=16'd10226;
      130107:data<=16'd9394;
      130108:data<=16'd8222;
      130109:data<=16'd9188;
      130110:data<=16'd10100;
      130111:data<=16'd9577;
      130112:data<=16'd10196;
      130113:data<=16'd12562;
      130114:data<=16'd12800;
      130115:data<=16'd11386;
      130116:data<=16'd11209;
      130117:data<=16'd10449;
      130118:data<=16'd9373;
      130119:data<=16'd9242;
      130120:data<=16'd8379;
      130121:data<=16'd7779;
      130122:data<=16'd7888;
      130123:data<=16'd7388;
      130124:data<=16'd7115;
      130125:data<=16'd6836;
      130126:data<=16'd7057;
      130127:data<=16'd8554;
      130128:data<=16'd8778;
      130129:data<=16'd7862;
      130130:data<=16'd7080;
      130131:data<=16'd5617;
      130132:data<=16'd4907;
      130133:data<=16'd4435;
      130134:data<=16'd3263;
      130135:data<=16'd3889;
      130136:data<=16'd2061;
      130137:data<=-16'd5962;
      130138:data<=-16'd11477;
      130139:data<=-16'd10795;
      130140:data<=-16'd10366;
      130141:data<=-16'd10871;
      130142:data<=-16'd10146;
      130143:data<=-16'd9080;
      130144:data<=-16'd7633;
      130145:data<=-16'd6730;
      130146:data<=-16'd7080;
      130147:data<=-16'd7092;
      130148:data<=-16'd6740;
      130149:data<=-16'd6407;
      130150:data<=-16'd6196;
      130151:data<=-16'd6554;
      130152:data<=-16'd6337;
      130153:data<=-16'd6034;
      130154:data<=-16'd6285;
      130155:data<=-16'd5521;
      130156:data<=-16'd5997;
      130157:data<=-16'd9022;
      130158:data<=-16'd10660;
      130159:data<=-16'd10041;
      130160:data<=-16'd8573;
      130161:data<=-16'd7453;
      130162:data<=-16'd7703;
      130163:data<=-16'd7420;
      130164:data<=-16'd7326;
      130165:data<=-16'd8484;
      130166:data<=-16'd7632;
      130167:data<=-16'd6176;
      130168:data<=-16'd5877;
      130169:data<=-16'd5278;
      130170:data<=-16'd6032;
      130171:data<=-16'd5729;
      130172:data<=-16'd4193;
      130173:data<=-16'd6056;
      130174:data<=-16'd3225;
      130175:data<=16'd6357;
      130176:data<=16'd9447;
      130177:data<=16'd8109;
      130178:data<=16'd9321;
      130179:data<=16'd8678;
      130180:data<=16'd7832;
      130181:data<=16'd8463;
      130182:data<=16'd7203;
      130183:data<=16'd6522;
      130184:data<=16'd6799;
      130185:data<=16'd5937;
      130186:data<=16'd5686;
      130187:data<=16'd5630;
      130188:data<=16'd4702;
      130189:data<=16'd3802;
      130190:data<=16'd3369;
      130191:data<=16'd3365;
      130192:data<=16'd2990;
      130193:data<=16'd3124;
      130194:data<=16'd3962;
      130195:data<=16'd3468;
      130196:data<=16'd3362;
      130197:data<=16'd4300;
      130198:data<=16'd3820;
      130199:data<=16'd2864;
      130200:data<=16'd2165;
      130201:data<=16'd3007;
      130202:data<=16'd6658;
      130203:data<=16'd8088;
      130204:data<=16'd6167;
      130205:data<=16'd5001;
      130206:data<=16'd4161;
      130207:data<=16'd3727;
      130208:data<=16'd3325;
      130209:data<=16'd2141;
      130210:data<=16'd3595;
      130211:data<=16'd3122;
      130212:data<=-16'd4698;
      130213:data<=-16'd10417;
      130214:data<=-16'd9577;
      130215:data<=-16'd8953;
      130216:data<=-16'd9189;
      130217:data<=-16'd8831;
      130218:data<=-16'd8821;
      130219:data<=-16'd8287;
      130220:data<=-16'd7937;
      130221:data<=-16'd8301;
      130222:data<=-16'd8084;
      130223:data<=-16'd7865;
      130224:data<=-16'd8026;
      130225:data<=-16'd8046;
      130226:data<=-16'd7917;
      130227:data<=-16'd7479;
      130228:data<=-16'd7413;
      130229:data<=-16'd7391;
      130230:data<=-16'd6526;
      130231:data<=-16'd6678;
      130232:data<=-16'd7410;
      130233:data<=-16'd6699;
      130234:data<=-16'd6548;
      130235:data<=-16'd6802;
      130236:data<=-16'd6003;
      130237:data<=-16'd6349;
      130238:data<=-16'd6678;
      130239:data<=-16'd5912;
      130240:data<=-16'd6757;
      130241:data<=-16'd7160;
      130242:data<=-16'd5958;
      130243:data<=-16'd5953;
      130244:data<=-16'd6385;
      130245:data<=-16'd7153;
      130246:data<=-16'd8622;
      130247:data<=-16'd10410;
      130248:data<=-16'd12815;
      130249:data<=-16'd8994;
      130250:data<=16'd1098;
      130251:data<=16'd4009;
      130252:data<=16'd1378;
      130253:data<=16'd2249;
      130254:data<=16'd2218;
      130255:data<=16'd1339;
      130256:data<=16'd2552;
      130257:data<=16'd1700;
      130258:data<=16'd622;
      130259:data<=16'd1445;
      130260:data<=16'd250;
      130261:data<=-16'd1968;
      130262:data<=-16'd2422;
      130263:data<=-16'd2300;
      130264:data<=-16'd2564;
      130265:data<=-16'd2569;
      130266:data<=-16'd2466;
      130267:data<=-16'd3065;
      130268:data<=-16'd3087;
      130269:data<=-16'd2366;
      130270:data<=-16'd2692;
      130271:data<=-16'd2952;
      130272:data<=-16'd2678;
      130273:data<=-16'd2793;
      130274:data<=-16'd2622;
      130275:data<=-16'd2701;
      130276:data<=-16'd2722;
      130277:data<=-16'd2766;
      130278:data<=-16'd4197;
      130279:data<=-16'd4496;
      130280:data<=-16'd4293;
      130281:data<=-16'd5724;
      130282:data<=-16'd5013;
      130283:data<=-16'd4140;
      130284:data<=-16'd5588;
      130285:data<=-16'd4402;
      130286:data<=-16'd4793;
      130287:data<=-16'd11852;
      130288:data<=-16'd17403;
      130289:data<=-16'd17443;
      130290:data<=-16'd15640;
      130291:data<=-16'd12875;
      130292:data<=-16'd10803;
      130293:data<=-16'd11288;
      130294:data<=-16'd12243;
      130295:data<=-16'd12146;
      130296:data<=-16'd11925;
      130297:data<=-16'd11370;
      130298:data<=-16'd10219;
      130299:data<=-16'd9831;
      130300:data<=-16'd9826;
      130301:data<=-16'd9250;
      130302:data<=-16'd8943;
      130303:data<=-16'd8693;
      130304:data<=-16'd8188;
      130305:data<=-16'd7999;
      130306:data<=-16'd7699;
      130307:data<=-16'd7225;
      130308:data<=-16'd6934;
      130309:data<=-16'd7019;
      130310:data<=-16'd7498;
      130311:data<=-16'd7726;
      130312:data<=-16'd7887;
      130313:data<=-16'd7946;
      130314:data<=-16'd7674;
      130315:data<=-16'd7691;
      130316:data<=-16'd7210;
      130317:data<=-16'd6279;
      130318:data<=-16'd5638;
      130319:data<=-16'd5037;
      130320:data<=-16'd5407;
      130321:data<=-16'd4754;
      130322:data<=-16'd3341;
      130323:data<=-16'd5159;
      130324:data<=-16'd2499;
      130325:data<=16'd7500;
      130326:data<=16'd10815;
      130327:data<=16'd7585;
      130328:data<=16'd7169;
      130329:data<=16'd6595;
      130330:data<=16'd6002;
      130331:data<=16'd7233;
      130332:data<=16'd6347;
      130333:data<=16'd5435;
      130334:data<=16'd6065;
      130335:data<=16'd4273;
      130336:data<=16'd1304;
      130337:data<=16'd566;
      130338:data<=16'd873;
      130339:data<=16'd376;
      130340:data<=16'd74;
      130341:data<=16'd693;
      130342:data<=16'd781;
      130343:data<=-16'd14;
      130344:data<=-16'd1119;
      130345:data<=-16'd1853;
      130346:data<=-16'd1389;
      130347:data<=-16'd1063;
      130348:data<=-16'd1509;
      130349:data<=-16'd1492;
      130350:data<=-16'd1145;
      130351:data<=-16'd588;
      130352:data<=16'd18;
      130353:data<=16'd276;
      130354:data<=16'd435;
      130355:data<=-16'd165;
      130356:data<=-16'd945;
      130357:data<=-16'd775;
      130358:data<=-16'd655;
      130359:data<=-16'd405;
      130360:data<=-16'd153;
      130361:data<=-16'd3030;
      130362:data<=-16'd10035;
      130363:data<=-16'd15898;
      130364:data<=-16'd15667;
      130365:data<=-16'd13700;
      130366:data<=-16'd14237;
      130367:data<=-16'd13769;
      130368:data<=-16'd12395;
      130369:data<=-16'd11956;
      130370:data<=-16'd10801;
      130371:data<=-16'd10313;
      130372:data<=-16'd10178;
      130373:data<=-16'd8746;
      130374:data<=-16'd8436;
      130375:data<=-16'd8410;
      130376:data<=-16'd7338;
      130377:data<=-16'd7544;
      130378:data<=-16'd8492;
      130379:data<=-16'd7723;
      130380:data<=-16'd4830;
      130381:data<=-16'd2769;
      130382:data<=-16'd3098;
      130383:data<=-16'd2599;
      130384:data<=-16'd1633;
      130385:data<=-16'd1644;
      130386:data<=-16'd814;
      130387:data<=-16'd558;
      130388:data<=-16'd776;
      130389:data<=-16'd118;
      130390:data<=-16'd500;
      130391:data<=-16'd522;
      130392:data<=16'd526;
      130393:data<=16'd883;
      130394:data<=16'd635;
      130395:data<=-16'd801;
      130396:data<=-16'd561;
      130397:data<=16'd978;
      130398:data<=-16'd923;
      130399:data<=16'd1973;
      130400:data<=16'd12119;
      130401:data<=16'd15417;
      130402:data<=16'd12944;
      130403:data<=16'd13624;
      130404:data<=16'd13556;
      130405:data<=16'd12022;
      130406:data<=16'd12348;
      130407:data<=16'd12575;
      130408:data<=16'd12269;
      130409:data<=16'd12019;
      130410:data<=16'd10423;
      130411:data<=16'd8654;
      130412:data<=16'd8728;
      130413:data<=16'd8846;
      130414:data<=16'd7873;
      130415:data<=16'd7645;
      130416:data<=16'd7686;
      130417:data<=16'd7322;
      130418:data<=16'd7345;
      130419:data<=16'd7012;
      130420:data<=16'd6972;
      130421:data<=16'd7233;
      130422:data<=16'd6532;
      130423:data<=16'd6431;
      130424:data<=16'd5441;
      130425:data<=16'd2444;
      130426:data<=16'd1791;
      130427:data<=16'd2364;
      130428:data<=16'd1119;
      130429:data<=16'd493;
      130430:data<=16'd538;
      130431:data<=16'd311;
      130432:data<=16'd741;
      130433:data<=16'd658;
      130434:data<=16'd14;
      130435:data<=16'd619;
      130436:data<=16'd64;
      130437:data<=-16'd5771;
      130438:data<=-16'd12531;
      130439:data<=-16'd13273;
      130440:data<=-16'd11523;
      130441:data<=-16'd11154;
      130442:data<=-16'd10066;
      130443:data<=-16'd9664;
      130444:data<=-16'd10445;
      130445:data<=-16'd10528;
      130446:data<=-16'd10605;
      130447:data<=-16'd9752;
      130448:data<=-16'd8382;
      130449:data<=-16'd8275;
      130450:data<=-16'd7879;
      130451:data<=-16'd7272;
      130452:data<=-16'd7051;
      130453:data<=-16'd6581;
      130454:data<=-16'd6106;
      130455:data<=-16'd4989;
      130456:data<=-16'd4507;
      130457:data<=-16'd4943;
      130458:data<=-16'd4067;
      130459:data<=-16'd3692;
      130460:data<=-16'd3958;
      130461:data<=-16'd3595;
      130462:data<=-16'd4458;
      130463:data<=-16'd4661;
      130464:data<=-16'd3982;
      130465:data<=-16'd4182;
      130466:data<=-16'd3112;
      130467:data<=-16'd2805;
      130468:data<=-16'd2708;
      130469:data<=16'd705;
      130470:data<=16'd2315;
      130471:data<=16'd2326;
      130472:data<=16'd3466;
      130473:data<=16'd1889;
      130474:data<=16'd4726;
      130475:data<=16'd14756;
      130476:data<=16'd18125;
      130477:data<=16'd14998;
      130478:data<=16'd14566;
      130479:data<=16'd14475;
      130480:data<=16'd13606;
      130481:data<=16'd13849;
      130482:data<=16'd13527;
      130483:data<=16'd12721;
      130484:data<=16'd12407;
      130485:data<=16'd12266;
      130486:data<=16'd12041;
      130487:data<=16'd11503;
      130488:data<=16'd10969;
      130489:data<=16'd10616;
      130490:data<=16'd10496;
      130491:data<=16'd10669;
      130492:data<=16'd10334;
      130493:data<=16'd9746;
      130494:data<=16'd9677;
      130495:data<=16'd9471;
      130496:data<=16'd9348;
      130497:data<=16'd9633;
      130498:data<=16'd9121;
      130499:data<=16'd8407;
      130500:data<=16'd8539;
      130501:data<=16'd8367;
      130502:data<=16'd8072;
      130503:data<=16'd8234;
      130504:data<=16'd7923;
      130505:data<=16'd7530;
      130506:data<=16'd7112;
      130507:data<=16'd6590;
      130508:data<=16'd7028;
      130509:data<=16'd6845;
      130510:data<=16'd6302;
      130511:data<=16'd6690;
      130512:data<=16'd2481;
      130513:data<=-16'd5971;
      130514:data<=-16'd9706;
      130515:data<=-16'd9279;
      130516:data<=-16'd9229;
      130517:data<=-16'd8724;
      130518:data<=-16'd8393;
      130519:data<=-16'd8363;
      130520:data<=-16'd7732;
      130521:data<=-16'd7395;
      130522:data<=-16'd6749;
      130523:data<=-16'd6143;
      130524:data<=-16'd6260;
      130525:data<=-16'd5797;
      130526:data<=-16'd5366;
      130527:data<=-16'd4642;
      130528:data<=-16'd2811;
      130529:data<=-16'd2008;
      130530:data<=-16'd1974;
      130531:data<=-16'd1641;
      130532:data<=-16'd1412;
      130533:data<=-16'd634;
      130534:data<=-16'd813;
      130535:data<=-16'd1876;
      130536:data<=-16'd1149;
      130537:data<=-16'd485;
      130538:data<=-16'd610;
      130539:data<=-16'd47;
      130540:data<=-16'd218;
      130541:data<=-16'd479;
      130542:data<=-16'd361;
      130543:data<=-16'd381;
      130544:data<=16'd1206;
      130545:data<=16'd2353;
      130546:data<=16'd2426;
      130547:data<=16'd3084;
      130548:data<=16'd1626;
      130549:data<=16'd3762;
      130550:data<=16'd13417;
      130551:data<=16'd17323;
      130552:data<=16'd14240;
      130553:data<=16'd14973;
      130554:data<=16'd16299;
      130555:data<=16'd15854;
      130556:data<=16'd16269;
      130557:data<=16'd15158;
      130558:data<=16'd15048;
      130559:data<=16'd16659;
      130560:data<=16'd15711;
      130561:data<=16'd15262;
      130562:data<=16'd16478;
      130563:data<=16'd16083;
      130564:data<=16'd15347;
      130565:data<=16'd14543;
      130566:data<=16'd13446;
      130567:data<=16'd13406;
      130568:data<=16'd13033;
      130569:data<=16'd12185;
      130570:data<=16'd12157;
      130571:data<=16'd12208;
      130572:data<=16'd11674;
      130573:data<=16'd10528;
      130574:data<=16'd10075;
      130575:data<=16'd10621;
      130576:data<=16'd10011;
      130577:data<=16'd9230;
      130578:data<=16'd9818;
      130579:data<=16'd10061;
      130580:data<=16'd9705;
      130581:data<=16'd8978;
      130582:data<=16'd8020;
      130583:data<=16'd7921;
      130584:data<=16'd7376;
      130585:data<=16'd6965;
      130586:data<=16'd7188;
      130587:data<=16'd2017;
      130588:data<=-16'd6414;
      130589:data<=-16'd8088;
      130590:data<=-16'd6132;
      130591:data<=-16'd6586;
      130592:data<=-16'd6546;
      130593:data<=-16'd6387;
      130594:data<=-16'd6546;
      130595:data<=-16'd4919;
      130596:data<=-16'd4319;
      130597:data<=-16'd4640;
      130598:data<=-16'd3680;
      130599:data<=-16'd3580;
      130600:data<=-16'd3595;
      130601:data<=-16'd3005;
      130602:data<=-16'd3908;
      130603:data<=-16'd5124;
      130604:data<=-16'd5618;
      130605:data<=-16'd5535;
      130606:data<=-16'd5018;
      130607:data<=-16'd5175;
      130608:data<=-16'd5095;
      130609:data<=-16'd5081;
      130610:data<=-16'd5697;
      130611:data<=-16'd4625;
      130612:data<=-16'd3354;
      130613:data<=-16'd3310;
      130614:data<=-16'd2893;
      130615:data<=-16'd2937;
      130616:data<=-16'd2874;
      130617:data<=-16'd2590;
      130618:data<=-16'd2795;
      130619:data<=-16'd1782;
      130620:data<=-16'd1842;
      130621:data<=-16'd2469;
      130622:data<=-16'd1389;
      130623:data<=-16'd2778;
      130624:data<=-16'd506;
      130625:data<=16'd9344;
      130626:data<=16'd12548;
      130627:data<=16'd9662;
      130628:data<=16'd11188;
      130629:data<=16'd12237;
      130630:data<=16'd11556;
      130631:data<=16'd11926;
      130632:data<=16'd10875;
      130633:data<=16'd10604;
      130634:data<=16'd10880;
      130635:data<=16'd9303;
      130636:data<=16'd8924;
      130637:data<=16'd9063;
      130638:data<=16'd7958;
      130639:data<=16'd7417;
      130640:data<=16'd7147;
      130641:data<=16'd7050;
      130642:data<=16'd7030;
      130643:data<=16'd5961;
      130644:data<=16'd5648;
      130645:data<=16'd6746;
      130646:data<=16'd7166;
      130647:data<=16'd7464;
      130648:data<=16'd8487;
      130649:data<=16'd8705;
      130650:data<=16'd8270;
      130651:data<=16'd8152;
      130652:data<=16'd7497;
      130653:data<=16'd6539;
      130654:data<=16'd6226;
      130655:data<=16'd6094;
      130656:data<=16'd5570;
      130657:data<=16'd4749;
      130658:data<=16'd4399;
      130659:data<=16'd3753;
      130660:data<=16'd3030;
      130661:data<=16'd4184;
      130662:data<=16'd1495;
      130663:data<=-16'd6724;
      130664:data<=-16'd9253;
      130665:data<=-16'd7057;
      130666:data<=-16'd7961;
      130667:data<=-16'd7696;
      130668:data<=-16'd6983;
      130669:data<=-16'd8525;
      130670:data<=-16'd8210;
      130671:data<=-16'd7946;
      130672:data<=-16'd8311;
      130673:data<=-16'd7594;
      130674:data<=-16'd8117;
      130675:data<=-16'd7764;
      130676:data<=-16'd7028;
      130677:data<=-16'd7899;
      130678:data<=-16'd6570;
      130679:data<=-16'd4963;
      130680:data<=-16'd4811;
      130681:data<=-16'd3946;
      130682:data<=-16'd4710;
      130683:data<=-16'd5685;
      130684:data<=-16'd5209;
      130685:data<=-16'd5676;
      130686:data<=-16'd5520;
      130687:data<=-16'd5006;
      130688:data<=-16'd5438;
      130689:data<=-16'd5382;
      130690:data<=-16'd5087;
      130691:data<=-16'd4623;
      130692:data<=-16'd5560;
      130693:data<=-16'd7121;
      130694:data<=-16'd6072;
      130695:data<=-16'd5577;
      130696:data<=-16'd4968;
      130697:data<=-16'd3427;
      130698:data<=-16'd5603;
      130699:data<=-16'd3190;
      130700:data<=16'd6396;
      130701:data<=16'd9224;
      130702:data<=16'd7012;
      130703:data<=16'd7426;
      130704:data<=16'd7289;
      130705:data<=16'd6945;
      130706:data<=16'd6578;
      130707:data<=16'd5319;
      130708:data<=16'd5533;
      130709:data<=16'd5456;
      130710:data<=16'd4529;
      130711:data<=16'd4978;
      130712:data<=16'd5673;
      130713:data<=16'd5870;
      130714:data<=16'd5752;
      130715:data<=16'd5143;
      130716:data<=16'd4525;
      130717:data<=16'd4081;
      130718:data<=16'd3727;
      130719:data<=16'd3356;
      130720:data<=16'd3483;
      130721:data<=16'd3563;
      130722:data<=16'd2590;
      130723:data<=16'd2115;
      130724:data<=16'd2103;
      130725:data<=16'd1494;
      130726:data<=16'd1178;
      130727:data<=16'd614;
      130728:data<=16'd422;
      130729:data<=16'd1745;
      130730:data<=16'd2566;
      130731:data<=16'd1909;
      130732:data<=16'd1030;
      130733:data<=16'd1260;
      130734:data<=16'd1071;
      130735:data<=-16'd61;
      130736:data<=16'd1256;
      130737:data<=-16'd761;
      130738:data<=-16'd9520;
      130739:data<=-16'd12536;
      130740:data<=-16'd9928;
      130741:data<=-16'd10901;
      130742:data<=-16'd10986;
      130743:data<=-16'd9791;
      130744:data<=-16'd10257;
      130745:data<=-16'd9118;
      130746:data<=-16'd8066;
      130747:data<=-16'd7864;
      130748:data<=-16'd7377;
      130749:data<=-16'd7944;
      130750:data<=-16'd7720;
      130751:data<=-16'd7295;
      130752:data<=-16'd7447;
      130753:data<=-16'd6542;
      130754:data<=-16'd6733;
      130755:data<=-16'd7068;
      130756:data<=-16'd6366;
      130757:data<=-16'd6816;
      130758:data<=-16'd6915;
      130759:data<=-16'd6907;
      130760:data<=-16'd6966;
      130761:data<=-16'd5792;
      130762:data<=-16'd5950;
      130763:data<=-16'd6037;
      130764:data<=-16'd5477;
      130765:data<=-16'd6458;
      130766:data<=-16'd5808;
      130767:data<=-16'd5194;
      130768:data<=-16'd6028;
      130769:data<=-16'd5013;
      130770:data<=-16'd5409;
      130771:data<=-16'd5533;
      130772:data<=-16'd4100;
      130773:data<=-16'd6614;
      130774:data<=-16'd4349;
      130775:data<=16'd5309;
      130776:data<=16'd8555;
      130777:data<=16'd7247;
      130778:data<=16'd6868;
      130779:data<=16'd4382;
      130780:data<=16'd3594;
      130781:data<=16'd3903;
      130782:data<=16'd1923;
      130783:data<=16'd1895;
      130784:data<=16'd2340;
      130785:data<=16'd873;
      130786:data<=16'd1011;
      130787:data<=16'd1463;
      130788:data<=16'd837;
      130789:data<=16'd725;
      130790:data<=16'd3;
      130791:data<=-16'd441;
      130792:data<=16'd338;
      130793:data<=16'd152;
      130794:data<=-16'd91;
      130795:data<=-16'd193;
      130796:data<=-16'd1794;
      130797:data<=-16'd2502;
      130798:data<=-16'd2379;
      130799:data<=-16'd2960;
      130800:data<=-16'd2252;
      130801:data<=-16'd1895;
      130802:data<=-16'd2648;
      130803:data<=-16'd2337;
      130804:data<=-16'd2722;
      130805:data<=-16'd2692;
      130806:data<=-16'd1920;
      130807:data<=-16'd3251;
      130808:data<=-16'd3275;
      130809:data<=-16'd2792;
      130810:data<=-16'd3250;
      130811:data<=-16'd1028;
      130812:data<=-16'd5150;
      130813:data<=-16'd16287;
      130814:data<=-16'd18440;
      130815:data<=-16'd15506;
      130816:data<=-16'd16139;
      130817:data<=-16'd15133;
      130818:data<=-16'd14186;
      130819:data<=-16'd14407;
      130820:data<=-16'd13341;
      130821:data<=-16'd13584;
      130822:data<=-16'd13342;
      130823:data<=-16'd12420;
      130824:data<=-16'd12834;
      130825:data<=-16'd11411;
      130826:data<=-16'd9342;
      130827:data<=-16'd8457;
      130828:data<=-16'd7928;
      130829:data<=-16'd9033;
      130830:data<=-16'd9312;
      130831:data<=-16'd8325;
      130832:data<=-16'd8760;
      130833:data<=-16'd8432;
      130834:data<=-16'd7809;
      130835:data<=-16'd8217;
      130836:data<=-16'd7653;
      130837:data<=-16'd7162;
      130838:data<=-16'd6951;
      130839:data<=-16'd6467;
      130840:data<=-16'd6467;
      130841:data<=-16'd5888;
      130842:data<=-16'd5670;
      130843:data<=-16'd5371;
      130844:data<=-16'd3780;
      130845:data<=-16'd4585;
      130846:data<=-16'd5970;
      130847:data<=-16'd5436;
      130848:data<=-16'd6681;
      130849:data<=-16'd4167;
      130850:data<=16'd4877;
      130851:data<=16'd8865;
      130852:data<=16'd7300;
      130853:data<=16'd7808;
      130854:data<=16'd7715;
      130855:data<=16'd6625;
      130856:data<=16'd7266;
      130857:data<=16'd7151;
      130858:data<=16'd6855;
      130859:data<=16'd7418;
      130860:data<=16'd6927;
      130861:data<=16'd6601;
      130862:data<=16'd5943;
      130863:data<=16'd3786;
      130864:data<=16'd3095;
      130865:data<=16'd3424;
      130866:data<=16'd3183;
      130867:data<=16'd3479;
      130868:data<=16'd3457;
      130869:data<=16'd3301;
      130870:data<=16'd2870;
      130871:data<=16'd1128;
      130872:data<=16'd983;
      130873:data<=16'd1868;
      130874:data<=16'd1406;
      130875:data<=16'd1630;
      130876:data<=16'd1485;
      130877:data<=16'd869;
      130878:data<=16'd1236;
      130879:data<=-16'd183;
      130880:data<=-16'd1236;
      130881:data<=-16'd546;
      130882:data<=-16'd1206;
      130883:data<=-16'd597;
      130884:data<=-16'd359;
      130885:data<=-16'd1600;
      130886:data<=16'd566;
      130887:data<=-16'd2513;
      130888:data<=-16'd12698;
      130889:data<=-16'd14583;
      130890:data<=-16'd11291;
      130891:data<=-16'd11958;
      130892:data<=-16'd11439;
      130893:data<=-16'd10355;
      130894:data<=-16'd10643;
      130895:data<=-16'd10228;
      130896:data<=-16'd11260;
      130897:data<=-16'd11996;
      130898:data<=-16'd10975;
      130899:data<=-16'd10981;
      130900:data<=-16'd10671;
      130901:data<=-16'd9699;
      130902:data<=-16'd8887;
      130903:data<=-16'd7592;
      130904:data<=-16'd7435;
      130905:data<=-16'd7586;
      130906:data<=-16'd6710;
      130907:data<=-16'd5890;
      130908:data<=-16'd4760;
      130909:data<=-16'd4860;
      130910:data<=-16'd5914;
      130911:data<=-16'd4971;
      130912:data<=-16'd4834;
      130913:data<=-16'd6346;
      130914:data<=-16'd5997;
      130915:data<=-16'd4487;
      130916:data<=-16'd3221;
      130917:data<=-16'd2855;
      130918:data<=-16'd2870;
      130919:data<=-16'd1627;
      130920:data<=-16'd1315;
      130921:data<=-16'd1328;
      130922:data<=-16'd368;
      130923:data<=-16'd1760;
      130924:data<=16'd253;
      130925:data<=16'd9436;
      130926:data<=16'd14049;
      130927:data<=16'd12289;
      130928:data<=16'd12149;
      130929:data<=16'd11382;
      130930:data<=16'd9297;
      130931:data<=16'd9461;
      130932:data<=16'd9688;
      130933:data<=16'd9006;
      130934:data<=16'd8848;
      130935:data<=16'd8792;
      130936:data<=16'd8877;
      130937:data<=16'd8734;
      130938:data<=16'd8005;
      130939:data<=16'd7562;
      130940:data<=16'd7448;
      130941:data<=16'd7413;
      130942:data<=16'd7370;
      130943:data<=16'd7204;
      130944:data<=16'd7151;
      130945:data<=16'd6598;
      130946:data<=16'd5517;
      130947:data<=16'd4927;
      130948:data<=16'd4452;
      130949:data<=16'd4264;
      130950:data<=16'd4804;
      130951:data<=16'd4663;
      130952:data<=16'd4288;
      130953:data<=16'd4440;
      130954:data<=16'd4087;
      130955:data<=16'd4128;
      130956:data<=16'd3864;
      130957:data<=16'd2858;
      130958:data<=16'd3821;
      130959:data<=16'd3168;
      130960:data<=16'd782;
      130961:data<=16'd2585;
      130962:data<=-16'd802;
      130963:data<=-16'd12448;
      130964:data<=-16'd15640;
      130965:data<=-16'd12346;
      130966:data<=-16'd13238;
      130967:data<=-16'd12672;
      130968:data<=-16'd11077;
      130969:data<=-16'd11421;
      130970:data<=-16'd10113;
      130971:data<=-16'd9765;
      130972:data<=-16'd9859;
      130973:data<=-16'd8335;
      130974:data<=-16'd8675;
      130975:data<=-16'd8516;
      130976:data<=-16'd7141;
      130977:data<=-16'd7097;
      130978:data<=-16'd5997;
      130979:data<=-16'd5739;
      130980:data<=-16'd7366;
      130981:data<=-16'd7210;
      130982:data<=-16'd6664;
      130983:data<=-16'd6487;
      130984:data<=-16'd6055;
      130985:data<=-16'd6364;
      130986:data<=-16'd5943;
      130987:data<=-16'd5027;
      130988:data<=-16'd4449;
      130989:data<=-16'd3896;
      130990:data<=-16'd4138;
      130991:data<=-16'd3635;
      130992:data<=-16'd2893;
      130993:data<=-16'd3107;
      130994:data<=-16'd2130;
      130995:data<=-16'd1853;
      130996:data<=-16'd2385;
      130997:data<=-16'd2106;
      130998:data<=-16'd3656;
      130999:data<=-16'd1398;
      131000:data<=16'd7465;
      131001:data<=16'd11715;
      131002:data<=16'd10328;
      131003:data<=16'd10596;
      131004:data<=16'd11643;
      131005:data<=16'd12273;
      131006:data<=16'd12515;
      131007:data<=16'd12091;
      131008:data<=16'd12110;
      131009:data<=16'd11721;
      131010:data<=16'd11239;
      131011:data<=16'd11546;
      131012:data<=16'd10777;
      131013:data<=16'd8963;
      131014:data<=16'd7558;
      131015:data<=16'd6940;
      131016:data<=16'd7101;
      131017:data<=16'd7109;
      131018:data<=16'd6796;
      131019:data<=16'd6692;
      131020:data<=16'd6660;
      131021:data<=16'd7033;
      131022:data<=16'd7423;
      131023:data<=16'd6992;
      131024:data<=16'd6708;
      131025:data<=16'd6957;
      131026:data<=16'd6598;
      131027:data<=16'd6206;
      131028:data<=16'd6369;
      131029:data<=16'd6176;
      131030:data<=16'd6175;
      131031:data<=16'd5803;
      131032:data<=16'd4684;
      131033:data<=16'd5209;
      131034:data<=16'd5071;
      131035:data<=16'd4170;
      131036:data<=16'd6261;
      131037:data<=16'd2692;
      131038:data<=-16'd7873;
      131039:data<=-16'd10302;
      131040:data<=-16'd7162;
      131041:data<=-16'd7935;
      131042:data<=-16'd7683;
      131043:data<=-16'd6426;
      131044:data<=-16'd6686;
      131045:data<=-16'd6261;
      131046:data<=-16'd5647;
      131047:data<=-16'd4134;
      131048:data<=-16'd3692;
      131049:data<=-16'd5632;
      131050:data<=-16'd5203;
      131051:data<=-16'd4334;
      131052:data<=-16'd4915;
      131053:data<=-16'd3800;
      131054:data<=-16'd3119;
      131055:data<=-16'd3245;
      131056:data<=-16'd3042;
      131057:data<=-16'd3389;
      131058:data<=-16'd2557;
      131059:data<=-16'd2209;
      131060:data<=-16'd3031;
      131061:data<=-16'd2349;
      131062:data<=-16'd1710;
      131063:data<=-16'd566;
      131064:data<=16'd869;
      131065:data<=16'd296;
      131066:data<=16'd778;
      131067:data<=16'd1347;
      131068:data<=16'd532;
      131069:data<=16'd1366;
      131070:data<=16'd1539;
      131071:data<=16'd1569;
    endcase
end
assign dout =data;
endmodule
